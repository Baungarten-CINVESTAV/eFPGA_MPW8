magic
tech sky130A
magscale 1 2
timestamp 1672417572
<< viali >>
rect 1777 37417 1811 37451
rect 26341 37417 26375 37451
rect 5825 37349 5859 37383
rect 19441 37349 19475 37383
rect 25789 37349 25823 37383
rect 12357 37281 12391 37315
rect 22017 37281 22051 37315
rect 30665 37281 30699 37315
rect 32321 37281 32355 37315
rect 1593 37213 1627 37247
rect 2881 37213 2915 37247
rect 3985 37213 4019 37247
rect 4905 37213 4939 37247
rect 6009 37213 6043 37247
rect 6561 37213 6595 37247
rect 7941 37213 7975 37247
rect 9413 37213 9447 37247
rect 10241 37213 10275 37247
rect 10885 37213 10919 37247
rect 12633 37213 12667 37247
rect 14473 37213 14507 37247
rect 15117 37213 15151 37247
rect 15577 37213 15611 37247
rect 17049 37213 17083 37247
rect 17509 37213 17543 37247
rect 18705 37213 18739 37247
rect 19625 37213 19659 37247
rect 20085 37213 20119 37247
rect 21005 37213 21039 37247
rect 22293 37213 22327 37247
rect 23305 37213 23339 37247
rect 26525 37213 26559 37247
rect 27353 37213 27387 37247
rect 27813 37213 27847 37247
rect 28549 37213 28583 37247
rect 32597 37213 32631 37247
rect 33609 37213 33643 37247
rect 34897 37213 34931 37247
rect 36277 37213 36311 37247
rect 37565 37213 37599 37247
rect 25237 37145 25271 37179
rect 25329 37145 25363 37179
rect 30389 37145 30423 37179
rect 30481 37145 30515 37179
rect 2697 37077 2731 37111
rect 4169 37077 4203 37111
rect 4721 37077 4755 37111
rect 6745 37077 6779 37111
rect 8033 37077 8067 37111
rect 9505 37077 9539 37111
rect 10057 37077 10091 37111
rect 11069 37077 11103 37111
rect 14289 37077 14323 37111
rect 14933 37077 14967 37111
rect 15761 37077 15795 37111
rect 16865 37077 16899 37111
rect 17693 37077 17727 37111
rect 18797 37077 18831 37111
rect 20269 37077 20303 37111
rect 20821 37077 20855 37111
rect 23397 37077 23431 37111
rect 27169 37077 27203 37111
rect 27997 37077 28031 37111
rect 28641 37077 28675 37111
rect 33793 37077 33827 37111
rect 35081 37077 35115 37111
rect 36369 37077 36403 37111
rect 37657 37077 37691 37111
rect 20177 36873 20211 36907
rect 20821 36873 20855 36907
rect 22017 36873 22051 36907
rect 22661 36873 22695 36907
rect 27169 36873 27203 36907
rect 33241 36873 33275 36907
rect 24225 36805 24259 36839
rect 30389 36805 30423 36839
rect 38117 36805 38151 36839
rect 1777 36737 1811 36771
rect 2605 36737 2639 36771
rect 4721 36737 4755 36771
rect 7021 36737 7055 36771
rect 7665 36737 7699 36771
rect 10517 36737 10551 36771
rect 14933 36737 14967 36771
rect 16313 36737 16347 36771
rect 19441 36737 19475 36771
rect 20085 36737 20119 36771
rect 20729 36737 20763 36771
rect 22201 36737 22235 36771
rect 22845 36737 22879 36771
rect 23305 36737 23339 36771
rect 25881 36737 25915 36771
rect 26341 36737 26375 36771
rect 27353 36737 27387 36771
rect 32413 36737 32447 36771
rect 33057 36737 33091 36771
rect 35725 36737 35759 36771
rect 36921 36737 36955 36771
rect 7113 36669 7147 36703
rect 8493 36669 8527 36703
rect 8677 36669 8711 36703
rect 9689 36669 9723 36703
rect 12725 36669 12759 36703
rect 13001 36669 13035 36703
rect 16865 36669 16899 36703
rect 17141 36669 17175 36703
rect 19533 36669 19567 36703
rect 23397 36669 23431 36703
rect 24041 36669 24075 36703
rect 27905 36669 27939 36703
rect 28089 36669 28123 36703
rect 29009 36669 29043 36703
rect 30297 36669 30331 36703
rect 30573 36669 30607 36703
rect 14473 36601 14507 36635
rect 35541 36601 35575 36635
rect 1593 36533 1627 36567
rect 2697 36533 2731 36567
rect 4813 36533 4847 36567
rect 7757 36533 7791 36567
rect 9137 36533 9171 36567
rect 10333 36533 10367 36567
rect 15025 36533 15059 36567
rect 16129 36533 16163 36567
rect 18613 36533 18647 36567
rect 26433 36533 26467 36567
rect 32505 36533 32539 36567
rect 36737 36533 36771 36567
rect 38209 36533 38243 36567
rect 2237 36329 2271 36363
rect 8493 36329 8527 36363
rect 13645 36329 13679 36363
rect 37473 36329 37507 36363
rect 1593 36261 1627 36295
rect 10793 36261 10827 36295
rect 26985 36261 27019 36295
rect 31677 36261 31711 36295
rect 6469 36193 6503 36227
rect 9781 36193 9815 36227
rect 10425 36193 10459 36227
rect 20453 36193 20487 36227
rect 22201 36193 22235 36227
rect 28365 36193 28399 36227
rect 30205 36193 30239 36227
rect 32413 36193 32447 36227
rect 1777 36125 1811 36159
rect 2421 36125 2455 36159
rect 8401 36125 8435 36159
rect 10609 36125 10643 36159
rect 11713 36125 11747 36159
rect 12909 36125 12943 36159
rect 13553 36125 13587 36159
rect 14565 36125 14599 36159
rect 16773 36125 16807 36159
rect 19717 36125 19751 36159
rect 23673 36125 23707 36159
rect 27169 36125 27203 36159
rect 31861 36125 31895 36159
rect 32321 36125 32355 36159
rect 36829 36125 36863 36159
rect 37289 36125 37323 36159
rect 38025 36125 38059 36159
rect 6561 36057 6595 36091
rect 7481 36057 7515 36091
rect 9321 36057 9355 36091
rect 9413 36057 9447 36091
rect 14657 36057 14691 36091
rect 17049 36057 17083 36091
rect 20545 36057 20579 36091
rect 21097 36057 21131 36091
rect 22293 36057 22327 36091
rect 23213 36057 23247 36091
rect 24685 36057 24719 36091
rect 24777 36057 24811 36091
rect 25329 36057 25363 36091
rect 25881 36057 25915 36091
rect 25973 36057 26007 36091
rect 26525 36057 26559 36091
rect 28089 36057 28123 36091
rect 28181 36057 28215 36091
rect 30297 36057 30331 36091
rect 31217 36057 31251 36091
rect 11529 35989 11563 36023
rect 13001 35989 13035 36023
rect 18521 35989 18555 36023
rect 19809 35989 19843 36023
rect 23765 35989 23799 36023
rect 36645 35989 36679 36023
rect 38209 35989 38243 36023
rect 10885 35785 10919 35819
rect 20177 35785 20211 35819
rect 20821 35785 20855 35819
rect 23213 35785 23247 35819
rect 25605 35785 25639 35819
rect 26249 35785 26283 35819
rect 30941 35785 30975 35819
rect 9321 35717 9355 35751
rect 27997 35717 28031 35751
rect 29193 35717 29227 35751
rect 1685 35649 1719 35683
rect 2605 35649 2639 35683
rect 3433 35649 3467 35683
rect 9045 35649 9079 35683
rect 11069 35649 11103 35683
rect 19441 35649 19475 35683
rect 20085 35649 20119 35683
rect 20729 35649 20763 35683
rect 22201 35649 22235 35683
rect 23121 35649 23155 35683
rect 23765 35649 23799 35683
rect 24409 35649 24443 35683
rect 24593 35649 24627 35683
rect 25513 35649 25547 35683
rect 26157 35649 26191 35683
rect 27169 35649 27203 35683
rect 30389 35649 30423 35683
rect 30849 35649 30883 35683
rect 32505 35649 32539 35683
rect 12449 35581 12483 35615
rect 12725 35581 12759 35615
rect 16865 35581 16899 35615
rect 17141 35581 17175 35615
rect 22017 35581 22051 35615
rect 23857 35581 23891 35615
rect 27905 35581 27939 35615
rect 28181 35581 28215 35615
rect 29101 35581 29135 35615
rect 31493 35581 31527 35615
rect 37473 35581 37507 35615
rect 37749 35581 37783 35615
rect 18613 35513 18647 35547
rect 19533 35513 19567 35547
rect 22661 35513 22695 35547
rect 25053 35513 25087 35547
rect 29653 35513 29687 35547
rect 30205 35513 30239 35547
rect 1777 35445 1811 35479
rect 2697 35445 2731 35479
rect 3525 35445 3559 35479
rect 14197 35445 14231 35479
rect 27261 35445 27295 35479
rect 32321 35445 32355 35479
rect 3341 35241 3375 35275
rect 4077 35241 4111 35275
rect 10333 35241 10367 35275
rect 11240 35241 11274 35275
rect 12725 35241 12759 35275
rect 23765 35241 23799 35275
rect 30481 35241 30515 35275
rect 31033 35241 31067 35275
rect 16405 35173 16439 35207
rect 1869 35105 1903 35139
rect 6285 35105 6319 35139
rect 10977 35105 11011 35139
rect 13369 35105 13403 35139
rect 14657 35105 14691 35139
rect 14933 35105 14967 35139
rect 17141 35105 17175 35139
rect 24685 35105 24719 35139
rect 26249 35105 26283 35139
rect 27813 35105 27847 35139
rect 28181 35105 28215 35139
rect 1593 35037 1627 35071
rect 3985 35037 4019 35071
rect 6009 35037 6043 35071
rect 10517 35037 10551 35071
rect 13277 35037 13311 35071
rect 16865 35037 16899 35071
rect 19441 35037 19475 35071
rect 20177 35037 20211 35071
rect 20821 35037 20855 35071
rect 21465 35037 21499 35071
rect 22133 35037 22167 35071
rect 22753 35037 22787 35071
rect 23673 35037 23707 35071
rect 24593 35037 24627 35071
rect 25237 35037 25271 35071
rect 28917 35037 28951 35071
rect 29929 35037 29963 35071
rect 30389 35037 30423 35071
rect 31217 35037 31251 35071
rect 37841 35037 37875 35071
rect 26341 34969 26375 35003
rect 27261 34969 27295 35003
rect 27905 34969 27939 35003
rect 7757 34901 7791 34935
rect 18613 34901 18647 34935
rect 19533 34901 19567 34935
rect 20269 34901 20303 34935
rect 20913 34901 20947 34935
rect 21557 34901 21591 34935
rect 22201 34901 22235 34935
rect 22845 34901 22879 34935
rect 25329 34901 25363 34935
rect 29009 34901 29043 34935
rect 29745 34901 29779 34935
rect 38025 34901 38059 34935
rect 1593 34697 1627 34731
rect 5365 34697 5399 34731
rect 6653 34697 6687 34731
rect 11713 34697 11747 34731
rect 15577 34697 15611 34731
rect 28549 34697 28583 34731
rect 29837 34697 29871 34731
rect 30481 34697 30515 34731
rect 20913 34629 20947 34663
rect 22477 34629 22511 34663
rect 25697 34629 25731 34663
rect 27905 34629 27939 34663
rect 1777 34561 1811 34595
rect 2237 34561 2271 34595
rect 2329 34561 2363 34595
rect 6561 34561 6595 34595
rect 8125 34561 8159 34595
rect 11897 34561 11931 34595
rect 12633 34561 12667 34595
rect 12725 34561 12759 34595
rect 22385 34561 22419 34595
rect 23029 34561 23063 34595
rect 23673 34561 23707 34595
rect 24317 34561 24351 34595
rect 24961 34561 24995 34595
rect 25605 34561 25639 34595
rect 26249 34561 26283 34595
rect 27169 34561 27203 34595
rect 27813 34561 27847 34595
rect 28457 34561 28491 34595
rect 29101 34561 29135 34595
rect 29745 34561 29779 34595
rect 30389 34561 30423 34595
rect 38025 34561 38059 34595
rect 3617 34493 3651 34527
rect 3893 34493 3927 34527
rect 8217 34493 8251 34527
rect 13829 34493 13863 34527
rect 14105 34493 14139 34527
rect 16865 34493 16899 34527
rect 18613 34493 18647 34527
rect 20821 34493 20855 34527
rect 21189 34493 21223 34527
rect 23121 34493 23155 34527
rect 23765 34493 23799 34527
rect 25053 34493 25087 34527
rect 26341 34493 26375 34527
rect 29193 34493 29227 34527
rect 17128 34357 17162 34391
rect 24409 34357 24443 34391
rect 27261 34357 27295 34391
rect 38209 34357 38243 34391
rect 4077 34153 4111 34187
rect 8493 34153 8527 34187
rect 22201 34153 22235 34187
rect 29009 34153 29043 34187
rect 37841 34153 37875 34187
rect 23581 34085 23615 34119
rect 28365 34085 28399 34119
rect 6745 34017 6779 34051
rect 11069 34017 11103 34051
rect 11989 34017 12023 34051
rect 13737 34017 13771 34051
rect 15025 34017 15059 34051
rect 15945 34017 15979 34051
rect 23213 34017 23247 34051
rect 24685 34017 24719 34051
rect 24961 34017 24995 34051
rect 27813 34017 27847 34051
rect 3985 33949 4019 33983
rect 14289 33949 14323 33983
rect 22109 33949 22143 33983
rect 23397 33949 23431 33983
rect 25789 33949 25823 33983
rect 27261 33949 27295 33983
rect 28917 33949 28951 33983
rect 30389 33949 30423 33983
rect 38025 33949 38059 33983
rect 7021 33881 7055 33915
rect 10517 33881 10551 33915
rect 10609 33881 10643 33915
rect 12265 33881 12299 33915
rect 16221 33881 16255 33915
rect 24777 33881 24811 33915
rect 26617 33881 26651 33915
rect 26709 33881 26743 33915
rect 27905 33881 27939 33915
rect 17693 33813 17727 33847
rect 25881 33813 25915 33847
rect 29745 33813 29779 33847
rect 30481 33813 30515 33847
rect 11805 33609 11839 33643
rect 14933 33609 14967 33643
rect 21097 33609 21131 33643
rect 23489 33609 23523 33643
rect 26433 33609 26467 33643
rect 7757 33541 7791 33575
rect 17233 33541 17267 33575
rect 25053 33541 25087 33575
rect 28917 33541 28951 33575
rect 29009 33541 29043 33575
rect 1593 33473 1627 33507
rect 2513 33473 2547 33507
rect 4997 33473 5031 33507
rect 11713 33473 11747 33507
rect 13185 33473 13219 33507
rect 21005 33473 21039 33507
rect 22017 33473 22051 33507
rect 22661 33473 22695 33507
rect 23397 33473 23431 33507
rect 24041 33473 24075 33507
rect 26617 33473 26651 33507
rect 27169 33473 27203 33507
rect 27813 33473 27847 33507
rect 2789 33405 2823 33439
rect 5641 33405 5675 33439
rect 7481 33405 7515 33439
rect 9505 33405 9539 33439
rect 13461 33405 13495 33439
rect 16957 33405 16991 33439
rect 24962 33393 24996 33427
rect 25973 33405 26007 33439
rect 29193 33405 29227 33439
rect 1777 33337 1811 33371
rect 22109 33337 22143 33371
rect 27261 33337 27295 33371
rect 4261 33269 4295 33303
rect 5089 33269 5123 33303
rect 18705 33269 18739 33303
rect 22753 33269 22787 33303
rect 24133 33269 24167 33303
rect 27905 33269 27939 33303
rect 1856 33065 1890 33099
rect 4537 33065 4571 33099
rect 14381 33065 14415 33099
rect 20453 33065 20487 33099
rect 23949 33065 23983 33099
rect 1593 32929 1627 32963
rect 5549 32929 5583 32963
rect 9965 32929 9999 32963
rect 23305 32929 23339 32963
rect 24685 32929 24719 32963
rect 25145 32929 25179 32963
rect 26801 32929 26835 32963
rect 27721 32929 27755 32963
rect 4721 32861 4755 32895
rect 6193 32861 6227 32895
rect 6837 32861 6871 32895
rect 7297 32861 7331 32895
rect 9689 32861 9723 32895
rect 11713 32861 11747 32895
rect 14289 32861 14323 32895
rect 16865 32861 16899 32895
rect 18889 32861 18923 32895
rect 20361 32861 20395 32895
rect 22569 32861 22603 32895
rect 23213 32861 23247 32895
rect 23857 32861 23891 32895
rect 28825 32861 28859 32895
rect 5641 32793 5675 32827
rect 15209 32793 15243 32827
rect 15945 32793 15979 32827
rect 17141 32793 17175 32827
rect 21097 32793 21131 32827
rect 21189 32793 21223 32827
rect 22109 32793 22143 32827
rect 22661 32793 22695 32827
rect 24777 32793 24811 32827
rect 26157 32793 26191 32827
rect 26249 32793 26283 32827
rect 27813 32793 27847 32827
rect 28365 32793 28399 32827
rect 38117 32793 38151 32827
rect 3341 32725 3375 32759
rect 6653 32725 6687 32759
rect 7389 32725 7423 32759
rect 28917 32725 28951 32759
rect 38209 32725 38243 32759
rect 5733 32521 5767 32555
rect 26341 32521 26375 32555
rect 27261 32521 27295 32555
rect 27905 32521 27939 32555
rect 38117 32521 38151 32555
rect 7481 32453 7515 32487
rect 13553 32453 13587 32487
rect 15301 32453 15335 32487
rect 17141 32453 17175 32487
rect 23305 32453 23339 32487
rect 24862 32453 24896 32487
rect 1593 32385 1627 32419
rect 2329 32385 2363 32419
rect 5641 32385 5675 32419
rect 6653 32385 6687 32419
rect 8953 32385 8987 32419
rect 13277 32385 13311 32419
rect 16865 32385 16899 32419
rect 19717 32385 19751 32419
rect 20361 32385 20395 32419
rect 21005 32385 21039 32419
rect 22017 32385 22051 32419
rect 26249 32385 26283 32419
rect 27169 32385 27203 32419
rect 27813 32385 27847 32419
rect 38301 32385 38335 32419
rect 9229 32317 9263 32351
rect 19809 32317 19843 32351
rect 23213 32317 23247 32351
rect 24225 32317 24259 32351
rect 24777 32317 24811 32351
rect 25053 32317 25087 32351
rect 18613 32249 18647 32283
rect 1777 32181 1811 32215
rect 2421 32181 2455 32215
rect 10701 32181 10735 32215
rect 20453 32181 20487 32215
rect 21097 32181 21131 32215
rect 22109 32181 22143 32215
rect 2973 31977 3007 32011
rect 4077 31977 4111 32011
rect 7573 31977 7607 32011
rect 12068 31977 12102 32011
rect 24685 31977 24719 32011
rect 25973 31909 26007 31943
rect 5089 31841 5123 31875
rect 13553 31841 13587 31875
rect 16773 31841 16807 31875
rect 18521 31841 18555 31875
rect 20729 31841 20763 31875
rect 21741 31841 21775 31875
rect 22477 31841 22511 31875
rect 23121 31841 23155 31875
rect 26801 31841 26835 31875
rect 27445 31841 27479 31875
rect 28917 31841 28951 31875
rect 1869 31773 1903 31807
rect 1961 31773 1995 31807
rect 3157 31773 3191 31807
rect 3985 31773 4019 31807
rect 7113 31773 7147 31807
rect 7757 31773 7791 31807
rect 11805 31773 11839 31807
rect 24593 31773 24627 31807
rect 25237 31773 25271 31807
rect 25329 31773 25363 31807
rect 25881 31773 25915 31807
rect 5365 31705 5399 31739
rect 10333 31705 10367 31739
rect 11161 31705 11195 31739
rect 17049 31705 17083 31739
rect 20821 31705 20855 31739
rect 22569 31705 22603 31739
rect 26893 31705 26927 31739
rect 27997 31705 28031 31739
rect 28089 31705 28123 31739
rect 1593 31433 1627 31467
rect 6745 31433 6779 31467
rect 23213 31433 23247 31467
rect 27261 31433 27295 31467
rect 27813 31433 27847 31467
rect 12357 31365 12391 31399
rect 16129 31365 16163 31399
rect 17141 31365 17175 31399
rect 21189 31365 21223 31399
rect 25697 31365 25731 31399
rect 30021 31365 30055 31399
rect 1777 31297 1811 31331
rect 3341 31297 3375 31331
rect 3985 31297 4019 31331
rect 6929 31297 6963 31331
rect 8125 31297 8159 31331
rect 12081 31297 12115 31331
rect 15393 31297 15427 31331
rect 16865 31297 16899 31331
rect 20453 31297 20487 31331
rect 21097 31297 21131 31331
rect 22753 31297 22787 31331
rect 23673 31297 23707 31331
rect 24317 31297 24351 31331
rect 25145 31297 25179 31331
rect 25605 31297 25639 31331
rect 26433 31297 26467 31331
rect 27169 31297 27203 31331
rect 27997 31297 28031 31331
rect 29101 31297 29135 31331
rect 29929 31297 29963 31331
rect 4261 31229 4295 31263
rect 6009 31229 6043 31263
rect 8401 31229 8435 31263
rect 14105 31229 14139 31263
rect 20545 31229 20579 31263
rect 22569 31229 22603 31263
rect 28457 31229 28491 31263
rect 24409 31161 24443 31195
rect 26249 31161 26283 31195
rect 3433 31093 3467 31127
rect 9873 31093 9907 31127
rect 18613 31093 18647 31127
rect 23765 31093 23799 31127
rect 24961 31093 24995 31127
rect 29193 31093 29227 31127
rect 16037 30889 16071 30923
rect 30389 30821 30423 30855
rect 34897 30821 34931 30855
rect 14289 30753 14323 30787
rect 14565 30753 14599 30787
rect 20453 30753 20487 30787
rect 25789 30753 25823 30787
rect 37749 30753 37783 30787
rect 19717 30685 19751 30719
rect 21557 30685 21591 30719
rect 22753 30685 22787 30719
rect 23673 30685 23707 30719
rect 24593 30685 24627 30719
rect 26617 30685 26651 30719
rect 27261 30685 27295 30719
rect 27905 30685 27939 30719
rect 28549 30685 28583 30719
rect 35081 30685 35115 30719
rect 37473 30685 37507 30719
rect 20545 30617 20579 30651
rect 21097 30617 21131 30651
rect 21833 30617 21867 30651
rect 23029 30617 23063 30651
rect 25513 30617 25547 30651
rect 25605 30617 25639 30651
rect 29837 30617 29871 30651
rect 29929 30617 29963 30651
rect 19809 30549 19843 30583
rect 23765 30549 23799 30583
rect 24685 30549 24719 30583
rect 26709 30549 26743 30583
rect 27353 30549 27387 30583
rect 27997 30549 28031 30583
rect 28641 30549 28675 30583
rect 19809 30345 19843 30379
rect 17233 30277 17267 30311
rect 22201 30277 22235 30311
rect 23765 30277 23799 30311
rect 24685 30277 24719 30311
rect 26065 30277 26099 30311
rect 28825 30277 28859 30311
rect 2053 30209 2087 30243
rect 16957 30209 16991 30243
rect 19717 30209 19751 30243
rect 20821 30209 20855 30243
rect 25145 30209 25179 30243
rect 25237 30209 25271 30243
rect 27629 30209 27663 30243
rect 28733 30209 28767 30243
rect 29377 30209 29411 30243
rect 11713 30141 11747 30175
rect 11989 30141 12023 30175
rect 22109 30141 22143 30175
rect 22385 30141 22419 30175
rect 23673 30141 23707 30175
rect 25973 30141 26007 30175
rect 27813 30141 27847 30175
rect 13461 30073 13495 30107
rect 26525 30073 26559 30107
rect 29469 30073 29503 30107
rect 2145 30005 2179 30039
rect 18705 30005 18739 30039
rect 20913 30005 20947 30039
rect 27997 30005 28031 30039
rect 18153 29801 18187 29835
rect 13369 29733 13403 29767
rect 26617 29733 26651 29767
rect 16405 29665 16439 29699
rect 21649 29665 21683 29699
rect 27629 29665 27663 29699
rect 1777 29597 1811 29631
rect 11621 29597 11655 29631
rect 18705 29597 18739 29631
rect 18797 29597 18831 29631
rect 19533 29597 19567 29631
rect 20269 29597 20303 29631
rect 20913 29597 20947 29631
rect 23121 29597 23155 29631
rect 23765 29597 23799 29631
rect 26433 29597 26467 29631
rect 38025 29597 38059 29631
rect 11897 29529 11931 29563
rect 16681 29529 16715 29563
rect 19625 29529 19659 29563
rect 21741 29529 21775 29563
rect 22661 29529 22695 29563
rect 24685 29529 24719 29563
rect 24777 29529 24811 29563
rect 25697 29529 25731 29563
rect 27721 29529 27755 29563
rect 28641 29529 28675 29563
rect 1593 29461 1627 29495
rect 20361 29461 20395 29495
rect 21005 29461 21039 29495
rect 23213 29461 23247 29495
rect 23857 29461 23891 29495
rect 38209 29461 38243 29495
rect 8309 29257 8343 29291
rect 8953 29257 8987 29291
rect 27813 29257 27847 29291
rect 10241 29189 10275 29223
rect 17141 29189 17175 29223
rect 20729 29189 20763 29223
rect 23581 29189 23615 29223
rect 23673 29189 23707 29223
rect 25789 29189 25823 29223
rect 26341 29189 26375 29223
rect 1777 29121 1811 29155
rect 3249 29121 3283 29155
rect 8861 29121 8895 29155
rect 9505 29121 9539 29155
rect 14289 29121 14323 29155
rect 22017 29121 22051 29155
rect 22293 29121 22327 29155
rect 27353 29121 27387 29155
rect 28273 29121 28307 29155
rect 30573 29121 30607 29155
rect 6561 29053 6595 29087
rect 11069 29053 11103 29087
rect 11713 29053 11747 29087
rect 13737 29053 13771 29087
rect 16865 29053 16899 29087
rect 18613 29053 18647 29087
rect 20637 29053 20671 29087
rect 23857 29053 23891 29087
rect 25697 29053 25731 29087
rect 27169 29053 27203 29087
rect 28457 29053 28491 29087
rect 3341 28985 3375 29019
rect 9597 28985 9631 29019
rect 16037 28985 16071 29019
rect 21189 28985 21223 29019
rect 1593 28917 1627 28951
rect 6824 28917 6858 28951
rect 11976 28917 12010 28951
rect 14552 28917 14586 28951
rect 28641 28917 28675 28951
rect 30665 28917 30699 28951
rect 14289 28713 14323 28747
rect 28181 28713 28215 28747
rect 26433 28645 26467 28679
rect 21649 28577 21683 28611
rect 23029 28577 23063 28611
rect 25881 28577 25915 28611
rect 27721 28577 27755 28611
rect 28733 28577 28767 28611
rect 1869 28509 1903 28543
rect 2789 28509 2823 28543
rect 6929 28509 6963 28543
rect 11253 28509 11287 28543
rect 13553 28509 13587 28543
rect 14473 28509 14507 28543
rect 15198 28509 15232 28543
rect 18245 28509 18279 28543
rect 19993 28509 20027 28543
rect 20637 28509 20671 28543
rect 21557 28509 21591 28543
rect 22201 28509 22235 28543
rect 24593 28509 24627 28543
rect 27537 28509 27571 28543
rect 28641 28509 28675 28543
rect 29745 28509 29779 28543
rect 31493 28509 31527 28543
rect 1961 28441 1995 28475
rect 6193 28441 6227 28475
rect 11529 28441 11563 28475
rect 15485 28441 15519 28475
rect 17509 28441 17543 28475
rect 20913 28441 20947 28475
rect 23121 28441 23155 28475
rect 24041 28441 24075 28475
rect 25973 28441 26007 28475
rect 29837 28441 29871 28475
rect 2881 28373 2915 28407
rect 13001 28373 13035 28407
rect 13645 28373 13679 28407
rect 16957 28373 16991 28407
rect 20085 28373 20119 28407
rect 22293 28373 22327 28407
rect 24685 28373 24719 28407
rect 31309 28373 31343 28407
rect 29009 28169 29043 28203
rect 6009 28101 6043 28135
rect 21005 28101 21039 28135
rect 22201 28101 22235 28135
rect 23765 28101 23799 28135
rect 24317 28101 24351 28135
rect 25697 28101 25731 28135
rect 26617 28101 26651 28135
rect 27353 28101 27387 28135
rect 27905 28101 27939 28135
rect 1777 28033 1811 28067
rect 8217 28033 8251 28067
rect 12817 28033 12851 28067
rect 19073 28033 19107 28067
rect 19165 28033 19199 28067
rect 20913 28033 20947 28067
rect 24777 28033 24811 28067
rect 28365 28033 28399 28067
rect 29193 28033 29227 28067
rect 38025 28033 38059 28067
rect 3985 27965 4019 27999
rect 4261 27965 4295 27999
rect 8493 27965 8527 27999
rect 13093 27965 13127 27999
rect 16865 27965 16899 27999
rect 17141 27965 17175 27999
rect 22109 27965 22143 27999
rect 23121 27965 23155 27999
rect 23673 27965 23707 27999
rect 25605 27965 25639 27999
rect 27261 27965 27295 27999
rect 24869 27897 24903 27931
rect 38209 27897 38243 27931
rect 1593 27829 1627 27863
rect 9965 27829 9999 27863
rect 14565 27829 14599 27863
rect 18613 27829 18647 27863
rect 28457 27829 28491 27863
rect 1850 27625 1884 27659
rect 27169 27625 27203 27659
rect 3341 27557 3375 27591
rect 24685 27557 24719 27591
rect 25973 27557 26007 27591
rect 28457 27557 28491 27591
rect 32413 27557 32447 27591
rect 1593 27489 1627 27523
rect 15853 27489 15887 27523
rect 16116 27489 16150 27523
rect 21925 27489 21959 27523
rect 4445 27421 4479 27455
rect 18337 27421 18371 27455
rect 19533 27421 19567 27455
rect 23397 27421 23431 27455
rect 24593 27421 24627 27455
rect 25237 27421 25271 27455
rect 25329 27421 25363 27455
rect 25881 27421 25915 27455
rect 26525 27421 26559 27455
rect 27353 27421 27387 27455
rect 27813 27421 27847 27455
rect 28641 27421 28675 27455
rect 29745 27421 29779 27455
rect 30389 27421 30423 27455
rect 32597 27421 32631 27455
rect 38025 27421 38059 27455
rect 10241 27353 10275 27387
rect 17877 27353 17911 27387
rect 18429 27353 18463 27387
rect 19717 27353 19751 27387
rect 21373 27353 21407 27387
rect 22017 27353 22051 27387
rect 22937 27353 22971 27387
rect 4537 27285 4571 27319
rect 11529 27285 11563 27319
rect 23489 27285 23523 27319
rect 26617 27285 26651 27319
rect 27905 27285 27939 27319
rect 29837 27285 29871 27319
rect 30481 27285 30515 27319
rect 38209 27285 38243 27319
rect 20085 27081 20119 27115
rect 31585 27081 31619 27115
rect 37841 27081 37875 27115
rect 3709 27013 3743 27047
rect 13737 27013 13771 27047
rect 17141 27013 17175 27047
rect 22201 27013 22235 27047
rect 24501 27013 24535 27047
rect 27353 27013 27387 27047
rect 1685 26945 1719 26979
rect 11713 26945 11747 26979
rect 14197 26945 14231 26979
rect 16865 26945 16899 26979
rect 19073 26945 19107 26979
rect 19993 26945 20027 26979
rect 25881 26945 25915 26979
rect 31493 26945 31527 26979
rect 38025 26945 38059 26979
rect 3433 26877 3467 26911
rect 11989 26877 12023 26911
rect 19349 26877 19383 26911
rect 22017 26877 22051 26911
rect 23857 26877 23891 26911
rect 24409 26877 24443 26911
rect 25421 26877 25455 26911
rect 27261 26877 27295 26911
rect 28181 26877 28215 26911
rect 1869 26809 1903 26843
rect 5181 26741 5215 26775
rect 14289 26741 14323 26775
rect 18613 26741 18647 26775
rect 25973 26741 26007 26775
rect 21097 26537 21131 26571
rect 24685 26537 24719 26571
rect 26893 26537 26927 26571
rect 29193 26537 29227 26571
rect 38117 26537 38151 26571
rect 11989 26469 12023 26503
rect 19533 26469 19567 26503
rect 29745 26469 29779 26503
rect 2421 26401 2455 26435
rect 8033 26401 8067 26435
rect 10241 26401 10275 26435
rect 16589 26401 16623 26435
rect 26433 26401 26467 26435
rect 6285 26333 6319 26367
rect 19433 26333 19467 26367
rect 20361 26333 20395 26367
rect 21005 26333 21039 26367
rect 21649 26333 21683 26367
rect 22661 26333 22695 26367
rect 23305 26333 23339 26367
rect 23397 26333 23431 26367
rect 24593 26333 24627 26367
rect 25237 26333 25271 26367
rect 26249 26333 26283 26367
rect 28549 26333 28583 26367
rect 28733 26333 28767 26367
rect 29929 26333 29963 26367
rect 38301 26333 38335 26367
rect 2513 26265 2547 26299
rect 3433 26265 3467 26299
rect 6561 26265 6595 26299
rect 10517 26265 10551 26299
rect 16865 26265 16899 26299
rect 18613 26265 18647 26299
rect 20453 26265 20487 26299
rect 21741 26265 21775 26299
rect 22753 26265 22787 26299
rect 25329 26197 25363 26231
rect 10793 25993 10827 26027
rect 19165 25993 19199 26027
rect 28733 25993 28767 26027
rect 24777 25925 24811 25959
rect 25697 25925 25731 25959
rect 29929 25925 29963 25959
rect 3525 25857 3559 25891
rect 12265 25857 12299 25891
rect 19073 25857 19107 25891
rect 19717 25857 19751 25891
rect 22293 25857 22327 25891
rect 26157 25857 26191 25891
rect 4169 25789 4203 25823
rect 4445 25789 4479 25823
rect 9045 25789 9079 25823
rect 9321 25789 9355 25823
rect 12541 25789 12575 25823
rect 14289 25789 14323 25823
rect 16865 25789 16899 25823
rect 17141 25789 17175 25823
rect 22477 25789 22511 25823
rect 24133 25789 24167 25823
rect 24685 25789 24719 25823
rect 29837 25789 29871 25823
rect 30849 25789 30883 25823
rect 3617 25653 3651 25687
rect 5917 25653 5951 25687
rect 18613 25653 18647 25687
rect 19809 25653 19843 25687
rect 26249 25653 26283 25687
rect 15012 25449 15046 25483
rect 22385 25449 22419 25483
rect 28825 25449 28859 25483
rect 26525 25381 26559 25415
rect 6101 25313 6135 25347
rect 20178 25313 20212 25347
rect 29929 25313 29963 25347
rect 1593 25245 1627 25279
rect 4905 25245 4939 25279
rect 14749 25245 14783 25279
rect 18061 25245 18095 25279
rect 19441 25245 19475 25279
rect 21649 25245 21683 25279
rect 22293 25245 22327 25279
rect 22937 25245 22971 25279
rect 23581 25245 23615 25279
rect 25329 25245 25363 25279
rect 25789 25245 25823 25279
rect 26433 25245 26467 25279
rect 27077 25245 27111 25279
rect 28365 25245 28399 25279
rect 29009 25245 29043 25279
rect 31493 25245 31527 25279
rect 4169 25177 4203 25211
rect 6377 25177 6411 25211
rect 18153 25177 18187 25211
rect 20269 25177 20303 25211
rect 21189 25177 21223 25211
rect 23673 25177 23707 25211
rect 24685 25177 24719 25211
rect 24777 25177 24811 25211
rect 1777 25109 1811 25143
rect 7849 25109 7883 25143
rect 16497 25109 16531 25143
rect 19533 25109 19567 25143
rect 21741 25109 21775 25143
rect 23029 25109 23063 25143
rect 25881 25109 25915 25143
rect 27169 25109 27203 25143
rect 28181 25109 28215 25143
rect 31585 25109 31619 25143
rect 5365 24905 5399 24939
rect 20453 24837 20487 24871
rect 24041 24837 24075 24871
rect 24961 24837 24995 24871
rect 1777 24769 1811 24803
rect 16865 24769 16899 24803
rect 18337 24769 18371 24803
rect 18981 24769 19015 24803
rect 19625 24769 19659 24803
rect 22201 24769 22235 24803
rect 22661 24769 22695 24803
rect 25513 24769 25547 24803
rect 25697 24769 25731 24803
rect 27353 24769 27387 24803
rect 27997 24769 28031 24803
rect 29009 24769 29043 24803
rect 38025 24769 38059 24803
rect 3617 24701 3651 24735
rect 3893 24701 3927 24735
rect 13277 24701 13311 24735
rect 13553 24701 13587 24735
rect 15025 24701 15059 24735
rect 17601 24701 17635 24735
rect 19073 24701 19107 24735
rect 20361 24701 20395 24735
rect 21189 24701 21223 24735
rect 23949 24701 23983 24735
rect 19717 24633 19751 24667
rect 22753 24633 22787 24667
rect 1593 24565 1627 24599
rect 18429 24565 18463 24599
rect 22017 24565 22051 24599
rect 25881 24565 25915 24599
rect 27169 24565 27203 24599
rect 28089 24565 28123 24599
rect 29101 24565 29135 24599
rect 38209 24565 38243 24599
rect 6837 24361 6871 24395
rect 26249 24361 26283 24395
rect 38117 24361 38151 24395
rect 2237 24293 2271 24327
rect 20085 24293 20119 24327
rect 21925 24293 21959 24327
rect 5089 24225 5123 24259
rect 5365 24225 5399 24259
rect 9873 24225 9907 24259
rect 12173 24225 12207 24259
rect 16497 24225 16531 24259
rect 1593 24157 1627 24191
rect 4445 24157 4479 24191
rect 18705 24157 18739 24191
rect 19993 24157 20027 24191
rect 21373 24157 21407 24191
rect 21833 24157 21867 24191
rect 22661 24157 22695 24191
rect 23121 24157 23155 24191
rect 23765 24157 23799 24191
rect 26157 24157 26191 24191
rect 26801 24157 26835 24191
rect 38301 24157 38335 24191
rect 9137 24089 9171 24123
rect 11345 24089 11379 24123
rect 16773 24089 16807 24123
rect 20729 24089 20763 24123
rect 20821 24089 20855 24123
rect 24685 24089 24719 24123
rect 24777 24089 24811 24123
rect 25697 24089 25731 24123
rect 1777 24021 1811 24055
rect 4537 24021 4571 24055
rect 18245 24021 18279 24055
rect 18797 24021 18831 24055
rect 22477 24021 22511 24055
rect 23213 24021 23247 24055
rect 23857 24021 23891 24055
rect 26893 24021 26927 24055
rect 1869 23817 1903 23851
rect 9229 23817 9263 23851
rect 15025 23817 15059 23851
rect 18613 23817 18647 23851
rect 25513 23817 25547 23851
rect 5365 23749 5399 23783
rect 20545 23749 20579 23783
rect 22569 23749 22603 23783
rect 1777 23681 1811 23715
rect 5273 23681 5307 23715
rect 6561 23681 6595 23715
rect 7481 23681 7515 23715
rect 12265 23681 12299 23715
rect 16865 23681 16899 23715
rect 23949 23681 23983 23715
rect 25053 23681 25087 23715
rect 25973 23681 26007 23715
rect 2421 23613 2455 23647
rect 2697 23613 2731 23647
rect 7757 23613 7791 23647
rect 13277 23613 13311 23647
rect 13553 23613 13587 23647
rect 17141 23613 17175 23647
rect 20442 23613 20476 23647
rect 21465 23613 21499 23647
rect 22477 23613 22511 23647
rect 22937 23613 22971 23647
rect 24869 23613 24903 23647
rect 31217 23613 31251 23647
rect 4169 23545 4203 23579
rect 6653 23477 6687 23511
rect 12357 23477 12391 23511
rect 24041 23477 24075 23511
rect 26065 23477 26099 23511
rect 21557 23273 21591 23307
rect 29837 23273 29871 23307
rect 25237 23205 25271 23239
rect 6653 23137 6687 23171
rect 10425 23137 10459 23171
rect 14565 23137 14599 23171
rect 18705 23137 18739 23171
rect 20545 23137 20579 23171
rect 31125 23137 31159 23171
rect 1869 23069 1903 23103
rect 5273 23069 5307 23103
rect 5917 23069 5951 23103
rect 7297 23069 7331 23103
rect 13093 23069 13127 23103
rect 14289 23069 14323 23103
rect 17969 23069 18003 23103
rect 20085 23069 20119 23103
rect 21465 23069 21499 23103
rect 25789 23069 25823 23103
rect 29745 23069 29779 23103
rect 38025 23069 38059 23103
rect 10701 23001 10735 23035
rect 13645 23001 13679 23035
rect 22661 23001 22695 23035
rect 22753 23001 22787 23035
rect 23673 23001 23707 23035
rect 24685 23001 24719 23035
rect 24777 23001 24811 23035
rect 31217 23001 31251 23035
rect 32137 23001 32171 23035
rect 1961 22933 1995 22967
rect 5365 22933 5399 22967
rect 7389 22933 7423 22967
rect 12173 22933 12207 22967
rect 16037 22933 16071 22967
rect 25881 22933 25915 22967
rect 26433 22933 26467 22967
rect 37841 22933 37875 22967
rect 36093 22729 36127 22763
rect 8033 22661 8067 22695
rect 12541 22661 12575 22695
rect 14289 22661 14323 22695
rect 24409 22661 24443 22695
rect 24961 22661 24995 22695
rect 25605 22661 25639 22695
rect 25697 22661 25731 22695
rect 27261 22661 27295 22695
rect 1777 22593 1811 22627
rect 7757 22593 7791 22627
rect 12265 22593 12299 22627
rect 18613 22593 18647 22627
rect 27169 22593 27203 22627
rect 36001 22593 36035 22627
rect 38025 22593 38059 22627
rect 2053 22525 2087 22559
rect 9505 22525 9539 22559
rect 24317 22525 24351 22559
rect 26617 22525 26651 22559
rect 38209 22457 38243 22491
rect 3525 22389 3559 22423
rect 18705 22389 18739 22423
rect 4242 22185 4276 22219
rect 7100 22185 7134 22219
rect 3985 22049 4019 22083
rect 5733 22049 5767 22083
rect 6837 22049 6871 22083
rect 25881 22049 25915 22083
rect 1593 21981 1627 22015
rect 10241 21981 10275 22015
rect 15117 21981 15151 22015
rect 19441 21981 19475 22015
rect 21833 21981 21867 22015
rect 27353 21981 27387 22015
rect 27997 21981 28031 22015
rect 29745 21981 29779 22015
rect 15393 21913 15427 21947
rect 25973 21913 26007 21947
rect 26893 21913 26927 21947
rect 1777 21845 1811 21879
rect 8585 21845 8619 21879
rect 10333 21845 10367 21879
rect 16865 21845 16899 21879
rect 19533 21845 19567 21879
rect 21925 21845 21959 21879
rect 27445 21845 27479 21879
rect 28089 21845 28123 21879
rect 29837 21845 29871 21879
rect 14197 21573 14231 21607
rect 17141 21573 17175 21607
rect 20085 21573 20119 21607
rect 27997 21573 28031 21607
rect 1777 21505 1811 21539
rect 3985 21505 4019 21539
rect 11989 21505 12023 21539
rect 14933 21505 14967 21539
rect 16865 21505 16899 21539
rect 19165 21505 19199 21539
rect 19993 21505 20027 21539
rect 20729 21505 20763 21539
rect 23397 21505 23431 21539
rect 26525 21505 26559 21539
rect 38301 21505 38335 21539
rect 4261 21437 4295 21471
rect 6009 21437 6043 21471
rect 6929 21437 6963 21471
rect 7205 21437 7239 21471
rect 9137 21437 9171 21471
rect 9413 21437 9447 21471
rect 11161 21437 11195 21471
rect 20821 21437 20855 21471
rect 27905 21437 27939 21471
rect 28181 21437 28215 21471
rect 23489 21369 23523 21403
rect 1593 21301 1627 21335
rect 8677 21301 8711 21335
rect 12246 21301 12280 21335
rect 13737 21301 13771 21335
rect 18613 21301 18647 21335
rect 19257 21301 19291 21335
rect 26341 21301 26375 21335
rect 38117 21301 38151 21335
rect 1856 21097 1890 21131
rect 9781 21097 9815 21131
rect 17693 21097 17727 21131
rect 8585 21029 8619 21063
rect 1593 20961 1627 20995
rect 4629 20961 4663 20995
rect 4905 20961 4939 20995
rect 11253 20961 11287 20995
rect 15945 20961 15979 20995
rect 16221 20961 16255 20995
rect 26985 20961 27019 20995
rect 28273 20961 28307 20995
rect 29837 20961 29871 20995
rect 6837 20893 6871 20927
rect 9689 20893 9723 20927
rect 10333 20893 10367 20927
rect 10977 20893 11011 20927
rect 23673 20893 23707 20927
rect 29745 20893 29779 20927
rect 30389 20893 30423 20927
rect 38301 20893 38335 20927
rect 7113 20825 7147 20859
rect 19809 20825 19843 20859
rect 19901 20825 19935 20859
rect 20821 20825 20855 20859
rect 26341 20825 26375 20859
rect 26433 20825 26467 20859
rect 28365 20825 28399 20859
rect 28917 20825 28951 20859
rect 3341 20757 3375 20791
rect 6377 20757 6411 20791
rect 10425 20757 10459 20791
rect 12725 20757 12759 20791
rect 23489 20757 23523 20791
rect 30481 20757 30515 20791
rect 1777 20553 1811 20587
rect 24777 20553 24811 20587
rect 7757 20485 7791 20519
rect 8493 20485 8527 20519
rect 11897 20485 11931 20519
rect 22937 20485 22971 20519
rect 23765 20485 23799 20519
rect 25789 20485 25823 20519
rect 28273 20485 28307 20519
rect 29653 20485 29687 20519
rect 1685 20417 1719 20451
rect 13369 20417 13403 20451
rect 16865 20417 16899 20451
rect 19073 20417 19107 20451
rect 22017 20417 22051 20451
rect 24961 20417 24995 20451
rect 28181 20417 28215 20451
rect 29009 20417 29043 20451
rect 2421 20349 2455 20383
rect 2697 20349 2731 20383
rect 9137 20349 9171 20383
rect 9413 20349 9447 20383
rect 12633 20349 12667 20383
rect 13645 20349 13679 20383
rect 23673 20349 23707 20383
rect 24041 20349 24075 20383
rect 25697 20349 25731 20383
rect 29561 20349 29595 20383
rect 30389 20349 30423 20383
rect 23121 20281 23155 20315
rect 26249 20281 26283 20315
rect 4169 20213 4203 20247
rect 10885 20213 10919 20247
rect 15117 20213 15151 20247
rect 16957 20213 16991 20247
rect 19165 20213 19199 20247
rect 22109 20213 22143 20247
rect 28825 20213 28859 20247
rect 10872 20009 10906 20043
rect 5733 19941 5767 19975
rect 12357 19941 12391 19975
rect 1685 19873 1719 19907
rect 3985 19873 4019 19907
rect 4261 19873 4295 19907
rect 6561 19873 6595 19907
rect 10609 19873 10643 19907
rect 16589 19873 16623 19907
rect 20545 19873 20579 19907
rect 20913 19873 20947 19907
rect 23765 19873 23799 19907
rect 26157 19873 26191 19907
rect 26617 19873 26651 19907
rect 6285 19805 6319 19839
rect 12909 19805 12943 19839
rect 20361 19805 20395 19839
rect 24961 19805 24995 19839
rect 28365 19805 28399 19839
rect 29009 19805 29043 19839
rect 1961 19737 1995 19771
rect 13185 19737 13219 19771
rect 16865 19737 16899 19771
rect 22753 19737 22787 19771
rect 22845 19737 22879 19771
rect 26249 19737 26283 19771
rect 27721 19737 27755 19771
rect 3433 19669 3467 19703
rect 8033 19669 8067 19703
rect 18337 19669 18371 19703
rect 25053 19669 25087 19703
rect 27813 19669 27847 19703
rect 28457 19669 28491 19703
rect 29101 19669 29135 19703
rect 3341 19465 3375 19499
rect 6009 19465 6043 19499
rect 15853 19465 15887 19499
rect 18613 19465 18647 19499
rect 20361 19465 20395 19499
rect 38117 19465 38151 19499
rect 21097 19397 21131 19431
rect 22201 19397 22235 19431
rect 23121 19397 23155 19431
rect 24225 19397 24259 19431
rect 29009 19397 29043 19431
rect 29929 19397 29963 19431
rect 30573 19397 30607 19431
rect 4261 19329 4295 19363
rect 8217 19329 8251 19363
rect 14105 19329 14139 19363
rect 16865 19329 16899 19363
rect 21005 19329 21039 19363
rect 23581 19329 23615 19363
rect 24869 19329 24903 19363
rect 38301 19329 38335 19363
rect 1593 19261 1627 19295
rect 1869 19261 1903 19295
rect 4537 19261 4571 19295
rect 8493 19261 8527 19295
rect 11897 19261 11931 19295
rect 12173 19261 12207 19295
rect 13645 19261 13679 19295
rect 14381 19261 14415 19295
rect 17141 19261 17175 19295
rect 22109 19261 22143 19295
rect 23765 19261 23799 19295
rect 28917 19261 28951 19295
rect 30481 19261 30515 19295
rect 30757 19261 30791 19295
rect 24685 19193 24719 19227
rect 9965 19125 9999 19159
rect 12817 18921 12851 18955
rect 19533 18921 19567 18955
rect 22753 18921 22787 18955
rect 30113 18921 30147 18955
rect 25237 18853 25271 18887
rect 1961 18785 1995 18819
rect 4629 18785 4663 18819
rect 7113 18785 7147 18819
rect 8585 18785 8619 18819
rect 11345 18785 11379 18819
rect 14749 18785 14783 18819
rect 23949 18785 23983 18819
rect 24685 18785 24719 18819
rect 25789 18785 25823 18819
rect 1685 18717 1719 18751
rect 6837 18717 6871 18751
rect 11069 18717 11103 18751
rect 16773 18717 16807 18751
rect 19441 18717 19475 18751
rect 22109 18717 22143 18751
rect 22293 18717 22327 18751
rect 23213 18717 23247 18751
rect 23857 18717 23891 18751
rect 30021 18717 30055 18751
rect 4905 18649 4939 18683
rect 15025 18649 15059 18683
rect 24777 18649 24811 18683
rect 3433 18581 3467 18615
rect 6377 18581 6411 18615
rect 23305 18581 23339 18615
rect 6009 18377 6043 18411
rect 6653 18377 6687 18411
rect 11805 18377 11839 18411
rect 15301 18377 15335 18411
rect 18613 18377 18647 18411
rect 22661 18377 22695 18411
rect 23121 18377 23155 18411
rect 38117 18377 38151 18411
rect 17141 18309 17175 18343
rect 2053 18241 2087 18275
rect 4261 18241 4295 18275
rect 6561 18241 6595 18275
rect 11713 18241 11747 18275
rect 13553 18241 13587 18275
rect 16865 18241 16899 18275
rect 19809 18241 19843 18275
rect 20545 18241 20579 18275
rect 22017 18241 22051 18275
rect 22201 18241 22235 18275
rect 23305 18241 23339 18275
rect 24501 18241 24535 18275
rect 38301 18241 38335 18275
rect 2329 18173 2363 18207
rect 4537 18173 4571 18207
rect 7297 18173 7331 18207
rect 7573 18173 7607 18207
rect 9321 18173 9355 18207
rect 13829 18173 13863 18207
rect 24685 18173 24719 18207
rect 3801 18037 3835 18071
rect 19901 18037 19935 18071
rect 20637 18037 20671 18071
rect 5733 17833 5767 17867
rect 11529 17833 11563 17867
rect 22569 17833 22603 17867
rect 3985 17697 4019 17731
rect 4261 17697 4295 17731
rect 6377 17697 6411 17731
rect 9781 17697 9815 17731
rect 10057 17697 10091 17731
rect 12265 17697 12299 17731
rect 16313 17697 16347 17731
rect 19809 17697 19843 17731
rect 20821 17697 20855 17731
rect 22109 17697 22143 17731
rect 1777 17629 1811 17663
rect 2237 17629 2271 17663
rect 11989 17629 12023 17663
rect 18521 17629 18555 17663
rect 19625 17629 19659 17663
rect 21925 17629 21959 17663
rect 6653 17561 6687 17595
rect 16589 17561 16623 17595
rect 18613 17561 18647 17595
rect 1593 17493 1627 17527
rect 2329 17493 2363 17527
rect 8125 17493 8159 17527
rect 13737 17493 13771 17527
rect 18061 17493 18095 17527
rect 2329 17289 2363 17323
rect 3157 17289 3191 17323
rect 14013 17289 14047 17323
rect 17785 17289 17819 17323
rect 18429 17289 18463 17323
rect 19717 17289 19751 17323
rect 20729 17289 20763 17323
rect 29193 17289 29227 17323
rect 4445 17221 4479 17255
rect 11897 17221 11931 17255
rect 1685 17153 1719 17187
rect 2513 17153 2547 17187
rect 3065 17153 3099 17187
rect 3709 17153 3743 17187
rect 4353 17153 4387 17187
rect 5457 17153 5491 17187
rect 9413 17153 9447 17187
rect 12633 17153 12667 17187
rect 13921 17153 13955 17187
rect 16037 17153 16071 17187
rect 17693 17153 17727 17187
rect 18337 17153 18371 17187
rect 18981 17153 19015 17187
rect 20637 17153 20671 17187
rect 29101 17153 29135 17187
rect 37841 17153 37875 17187
rect 9689 17085 9723 17119
rect 1869 17017 1903 17051
rect 3801 16949 3835 16983
rect 5549 16949 5583 16983
rect 11161 16949 11195 16983
rect 16129 16949 16163 16983
rect 19073 16949 19107 16983
rect 37657 16949 37691 16983
rect 23305 16609 23339 16643
rect 1961 16541 1995 16575
rect 2605 16541 2639 16575
rect 3249 16541 3283 16575
rect 4077 16541 4111 16575
rect 5181 16541 5215 16575
rect 5825 16541 5859 16575
rect 6469 16541 6503 16575
rect 6561 16541 6595 16575
rect 7297 16541 7331 16575
rect 8033 16541 8067 16575
rect 9873 16541 9907 16575
rect 10701 16541 10735 16575
rect 11621 16541 11655 16575
rect 13553 16541 13587 16575
rect 13645 16541 13679 16575
rect 14749 16541 14783 16575
rect 14841 16541 14875 16575
rect 15577 16541 15611 16575
rect 16681 16541 16715 16575
rect 21281 16541 21315 16575
rect 37565 16541 37599 16575
rect 2053 16473 2087 16507
rect 4169 16473 4203 16507
rect 17417 16473 17451 16507
rect 17509 16473 17543 16507
rect 18061 16473 18095 16507
rect 23029 16473 23063 16507
rect 23121 16473 23155 16507
rect 38117 16473 38151 16507
rect 2697 16405 2731 16439
rect 3341 16405 3375 16439
rect 5273 16405 5307 16439
rect 5917 16405 5951 16439
rect 7389 16405 7423 16439
rect 8125 16405 8159 16439
rect 9965 16405 9999 16439
rect 10793 16405 10827 16439
rect 11713 16405 11747 16439
rect 15393 16405 15427 16439
rect 16773 16405 16807 16439
rect 21373 16405 21407 16439
rect 37381 16405 37415 16439
rect 38209 16405 38243 16439
rect 3341 16201 3375 16235
rect 6929 16201 6963 16235
rect 8217 16201 8251 16235
rect 8861 16201 8895 16235
rect 10425 16201 10459 16235
rect 11069 16201 11103 16235
rect 13737 16201 13771 16235
rect 16129 16201 16163 16235
rect 38117 16201 38151 16235
rect 4169 16133 4203 16167
rect 4261 16133 4295 16167
rect 11897 16133 11931 16167
rect 12633 16133 12667 16167
rect 17049 16133 17083 16167
rect 19165 16133 19199 16167
rect 20545 16133 20579 16167
rect 22845 16133 22879 16167
rect 1593 16065 1627 16099
rect 2605 16065 2639 16099
rect 3249 16065 3283 16099
rect 5825 16065 5859 16099
rect 6837 16065 6871 16099
rect 8125 16065 8159 16099
rect 8769 16065 8803 16099
rect 9689 16065 9723 16099
rect 10333 16065 10367 16099
rect 10977 16065 11011 16099
rect 13645 16065 13679 16099
rect 16313 16065 16347 16099
rect 22017 16065 22051 16099
rect 27445 16065 27479 16099
rect 33517 16065 33551 16099
rect 38301 16065 38335 16099
rect 2697 15997 2731 16031
rect 5181 15997 5215 16031
rect 5917 15997 5951 16031
rect 16957 15997 16991 16031
rect 17969 15997 18003 16031
rect 19073 15997 19107 16031
rect 19349 15997 19383 16031
rect 20453 15997 20487 16031
rect 20729 15997 20763 16031
rect 22753 15997 22787 16031
rect 23581 15997 23615 16031
rect 26249 15997 26283 16031
rect 1777 15861 1811 15895
rect 9781 15861 9815 15895
rect 22109 15861 22143 15895
rect 27537 15861 27571 15895
rect 33333 15861 33367 15895
rect 6653 15657 6687 15691
rect 9413 15657 9447 15691
rect 3157 15589 3191 15623
rect 5917 15589 5951 15623
rect 30021 15589 30055 15623
rect 2789 15521 2823 15555
rect 10333 15521 10367 15555
rect 23489 15521 23523 15555
rect 26157 15521 26191 15555
rect 26341 15521 26375 15555
rect 27905 15521 27939 15555
rect 1593 15453 1627 15487
rect 2973 15453 3007 15487
rect 5825 15453 5859 15487
rect 6561 15453 6595 15487
rect 9321 15453 9355 15487
rect 12909 15453 12943 15487
rect 13185 15453 13219 15487
rect 18705 15453 18739 15487
rect 19441 15453 19475 15487
rect 21097 15453 21131 15487
rect 21189 15453 21223 15487
rect 4353 15385 4387 15419
rect 4445 15385 4479 15419
rect 5365 15385 5399 15419
rect 7573 15385 7607 15419
rect 7665 15385 7699 15419
rect 8585 15385 8619 15419
rect 10057 15385 10091 15419
rect 10149 15385 10183 15419
rect 11437 15385 11471 15419
rect 11529 15385 11563 15419
rect 12449 15385 12483 15419
rect 16865 15385 16899 15419
rect 16957 15385 16991 15419
rect 17877 15385 17911 15419
rect 22845 15385 22879 15419
rect 22937 15385 22971 15419
rect 24685 15385 24719 15419
rect 24777 15385 24811 15419
rect 25697 15385 25731 15419
rect 29837 15385 29871 15419
rect 1777 15317 1811 15351
rect 18797 15317 18831 15351
rect 19533 15317 19567 15351
rect 12449 15113 12483 15147
rect 2053 15045 2087 15079
rect 6745 15045 6779 15079
rect 10241 15045 10275 15079
rect 11161 15045 11195 15079
rect 17049 15045 17083 15079
rect 22201 15045 22235 15079
rect 23121 15045 23155 15079
rect 23857 15045 23891 15079
rect 7297 14977 7331 15011
rect 7757 14977 7791 15011
rect 9137 14977 9171 15011
rect 11713 14977 11747 15011
rect 12357 14977 12391 15011
rect 18429 14977 18463 15011
rect 19073 14977 19107 15011
rect 21281 14977 21315 15011
rect 1869 14909 1903 14943
rect 3709 14909 3743 14943
rect 4169 14909 4203 14943
rect 4353 14909 4387 14943
rect 6009 14909 6043 14943
rect 6653 14909 6687 14943
rect 7941 14909 7975 14943
rect 10150 14909 10184 14943
rect 16957 14909 16991 14943
rect 17233 14909 17267 14943
rect 22109 14909 22143 14943
rect 23765 14909 23799 14943
rect 24317 14841 24351 14875
rect 8125 14773 8159 14807
rect 9229 14773 9263 14807
rect 11805 14773 11839 14807
rect 18521 14773 18555 14807
rect 19165 14773 19199 14807
rect 21373 14773 21407 14807
rect 1869 14569 1903 14603
rect 3065 14569 3099 14603
rect 5365 14569 5399 14603
rect 6009 14569 6043 14603
rect 8217 14569 8251 14603
rect 11253 14569 11287 14603
rect 15117 14569 15151 14603
rect 24593 14569 24627 14603
rect 38117 14569 38151 14603
rect 20269 14501 20303 14535
rect 9321 14433 9355 14467
rect 18153 14433 18187 14467
rect 1777 14365 1811 14399
rect 2421 14365 2455 14399
rect 2605 14365 2639 14399
rect 3985 14365 4019 14399
rect 4629 14365 4663 14399
rect 5273 14365 5307 14399
rect 5917 14365 5951 14399
rect 8125 14365 8159 14399
rect 11161 14365 11195 14399
rect 11805 14365 11839 14399
rect 15025 14365 15059 14399
rect 22477 14365 22511 14399
rect 24777 14365 24811 14399
rect 38301 14365 38335 14399
rect 4077 14297 4111 14331
rect 6745 14297 6779 14331
rect 6837 14297 6871 14331
rect 7389 14297 7423 14331
rect 9413 14297 9447 14331
rect 10333 14297 10367 14331
rect 17877 14297 17911 14331
rect 17969 14297 18003 14331
rect 19717 14297 19751 14331
rect 19809 14297 19843 14331
rect 4721 14229 4755 14263
rect 11897 14229 11931 14263
rect 22569 14229 22603 14263
rect 27629 14229 27663 14263
rect 7297 14025 7331 14059
rect 8401 14025 8435 14059
rect 24409 14025 24443 14059
rect 2513 13957 2547 13991
rect 10425 13957 10459 13991
rect 11897 13957 11931 13991
rect 12817 13957 12851 13991
rect 15393 13957 15427 13991
rect 18429 13957 18463 13991
rect 19993 13957 20027 13991
rect 20177 13957 20211 13991
rect 27629 13957 27663 13991
rect 27721 13957 27755 13991
rect 1593 13889 1627 13923
rect 4445 13889 4479 13923
rect 5273 13889 5307 13923
rect 5733 13889 5767 13923
rect 6653 13889 6687 13923
rect 7757 13889 7791 13923
rect 8585 13889 8619 13923
rect 9229 13889 9263 13923
rect 9689 13889 9723 13923
rect 10333 13889 10367 13923
rect 10977 13889 11011 13923
rect 11069 13889 11103 13923
rect 13277 13889 13311 13923
rect 14565 13889 14599 13923
rect 18981 13889 19015 13923
rect 20637 13889 20671 13923
rect 24593 13889 24627 13923
rect 2421 13821 2455 13855
rect 3433 13821 3467 13855
rect 4537 13821 4571 13855
rect 6837 13821 6871 13855
rect 7849 13821 7883 13855
rect 11805 13821 11839 13855
rect 14657 13821 14691 13855
rect 15301 13821 15335 13855
rect 16313 13821 16347 13855
rect 18337 13821 18371 13855
rect 20729 13821 20763 13855
rect 27997 13821 28031 13855
rect 9045 13753 9079 13787
rect 1777 13685 1811 13719
rect 5089 13685 5123 13719
rect 5825 13685 5859 13719
rect 9781 13685 9815 13719
rect 13369 13685 13403 13719
rect 4077 13481 4111 13515
rect 5365 13481 5399 13515
rect 12081 13481 12115 13515
rect 12817 13481 12851 13515
rect 2053 13345 2087 13379
rect 2789 13345 2823 13379
rect 3433 13345 3467 13379
rect 6745 13345 6779 13379
rect 7021 13345 7055 13379
rect 9689 13345 9723 13379
rect 10241 13345 10275 13379
rect 14565 13345 14599 13379
rect 16405 13345 16439 13379
rect 16681 13345 16715 13379
rect 23305 13345 23339 13379
rect 30113 13345 30147 13379
rect 30573 13345 30607 13379
rect 3985 13277 4019 13311
rect 4813 13277 4847 13311
rect 5549 13277 5583 13311
rect 6009 13277 6043 13311
rect 8401 13277 8435 13311
rect 11437 13277 11471 13311
rect 11529 13277 11563 13311
rect 12265 13277 12299 13311
rect 12725 13277 12759 13311
rect 13553 13277 13587 13311
rect 14473 13277 14507 13311
rect 15669 13277 15703 13311
rect 17501 13279 17535 13313
rect 37289 13277 37323 13311
rect 38025 13277 38059 13311
rect 2881 13209 2915 13243
rect 6837 13209 6871 13243
rect 9781 13209 9815 13243
rect 13645 13209 13679 13243
rect 16497 13209 16531 13243
rect 23397 13209 23431 13243
rect 23949 13209 23983 13243
rect 30205 13209 30239 13243
rect 4629 13141 4663 13175
rect 6101 13141 6135 13175
rect 8493 13141 8527 13175
rect 15761 13141 15795 13175
rect 17601 13141 17635 13175
rect 37381 13141 37415 13175
rect 38209 13141 38243 13175
rect 2421 12937 2455 12971
rect 3157 12937 3191 12971
rect 3801 12937 3835 12971
rect 25881 12937 25915 12971
rect 4721 12869 4755 12903
rect 7573 12869 7607 12903
rect 10241 12869 10275 12903
rect 12357 12869 12391 12903
rect 17877 12869 17911 12903
rect 18797 12869 18831 12903
rect 23397 12869 23431 12903
rect 1593 12801 1627 12835
rect 2329 12801 2363 12835
rect 3065 12801 3099 12835
rect 3709 12801 3743 12835
rect 6745 12801 6779 12835
rect 13737 12801 13771 12835
rect 19901 12801 19935 12835
rect 22017 12801 22051 12835
rect 25789 12801 25823 12835
rect 38025 12801 38059 12835
rect 4629 12733 4663 12767
rect 5457 12733 5491 12767
rect 7389 12733 7423 12767
rect 8309 12733 8343 12767
rect 10149 12733 10183 12767
rect 10517 12733 10551 12767
rect 12265 12733 12299 12767
rect 12541 12733 12575 12767
rect 17785 12733 17819 12767
rect 23305 12733 23339 12767
rect 23581 12733 23615 12767
rect 1777 12597 1811 12631
rect 6837 12597 6871 12631
rect 13829 12597 13863 12631
rect 19993 12597 20027 12631
rect 22109 12597 22143 12631
rect 38209 12597 38243 12631
rect 2053 12393 2087 12427
rect 3985 12393 4019 12427
rect 7021 12393 7055 12427
rect 37841 12393 37875 12427
rect 8309 12325 8343 12359
rect 20729 12325 20763 12359
rect 3157 12257 3191 12291
rect 6837 12257 6871 12291
rect 7941 12257 7975 12291
rect 9229 12257 9263 12291
rect 9689 12257 9723 12291
rect 15945 12257 15979 12291
rect 16957 12257 16991 12291
rect 21925 12257 21959 12291
rect 23397 12257 23431 12291
rect 1961 12189 1995 12223
rect 4169 12189 4203 12223
rect 4721 12189 4755 12223
rect 5365 12189 5399 12223
rect 6009 12189 6043 12223
rect 6653 12189 6687 12223
rect 8125 12189 8159 12223
rect 10701 12189 10735 12223
rect 14289 12189 14323 12223
rect 15117 12189 15151 12223
rect 17785 12189 17819 12223
rect 19441 12189 19475 12223
rect 25053 12189 25087 12223
rect 25237 12189 25271 12223
rect 28457 12189 28491 12223
rect 38025 12189 38059 12223
rect 9321 12121 9355 12155
rect 10885 12121 10919 12155
rect 12541 12121 12575 12155
rect 13277 12121 13311 12155
rect 16037 12121 16071 12155
rect 20177 12121 20211 12155
rect 20269 12121 20303 12155
rect 22017 12121 22051 12155
rect 22937 12121 22971 12155
rect 28549 12121 28583 12155
rect 4813 12053 4847 12087
rect 5457 12053 5491 12087
rect 6101 12053 6135 12087
rect 13369 12053 13403 12087
rect 14381 12053 14415 12087
rect 15209 12053 15243 12087
rect 17877 12053 17911 12087
rect 19533 12053 19567 12087
rect 25697 12053 25731 12087
rect 3341 11849 3375 11883
rect 3985 11849 4019 11883
rect 9781 11849 9815 11883
rect 23765 11849 23799 11883
rect 25053 11849 25087 11883
rect 27813 11849 27847 11883
rect 5457 11781 5491 11815
rect 12265 11781 12299 11815
rect 13461 11781 13495 11815
rect 18429 11781 18463 11815
rect 19993 11781 20027 11815
rect 2053 11713 2087 11747
rect 2697 11713 2731 11747
rect 3525 11713 3559 11747
rect 4169 11713 4203 11747
rect 4629 11713 4663 11747
rect 6745 11713 6779 11747
rect 7205 11713 7239 11747
rect 8217 11713 8251 11747
rect 9689 11713 9723 11747
rect 10333 11713 10367 11747
rect 10977 11713 11011 11747
rect 14473 11713 14507 11747
rect 14657 11713 14691 11747
rect 15761 11713 15795 11747
rect 22477 11713 22511 11747
rect 22569 11713 22603 11747
rect 23305 11713 23339 11747
rect 24961 11713 24995 11747
rect 25789 11713 25823 11747
rect 28273 11713 28307 11747
rect 5365 11645 5399 11679
rect 5641 11645 5675 11679
rect 7757 11645 7791 11679
rect 8033 11645 8067 11679
rect 12173 11645 12207 11679
rect 13369 11645 13403 11679
rect 15117 11645 15151 11679
rect 18337 11645 18371 11679
rect 18981 11645 19015 11679
rect 19901 11645 19935 11679
rect 20545 11645 20579 11679
rect 23121 11645 23155 11679
rect 24317 11645 24351 11679
rect 27169 11645 27203 11679
rect 27353 11645 27387 11679
rect 7297 11577 7331 11611
rect 10425 11577 10459 11611
rect 12725 11577 12759 11611
rect 13921 11577 13955 11611
rect 2145 11509 2179 11543
rect 2789 11509 2823 11543
rect 4721 11509 4755 11543
rect 6837 11509 6871 11543
rect 8401 11509 8435 11543
rect 11069 11509 11103 11543
rect 15577 11509 15611 11543
rect 25605 11509 25639 11543
rect 28365 11509 28399 11543
rect 1777 11305 1811 11339
rect 3985 11305 4019 11339
rect 9689 11305 9723 11339
rect 26341 11305 26375 11339
rect 3341 11237 3375 11271
rect 6837 11237 6871 11271
rect 28089 11237 28123 11271
rect 5641 11169 5675 11203
rect 8585 11169 8619 11203
rect 11345 11169 11379 11203
rect 13645 11169 13679 11203
rect 19533 11169 19567 11203
rect 20361 11169 20395 11203
rect 22661 11169 22695 11203
rect 23397 11169 23431 11203
rect 24685 11169 24719 11203
rect 26985 11169 27019 11203
rect 37749 11169 37783 11203
rect 1961 11101 1995 11135
rect 2421 11101 2455 11135
rect 3249 11101 3283 11135
rect 4169 11101 4203 11135
rect 4629 11101 4663 11135
rect 7021 11101 7055 11135
rect 9137 11101 9171 11135
rect 9321 11101 9355 11135
rect 10333 11101 10367 11135
rect 15025 11101 15059 11135
rect 21097 11101 21131 11135
rect 22569 11101 22603 11135
rect 23213 11101 23247 11135
rect 26525 11101 26559 11135
rect 27997 11101 28031 11135
rect 31861 11101 31895 11135
rect 37473 11101 37507 11135
rect 5365 11033 5399 11067
rect 5457 11033 5491 11067
rect 7573 11033 7607 11067
rect 7665 11033 7699 11067
rect 10425 11033 10459 11067
rect 11069 11033 11103 11067
rect 11161 11033 11195 11067
rect 12633 11033 12667 11067
rect 12725 11033 12759 11067
rect 15577 11033 15611 11067
rect 15669 11033 15703 11067
rect 16221 11033 16255 11067
rect 19625 11033 19659 11067
rect 23857 11033 23891 11067
rect 24777 11033 24811 11067
rect 25329 11033 25363 11067
rect 31953 11033 31987 11067
rect 2513 10965 2547 10999
rect 4721 10965 4755 10999
rect 14841 10965 14875 10999
rect 21189 10965 21223 10999
rect 5365 10761 5399 10795
rect 7665 10761 7699 10795
rect 10977 10761 11011 10795
rect 13553 10761 13587 10795
rect 14197 10761 14231 10795
rect 19073 10761 19107 10795
rect 19901 10761 19935 10795
rect 23857 10761 23891 10795
rect 2605 10693 2639 10727
rect 3525 10693 3559 10727
rect 8493 10693 8527 10727
rect 9045 10693 9079 10727
rect 9689 10693 9723 10727
rect 10241 10693 10275 10727
rect 11897 10693 11931 10727
rect 17969 10693 18003 10727
rect 1777 10625 1811 10659
rect 4261 10625 4295 10659
rect 6745 10625 6779 10659
rect 7849 10625 7883 10659
rect 10885 10625 10919 10659
rect 12909 10625 12943 10659
rect 13737 10625 13771 10659
rect 14381 10625 14415 10659
rect 15117 10625 15151 10659
rect 17141 10625 17175 10659
rect 18981 10625 19015 10659
rect 19809 10625 19843 10659
rect 21005 10625 21039 10659
rect 23305 10625 23339 10659
rect 23765 10625 23799 10659
rect 25053 10625 25087 10659
rect 2513 10557 2547 10591
rect 4077 10557 4111 10591
rect 6561 10557 6595 10591
rect 8401 10557 8435 10591
rect 9597 10557 9631 10591
rect 11805 10557 11839 10591
rect 12081 10557 12115 10591
rect 14933 10557 14967 10591
rect 17877 10557 17911 10591
rect 18153 10557 18187 10591
rect 20821 10557 20855 10591
rect 22017 10557 22051 10591
rect 22201 10557 22235 10591
rect 22661 10557 22695 10591
rect 1869 10421 1903 10455
rect 4445 10421 4479 10455
rect 6929 10421 6963 10455
rect 13001 10421 13035 10455
rect 15301 10421 15335 10455
rect 17233 10421 17267 10455
rect 21189 10421 21223 10455
rect 23121 10421 23155 10455
rect 24869 10421 24903 10455
rect 9597 10217 9631 10251
rect 13369 10217 13403 10251
rect 19901 10217 19935 10251
rect 22293 10217 22327 10251
rect 25237 10217 25271 10251
rect 2881 10149 2915 10183
rect 12449 10149 12483 10183
rect 2329 10081 2363 10115
rect 7665 10081 7699 10115
rect 18337 10081 18371 10115
rect 1777 10013 1811 10047
rect 5181 10013 5215 10047
rect 6837 10013 6871 10047
rect 8401 10013 8435 10047
rect 9781 10013 9815 10047
rect 11069 10013 11103 10047
rect 12357 10013 12391 10047
rect 13277 10013 13311 10047
rect 19809 10013 19843 10047
rect 22477 10013 22511 10047
rect 24777 10013 24811 10047
rect 25421 10013 25455 10047
rect 38025 10013 38059 10047
rect 2421 9945 2455 9979
rect 6929 9945 6963 9979
rect 17325 9945 17359 9979
rect 17417 9945 17451 9979
rect 1593 9877 1627 9911
rect 4997 9877 5031 9911
rect 8493 9877 8527 9911
rect 11161 9877 11195 9911
rect 24593 9877 24627 9911
rect 38209 9877 38243 9911
rect 2053 9673 2087 9707
rect 21005 9673 21039 9707
rect 8217 9605 8251 9639
rect 9229 9605 9263 9639
rect 11897 9605 11931 9639
rect 32413 9605 32447 9639
rect 1961 9537 1995 9571
rect 2789 9537 2823 9571
rect 3985 9537 4019 9571
rect 4629 9537 4663 9571
rect 5825 9537 5859 9571
rect 5917 9537 5951 9571
rect 6561 9537 6595 9571
rect 7205 9537 7239 9571
rect 8125 9537 8159 9571
rect 10241 9537 10275 9571
rect 19717 9537 19751 9571
rect 32321 9537 32355 9571
rect 34897 9537 34931 9571
rect 9137 9469 9171 9503
rect 10517 9469 10551 9503
rect 11805 9469 11839 9503
rect 20361 9469 20395 9503
rect 20545 9469 20579 9503
rect 34345 9469 34379 9503
rect 2605 9401 2639 9435
rect 4445 9401 4479 9435
rect 9689 9401 9723 9435
rect 12357 9401 12391 9435
rect 34713 9401 34747 9435
rect 3801 9333 3835 9367
rect 6653 9333 6687 9367
rect 7297 9333 7331 9367
rect 19809 9333 19843 9367
rect 1593 9129 1627 9163
rect 9229 9129 9263 9163
rect 11437 9129 11471 9163
rect 12081 9129 12115 9163
rect 26341 9129 26375 9163
rect 2329 9061 2363 9095
rect 5457 9061 5491 9095
rect 20453 8993 20487 9027
rect 1777 8925 1811 8959
rect 2237 8925 2271 8959
rect 4169 8925 4203 8959
rect 5641 8925 5675 8959
rect 9137 8925 9171 8959
rect 11345 8925 11379 8959
rect 11989 8925 12023 8959
rect 24593 8925 24627 8959
rect 26341 8925 26375 8959
rect 32597 8925 32631 8959
rect 2881 8789 2915 8823
rect 3985 8789 4019 8823
rect 4629 8789 4663 8823
rect 24685 8789 24719 8823
rect 32413 8789 32447 8823
rect 2237 8585 2271 8619
rect 3525 8585 3559 8619
rect 4629 8585 4663 8619
rect 2145 8449 2179 8483
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 3985 8449 4019 8483
rect 14565 8449 14599 8483
rect 21005 8449 21039 8483
rect 27169 8449 27203 8483
rect 38117 8449 38151 8483
rect 4169 8381 4203 8415
rect 38301 8381 38335 8415
rect 14657 8313 14691 8347
rect 27261 8313 27295 8347
rect 20821 8245 20855 8279
rect 4077 8041 4111 8075
rect 14841 8041 14875 8075
rect 20821 8041 20855 8075
rect 1869 7905 1903 7939
rect 1593 7837 1627 7871
rect 3157 7837 3191 7871
rect 3985 7837 4019 7871
rect 11069 7837 11103 7871
rect 14749 7837 14783 7871
rect 18889 7837 18923 7871
rect 21005 7837 21039 7871
rect 24777 7837 24811 7871
rect 29193 7837 29227 7871
rect 33793 7837 33827 7871
rect 38025 7837 38059 7871
rect 3249 7701 3283 7735
rect 10885 7701 10919 7735
rect 18705 7701 18739 7735
rect 24593 7701 24627 7735
rect 29009 7701 29043 7735
rect 33885 7701 33919 7735
rect 38209 7701 38243 7735
rect 2421 7429 2455 7463
rect 2513 7429 2547 7463
rect 1685 7361 1719 7395
rect 4629 7361 4663 7395
rect 14197 7361 14231 7395
rect 16865 7361 16899 7395
rect 35081 7361 35115 7395
rect 2973 7225 3007 7259
rect 14013 7225 14047 7259
rect 1777 7157 1811 7191
rect 4445 7157 4479 7191
rect 16957 7157 16991 7191
rect 34897 7157 34931 7191
rect 2329 6817 2363 6851
rect 1777 6749 1811 6783
rect 2237 6749 2271 6783
rect 35081 6749 35115 6783
rect 1593 6613 1627 6647
rect 34897 6613 34931 6647
rect 37749 6273 37783 6307
rect 15209 6205 15243 6239
rect 37473 6205 37507 6239
rect 2881 5865 2915 5899
rect 15209 5729 15243 5763
rect 15485 5729 15519 5763
rect 1593 5661 1627 5695
rect 2789 5661 2823 5695
rect 4445 5661 4479 5695
rect 23857 5661 23891 5695
rect 15301 5593 15335 5627
rect 1777 5525 1811 5559
rect 4537 5525 4571 5559
rect 23949 5525 23983 5559
rect 4721 5185 4755 5219
rect 9505 5185 9539 5219
rect 24777 5185 24811 5219
rect 38025 5185 38059 5219
rect 4537 4981 4571 5015
rect 9321 4981 9355 5015
rect 24593 4981 24627 5015
rect 38209 4981 38243 5015
rect 33149 4573 33183 4607
rect 33241 4573 33275 4607
rect 35541 4573 35575 4607
rect 38025 4573 38059 4607
rect 1685 4505 1719 4539
rect 1777 4437 1811 4471
rect 35357 4437 35391 4471
rect 38209 4437 38243 4471
rect 38025 4097 38059 4131
rect 38209 3893 38243 3927
rect 1593 3689 1627 3723
rect 1777 3485 1811 3519
rect 37565 3485 37599 3519
rect 38025 3485 38059 3519
rect 37381 3349 37415 3383
rect 38209 3349 38243 3383
rect 2329 3145 2363 3179
rect 36737 3145 36771 3179
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 3525 3009 3559 3043
rect 11989 3009 12023 3043
rect 17049 3009 17083 3043
rect 18889 3009 18923 3043
rect 25789 3009 25823 3043
rect 36921 3009 36955 3043
rect 37749 3009 37783 3043
rect 11713 2941 11747 2975
rect 37473 2941 37507 2975
rect 3341 2873 3375 2907
rect 1777 2805 1811 2839
rect 16865 2805 16899 2839
rect 18705 2805 18739 2839
rect 25605 2805 25639 2839
rect 7205 2601 7239 2635
rect 9781 2601 9815 2635
rect 14289 2601 14323 2635
rect 18245 2601 18279 2635
rect 22017 2601 22051 2635
rect 24593 2601 24627 2635
rect 27169 2601 27203 2635
rect 28641 2601 28675 2635
rect 3249 2533 3283 2567
rect 13185 2465 13219 2499
rect 19717 2465 19751 2499
rect 37749 2465 37783 2499
rect 2329 2397 2363 2431
rect 3065 2397 3099 2431
rect 3985 2397 4019 2431
rect 4997 2397 5031 2431
rect 5273 2397 5307 2431
rect 6745 2397 6779 2431
rect 7389 2397 7423 2431
rect 9321 2397 9355 2431
rect 9965 2397 9999 2431
rect 11713 2397 11747 2431
rect 12909 2397 12943 2431
rect 14473 2397 14507 2431
rect 14933 2397 14967 2431
rect 16037 2397 16071 2431
rect 17509 2397 17543 2431
rect 18429 2397 18463 2431
rect 19441 2397 19475 2431
rect 20729 2397 20763 2431
rect 22201 2397 22235 2431
rect 22661 2397 22695 2431
rect 24777 2397 24811 2431
rect 25237 2397 25271 2431
rect 25973 2397 26007 2431
rect 27353 2397 27387 2431
rect 29745 2397 29779 2431
rect 30481 2397 30515 2431
rect 32321 2397 32355 2431
rect 33057 2397 33091 2431
rect 33793 2397 33827 2431
rect 34897 2397 34931 2431
rect 36185 2397 36219 2431
rect 37473 2397 37507 2431
rect 1685 2329 1719 2363
rect 28549 2329 28583 2363
rect 1777 2261 1811 2295
rect 2513 2261 2547 2295
rect 4169 2261 4203 2295
rect 5457 2261 5491 2295
rect 6561 2261 6595 2295
rect 9137 2261 9171 2295
rect 11897 2261 11931 2295
rect 15117 2261 15151 2295
rect 16221 2261 16255 2295
rect 17693 2261 17727 2295
rect 20913 2261 20947 2295
rect 22845 2261 22879 2295
rect 25421 2261 25455 2295
rect 26157 2261 26191 2295
rect 29929 2261 29963 2295
rect 30665 2261 30699 2295
rect 32505 2261 32539 2295
rect 33241 2261 33275 2295
rect 33977 2261 34011 2295
rect 35081 2261 35115 2295
rect 36369 2261 36403 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1762 37448 1768 37460
rect 1723 37420 1768 37448
rect 1762 37408 1768 37420
rect 1820 37408 1826 37460
rect 25038 37408 25044 37460
rect 25096 37448 25102 37460
rect 26329 37451 26387 37457
rect 26329 37448 26341 37451
rect 25096 37420 26341 37448
rect 25096 37408 25102 37420
rect 26329 37417 26341 37420
rect 26375 37417 26387 37451
rect 26329 37411 26387 37417
rect 5813 37383 5871 37389
rect 5813 37349 5825 37383
rect 5859 37380 5871 37383
rect 6086 37380 6092 37392
rect 5859 37352 6092 37380
rect 5859 37349 5871 37352
rect 5813 37343 5871 37349
rect 6086 37340 6092 37352
rect 6144 37340 6150 37392
rect 19429 37383 19487 37389
rect 19429 37349 19441 37383
rect 19475 37380 19487 37383
rect 25406 37380 25412 37392
rect 19475 37352 25412 37380
rect 19475 37349 19487 37352
rect 19429 37343 19487 37349
rect 25406 37340 25412 37352
rect 25464 37340 25470 37392
rect 25777 37383 25835 37389
rect 25777 37349 25789 37383
rect 25823 37380 25835 37383
rect 26234 37380 26240 37392
rect 25823 37352 26240 37380
rect 25823 37349 25835 37352
rect 25777 37343 25835 37349
rect 26234 37340 26240 37352
rect 26292 37340 26298 37392
rect 12250 37272 12256 37324
rect 12308 37312 12314 37324
rect 12345 37315 12403 37321
rect 12345 37312 12357 37315
rect 12308 37284 12357 37312
rect 12308 37272 12314 37284
rect 12345 37281 12357 37284
rect 12391 37281 12403 37315
rect 12345 37275 12403 37281
rect 16960 37284 18828 37312
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37244 1639 37247
rect 2314 37244 2320 37256
rect 1627 37216 2320 37244
rect 1627 37213 1639 37216
rect 1581 37207 1639 37213
rect 2314 37204 2320 37216
rect 2372 37204 2378 37256
rect 2774 37204 2780 37256
rect 2832 37244 2838 37256
rect 2869 37247 2927 37253
rect 2869 37244 2881 37247
rect 2832 37216 2881 37244
rect 2832 37204 2838 37216
rect 2869 37213 2881 37216
rect 2915 37213 2927 37247
rect 2869 37207 2927 37213
rect 2958 37204 2964 37256
rect 3016 37244 3022 37256
rect 3973 37247 4031 37253
rect 3973 37244 3985 37247
rect 3016 37216 3985 37244
rect 3016 37204 3022 37216
rect 3973 37213 3985 37216
rect 4019 37213 4031 37247
rect 3973 37207 4031 37213
rect 4614 37204 4620 37256
rect 4672 37244 4678 37256
rect 4893 37247 4951 37253
rect 4893 37244 4905 37247
rect 4672 37216 4905 37244
rect 4672 37204 4678 37216
rect 4893 37213 4905 37216
rect 4939 37213 4951 37247
rect 4893 37207 4951 37213
rect 5997 37247 6055 37253
rect 5997 37213 6009 37247
rect 6043 37244 6055 37247
rect 6454 37244 6460 37256
rect 6043 37216 6460 37244
rect 6043 37213 6055 37216
rect 5997 37207 6055 37213
rect 6454 37204 6460 37216
rect 6512 37204 6518 37256
rect 6546 37204 6552 37256
rect 6604 37244 6610 37256
rect 6604 37216 6649 37244
rect 6604 37204 6610 37216
rect 7742 37204 7748 37256
rect 7800 37244 7806 37256
rect 7929 37247 7987 37253
rect 7929 37244 7941 37247
rect 7800 37216 7941 37244
rect 7800 37204 7806 37216
rect 7929 37213 7941 37216
rect 7975 37213 7987 37247
rect 7929 37207 7987 37213
rect 9401 37247 9459 37253
rect 9401 37213 9413 37247
rect 9447 37213 9459 37247
rect 9401 37207 9459 37213
rect 9416 37176 9444 37207
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 10229 37247 10287 37253
rect 10229 37244 10241 37247
rect 9732 37216 10241 37244
rect 9732 37204 9738 37216
rect 10229 37213 10241 37216
rect 10275 37213 10287 37247
rect 10229 37207 10287 37213
rect 10873 37247 10931 37253
rect 10873 37213 10885 37247
rect 10919 37244 10931 37247
rect 12621 37247 12679 37253
rect 10919 37216 12434 37244
rect 10919 37213 10931 37216
rect 10873 37207 10931 37213
rect 2700 37148 9444 37176
rect 2700 37117 2728 37148
rect 2685 37111 2743 37117
rect 2685 37077 2697 37111
rect 2731 37077 2743 37111
rect 2685 37071 2743 37077
rect 3234 37068 3240 37120
rect 3292 37108 3298 37120
rect 4157 37111 4215 37117
rect 4157 37108 4169 37111
rect 3292 37080 4169 37108
rect 3292 37068 3298 37080
rect 4157 37077 4169 37080
rect 4203 37077 4215 37111
rect 4157 37071 4215 37077
rect 4709 37111 4767 37117
rect 4709 37077 4721 37111
rect 4755 37108 4767 37111
rect 5718 37108 5724 37120
rect 4755 37080 5724 37108
rect 4755 37077 4767 37080
rect 4709 37071 4767 37077
rect 5718 37068 5724 37080
rect 5776 37068 5782 37120
rect 5994 37068 6000 37120
rect 6052 37108 6058 37120
rect 6733 37111 6791 37117
rect 6733 37108 6745 37111
rect 6052 37080 6745 37108
rect 6052 37068 6058 37080
rect 6733 37077 6745 37080
rect 6779 37077 6791 37111
rect 8018 37108 8024 37120
rect 7979 37080 8024 37108
rect 6733 37071 6791 37077
rect 8018 37068 8024 37080
rect 8076 37068 8082 37120
rect 9490 37108 9496 37120
rect 9451 37080 9496 37108
rect 9490 37068 9496 37080
rect 9548 37068 9554 37120
rect 10045 37111 10103 37117
rect 10045 37077 10057 37111
rect 10091 37108 10103 37111
rect 10870 37108 10876 37120
rect 10091 37080 10876 37108
rect 10091 37077 10103 37080
rect 10045 37071 10103 37077
rect 10870 37068 10876 37080
rect 10928 37068 10934 37120
rect 11054 37108 11060 37120
rect 11015 37080 11060 37108
rect 11054 37068 11060 37080
rect 11112 37068 11118 37120
rect 12406 37108 12434 37216
rect 12621 37213 12633 37247
rect 12667 37244 12679 37247
rect 13998 37244 14004 37256
rect 12667 37216 14004 37244
rect 12667 37213 12679 37216
rect 12621 37207 12679 37213
rect 13998 37204 14004 37216
rect 14056 37204 14062 37256
rect 14182 37204 14188 37256
rect 14240 37244 14246 37256
rect 14461 37247 14519 37253
rect 14461 37244 14473 37247
rect 14240 37216 14473 37244
rect 14240 37204 14246 37216
rect 14461 37213 14473 37216
rect 14507 37213 14519 37247
rect 14461 37207 14519 37213
rect 15105 37247 15163 37253
rect 15105 37213 15117 37247
rect 15151 37213 15163 37247
rect 15562 37244 15568 37256
rect 15523 37216 15568 37244
rect 15105 37207 15163 37213
rect 13538 37136 13544 37188
rect 13596 37176 13602 37188
rect 15120 37176 15148 37207
rect 15562 37204 15568 37216
rect 15620 37204 15626 37256
rect 16960 37176 16988 37284
rect 17037 37247 17095 37253
rect 17037 37213 17049 37247
rect 17083 37213 17095 37247
rect 17037 37207 17095 37213
rect 17497 37247 17555 37253
rect 17497 37213 17509 37247
rect 17543 37244 17555 37247
rect 17770 37244 17776 37256
rect 17543 37216 17776 37244
rect 17543 37213 17555 37216
rect 17497 37207 17555 37213
rect 13596 37148 15148 37176
rect 15212 37148 16988 37176
rect 17052 37176 17080 37207
rect 17770 37204 17776 37216
rect 17828 37204 17834 37256
rect 17862 37204 17868 37256
rect 17920 37244 17926 37256
rect 18693 37247 18751 37253
rect 18693 37244 18705 37247
rect 17920 37216 18705 37244
rect 17920 37204 17926 37216
rect 18693 37213 18705 37216
rect 18739 37213 18751 37247
rect 18800 37244 18828 37284
rect 21266 37272 21272 37324
rect 21324 37312 21330 37324
rect 22005 37315 22063 37321
rect 22005 37312 22017 37315
rect 21324 37284 22017 37312
rect 21324 37272 21330 37284
rect 22005 37281 22017 37284
rect 22051 37281 22063 37315
rect 22005 37275 22063 37281
rect 23198 37272 23204 37324
rect 23256 37312 23262 37324
rect 23256 37284 26096 37312
rect 23256 37272 23262 37284
rect 19426 37244 19432 37256
rect 18800 37216 19432 37244
rect 18693 37207 18751 37213
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 19613 37247 19671 37253
rect 19613 37213 19625 37247
rect 19659 37213 19671 37247
rect 19613 37207 19671 37213
rect 20073 37247 20131 37253
rect 20073 37213 20085 37247
rect 20119 37244 20131 37247
rect 20990 37244 20996 37256
rect 20119 37216 20852 37244
rect 20951 37216 20996 37244
rect 20119 37213 20131 37216
rect 20073 37207 20131 37213
rect 18598 37176 18604 37188
rect 17052 37148 18604 37176
rect 13596 37136 13602 37148
rect 14090 37108 14096 37120
rect 12406 37080 14096 37108
rect 14090 37068 14096 37080
rect 14148 37068 14154 37120
rect 14274 37108 14280 37120
rect 14235 37080 14280 37108
rect 14274 37068 14280 37080
rect 14332 37068 14338 37120
rect 14918 37108 14924 37120
rect 14879 37080 14924 37108
rect 14918 37068 14924 37080
rect 14976 37068 14982 37120
rect 15010 37068 15016 37120
rect 15068 37108 15074 37120
rect 15212 37108 15240 37148
rect 18598 37136 18604 37148
rect 18656 37136 18662 37188
rect 19628 37176 19656 37207
rect 20714 37176 20720 37188
rect 19628 37148 20720 37176
rect 20714 37136 20720 37148
rect 20772 37136 20778 37188
rect 15068 37080 15240 37108
rect 15068 37068 15074 37080
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 15749 37111 15807 37117
rect 15749 37108 15761 37111
rect 15528 37080 15761 37108
rect 15528 37068 15534 37080
rect 15749 37077 15761 37080
rect 15795 37077 15807 37111
rect 15749 37071 15807 37077
rect 16853 37111 16911 37117
rect 16853 37077 16865 37111
rect 16899 37108 16911 37111
rect 17218 37108 17224 37120
rect 16899 37080 17224 37108
rect 16899 37077 16911 37080
rect 16853 37071 16911 37077
rect 17218 37068 17224 37080
rect 17276 37068 17282 37120
rect 17402 37068 17408 37120
rect 17460 37108 17466 37120
rect 17681 37111 17739 37117
rect 17681 37108 17693 37111
rect 17460 37080 17693 37108
rect 17460 37068 17466 37080
rect 17681 37077 17693 37080
rect 17727 37077 17739 37111
rect 18782 37108 18788 37120
rect 18743 37080 18788 37108
rect 17681 37071 17739 37077
rect 18782 37068 18788 37080
rect 18840 37068 18846 37120
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20824 37117 20852 37216
rect 20990 37204 20996 37216
rect 21048 37204 21054 37256
rect 22281 37247 22339 37253
rect 22281 37213 22293 37247
rect 22327 37244 22339 37247
rect 22554 37244 22560 37256
rect 22327 37216 22560 37244
rect 22327 37213 22339 37216
rect 22281 37207 22339 37213
rect 22554 37204 22560 37216
rect 22612 37204 22618 37256
rect 23106 37204 23112 37256
rect 23164 37244 23170 37256
rect 23293 37247 23351 37253
rect 23293 37244 23305 37247
rect 23164 37216 23305 37244
rect 23164 37204 23170 37216
rect 23293 37213 23305 37216
rect 23339 37213 23351 37247
rect 23293 37207 23351 37213
rect 23382 37204 23388 37256
rect 23440 37244 23446 37256
rect 25038 37244 25044 37256
rect 23440 37216 25044 37244
rect 23440 37204 23446 37216
rect 25038 37204 25044 37216
rect 25096 37204 25102 37256
rect 26068 37244 26096 37284
rect 27264 37284 27936 37312
rect 26513 37247 26571 37253
rect 26513 37244 26525 37247
rect 26068 37216 26525 37244
rect 26513 37213 26525 37216
rect 26559 37213 26571 37247
rect 26513 37207 26571 37213
rect 26602 37204 26608 37256
rect 26660 37244 26666 37256
rect 27264 37244 27292 37284
rect 26660 37216 27292 37244
rect 27341 37247 27399 37253
rect 26660 37204 26666 37216
rect 27341 37213 27353 37247
rect 27387 37213 27399 37247
rect 27798 37244 27804 37256
rect 27759 37216 27804 37244
rect 27341 37207 27399 37213
rect 20898 37136 20904 37188
rect 20956 37176 20962 37188
rect 21910 37176 21916 37188
rect 20956 37148 21916 37176
rect 20956 37136 20962 37148
rect 21910 37136 21916 37148
rect 21968 37136 21974 37188
rect 25222 37176 25228 37188
rect 25183 37148 25228 37176
rect 25222 37136 25228 37148
rect 25280 37136 25286 37188
rect 25314 37136 25320 37188
rect 25372 37176 25378 37188
rect 27356 37176 27384 37207
rect 27798 37204 27804 37216
rect 27856 37204 27862 37256
rect 27908 37244 27936 37284
rect 28460 37284 28764 37312
rect 28460 37244 28488 37284
rect 27908 37216 28488 37244
rect 28534 37204 28540 37256
rect 28592 37244 28598 37256
rect 28736 37244 28764 37284
rect 30374 37272 30380 37324
rect 30432 37312 30438 37324
rect 30653 37315 30711 37321
rect 30653 37312 30665 37315
rect 30432 37284 30665 37312
rect 30432 37272 30438 37284
rect 30653 37281 30665 37284
rect 30699 37281 30711 37315
rect 30653 37275 30711 37281
rect 30926 37272 30932 37324
rect 30984 37312 30990 37324
rect 32309 37315 32367 37321
rect 32309 37312 32321 37315
rect 30984 37284 32321 37312
rect 30984 37272 30990 37284
rect 32309 37281 32321 37284
rect 32355 37281 32367 37315
rect 32309 37275 32367 37281
rect 32582 37244 32588 37256
rect 28592 37216 28637 37244
rect 28736 37216 29040 37244
rect 32543 37216 32588 37244
rect 28592 37204 28598 37216
rect 28902 37176 28908 37188
rect 25372 37148 25417 37176
rect 26252 37148 27384 37176
rect 27632 37148 28908 37176
rect 25372 37136 25378 37148
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 20809 37111 20867 37117
rect 20809 37077 20821 37111
rect 20855 37077 20867 37111
rect 20809 37071 20867 37077
rect 23382 37068 23388 37120
rect 23440 37108 23446 37120
rect 23440 37080 23485 37108
rect 23440 37068 23446 37080
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 26252 37108 26280 37148
rect 24544 37080 26280 37108
rect 27157 37111 27215 37117
rect 24544 37068 24550 37080
rect 27157 37077 27169 37111
rect 27203 37108 27215 37111
rect 27632 37108 27660 37148
rect 28902 37136 28908 37148
rect 28960 37136 28966 37188
rect 29012 37176 29040 37216
rect 32582 37204 32588 37216
rect 32640 37204 32646 37256
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 34848 37216 34897 37244
rect 34848 37204 34854 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 36078 37204 36084 37256
rect 36136 37244 36142 37256
rect 36265 37247 36323 37253
rect 36265 37244 36277 37247
rect 36136 37216 36277 37244
rect 36136 37204 36142 37216
rect 36265 37213 36277 37216
rect 36311 37213 36323 37247
rect 36265 37207 36323 37213
rect 37366 37204 37372 37256
rect 37424 37244 37430 37256
rect 37553 37247 37611 37253
rect 37553 37244 37565 37247
rect 37424 37216 37565 37244
rect 37424 37204 37430 37216
rect 37553 37213 37565 37216
rect 37599 37213 37611 37247
rect 37553 37207 37611 37213
rect 30377 37179 30435 37185
rect 30377 37176 30389 37179
rect 29012 37148 30389 37176
rect 30377 37145 30389 37148
rect 30423 37145 30435 37179
rect 30377 37139 30435 37145
rect 30466 37136 30472 37188
rect 30524 37176 30530 37188
rect 30524 37148 30569 37176
rect 30524 37136 30530 37148
rect 27203 37080 27660 37108
rect 27203 37077 27215 37080
rect 27157 37071 27215 37077
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 27985 37111 28043 37117
rect 27985 37108 27997 37111
rect 27764 37080 27997 37108
rect 27764 37068 27770 37080
rect 27985 37077 27997 37080
rect 28031 37077 28043 37111
rect 28626 37108 28632 37120
rect 28587 37080 28632 37108
rect 27985 37071 28043 37077
rect 28626 37068 28632 37080
rect 28684 37068 28690 37120
rect 33134 37068 33140 37120
rect 33192 37108 33198 37120
rect 33781 37111 33839 37117
rect 33781 37108 33793 37111
rect 33192 37080 33793 37108
rect 33192 37068 33198 37080
rect 33781 37077 33793 37080
rect 33827 37077 33839 37111
rect 33781 37071 33839 37077
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 35069 37111 35127 37117
rect 35069 37108 35081 37111
rect 34572 37080 35081 37108
rect 34572 37068 34578 37080
rect 35069 37077 35081 37080
rect 35115 37077 35127 37111
rect 36354 37108 36360 37120
rect 36315 37080 36360 37108
rect 35069 37071 35127 37077
rect 36354 37068 36360 37080
rect 36412 37068 36418 37120
rect 37642 37108 37648 37120
rect 37603 37080 37648 37108
rect 37642 37068 37648 37080
rect 37700 37068 37706 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 6546 36864 6552 36916
rect 6604 36904 6610 36916
rect 10134 36904 10140 36916
rect 6604 36876 10140 36904
rect 6604 36864 6610 36876
rect 10134 36864 10140 36876
rect 10192 36864 10198 36916
rect 10870 36864 10876 36916
rect 10928 36904 10934 36916
rect 10928 36876 12112 36904
rect 10928 36864 10934 36876
rect 6086 36796 6092 36848
rect 6144 36836 6150 36848
rect 11974 36836 11980 36848
rect 6144 36808 11980 36836
rect 6144 36796 6150 36808
rect 11974 36796 11980 36808
rect 12032 36796 12038 36848
rect 1302 36728 1308 36780
rect 1360 36768 1366 36780
rect 1765 36771 1823 36777
rect 1765 36768 1777 36771
rect 1360 36740 1777 36768
rect 1360 36728 1366 36740
rect 1765 36737 1777 36740
rect 1811 36737 1823 36771
rect 1765 36731 1823 36737
rect 2593 36771 2651 36777
rect 2593 36737 2605 36771
rect 2639 36768 2651 36771
rect 4706 36768 4712 36780
rect 2639 36740 2774 36768
rect 4667 36740 4712 36768
rect 2639 36737 2651 36740
rect 2593 36731 2651 36737
rect 2746 36632 2774 36740
rect 4706 36728 4712 36740
rect 4764 36728 4770 36780
rect 5718 36728 5724 36780
rect 5776 36768 5782 36780
rect 7009 36771 7067 36777
rect 7009 36768 7021 36771
rect 5776 36740 7021 36768
rect 5776 36728 5782 36740
rect 7009 36737 7021 36740
rect 7055 36737 7067 36771
rect 7650 36768 7656 36780
rect 7611 36740 7656 36768
rect 7009 36731 7067 36737
rect 7650 36728 7656 36740
rect 7708 36728 7714 36780
rect 9030 36728 9036 36780
rect 9088 36768 9094 36780
rect 10505 36771 10563 36777
rect 10505 36768 10517 36771
rect 9088 36740 10517 36768
rect 9088 36728 9094 36740
rect 10505 36737 10517 36740
rect 10551 36737 10563 36771
rect 10505 36731 10563 36737
rect 7101 36703 7159 36709
rect 7101 36669 7113 36703
rect 7147 36700 7159 36703
rect 8481 36703 8539 36709
rect 8481 36700 8493 36703
rect 7147 36672 8493 36700
rect 7147 36669 7159 36672
rect 7101 36663 7159 36669
rect 8481 36669 8493 36672
rect 8527 36669 8539 36703
rect 8662 36700 8668 36712
rect 8623 36672 8668 36700
rect 8481 36663 8539 36669
rect 8662 36660 8668 36672
rect 8720 36660 8726 36712
rect 9677 36703 9735 36709
rect 9677 36669 9689 36703
rect 9723 36700 9735 36703
rect 10410 36700 10416 36712
rect 9723 36672 10416 36700
rect 9723 36669 9735 36672
rect 9677 36663 9735 36669
rect 10410 36660 10416 36672
rect 10468 36660 10474 36712
rect 3418 36632 3424 36644
rect 2746 36604 3424 36632
rect 3418 36592 3424 36604
rect 3476 36632 3482 36644
rect 11882 36632 11888 36644
rect 3476 36604 11888 36632
rect 3476 36592 3482 36604
rect 11882 36592 11888 36604
rect 11940 36592 11946 36644
rect 12084 36632 12112 36876
rect 12894 36864 12900 36916
rect 12952 36904 12958 36916
rect 13906 36904 13912 36916
rect 12952 36876 13912 36904
rect 12952 36864 12958 36876
rect 13906 36864 13912 36876
rect 13964 36904 13970 36916
rect 14826 36904 14832 36916
rect 13964 36876 14832 36904
rect 13964 36864 13970 36876
rect 14826 36864 14832 36876
rect 14884 36864 14890 36916
rect 14918 36864 14924 36916
rect 14976 36904 14982 36916
rect 20070 36904 20076 36916
rect 14976 36876 20076 36904
rect 14976 36864 14982 36876
rect 20070 36864 20076 36876
rect 20128 36864 20134 36916
rect 20165 36907 20223 36913
rect 20165 36873 20177 36907
rect 20211 36904 20223 36907
rect 20622 36904 20628 36916
rect 20211 36876 20628 36904
rect 20211 36873 20223 36876
rect 20165 36867 20223 36873
rect 20622 36864 20628 36876
rect 20680 36864 20686 36916
rect 20809 36907 20867 36913
rect 20809 36873 20821 36907
rect 20855 36904 20867 36907
rect 20990 36904 20996 36916
rect 20855 36876 20996 36904
rect 20855 36873 20867 36876
rect 20809 36867 20867 36873
rect 20990 36864 20996 36876
rect 21048 36864 21054 36916
rect 21910 36864 21916 36916
rect 21968 36904 21974 36916
rect 22005 36907 22063 36913
rect 22005 36904 22017 36907
rect 21968 36876 22017 36904
rect 21968 36864 21974 36876
rect 22005 36873 22017 36876
rect 22051 36873 22063 36907
rect 22646 36904 22652 36916
rect 22607 36876 22652 36904
rect 22005 36867 22063 36873
rect 22646 36864 22652 36876
rect 22704 36864 22710 36916
rect 23308 36876 25176 36904
rect 16758 36836 16764 36848
rect 14214 36808 16252 36836
rect 14921 36771 14979 36777
rect 14921 36737 14933 36771
rect 14967 36737 14979 36771
rect 14921 36731 14979 36737
rect 12434 36660 12440 36712
rect 12492 36700 12498 36712
rect 12713 36703 12771 36709
rect 12713 36700 12725 36703
rect 12492 36672 12725 36700
rect 12492 36660 12498 36672
rect 12713 36669 12725 36672
rect 12759 36669 12771 36703
rect 12986 36700 12992 36712
rect 12947 36672 12992 36700
rect 12713 36663 12771 36669
rect 12986 36660 12992 36672
rect 13044 36660 13050 36712
rect 14936 36700 14964 36731
rect 14016 36672 14964 36700
rect 16224 36700 16252 36808
rect 16316 36808 16764 36836
rect 16316 36777 16344 36808
rect 16758 36796 16764 36808
rect 16816 36796 16822 36848
rect 17402 36836 17408 36848
rect 16868 36808 17408 36836
rect 16301 36771 16359 36777
rect 16301 36737 16313 36771
rect 16347 36737 16359 36771
rect 16868 36768 16896 36808
rect 17402 36796 17408 36808
rect 17460 36796 17466 36848
rect 18414 36796 18420 36848
rect 18472 36836 18478 36848
rect 23308 36836 23336 36876
rect 24210 36836 24216 36848
rect 18472 36808 23336 36836
rect 24171 36808 24216 36836
rect 18472 36796 18478 36808
rect 16301 36731 16359 36737
rect 16684 36740 16896 36768
rect 16684 36700 16712 36740
rect 18230 36728 18236 36780
rect 18288 36728 18294 36780
rect 19334 36728 19340 36780
rect 19392 36768 19398 36780
rect 19429 36771 19487 36777
rect 19429 36768 19441 36771
rect 19392 36740 19441 36768
rect 19392 36728 19398 36740
rect 19429 36737 19441 36740
rect 19475 36737 19487 36771
rect 20070 36768 20076 36780
rect 20031 36740 20076 36768
rect 19429 36731 19487 36737
rect 20070 36728 20076 36740
rect 20128 36728 20134 36780
rect 20714 36768 20720 36780
rect 20675 36740 20720 36768
rect 20714 36728 20720 36740
rect 20772 36728 20778 36780
rect 22189 36771 22247 36777
rect 22189 36737 22201 36771
rect 22235 36768 22247 36771
rect 22278 36768 22284 36780
rect 22235 36740 22284 36768
rect 22235 36737 22247 36740
rect 22189 36731 22247 36737
rect 22278 36728 22284 36740
rect 22336 36728 22342 36780
rect 22738 36728 22744 36780
rect 22796 36768 22802 36780
rect 22833 36771 22891 36777
rect 22833 36768 22845 36771
rect 22796 36740 22845 36768
rect 22796 36728 22802 36740
rect 22833 36737 22845 36740
rect 22879 36768 22891 36771
rect 23198 36768 23204 36780
rect 22879 36740 23204 36768
rect 22879 36737 22891 36740
rect 22833 36731 22891 36737
rect 23198 36728 23204 36740
rect 23256 36728 23262 36780
rect 23308 36777 23336 36808
rect 24210 36796 24216 36808
rect 24268 36796 24274 36848
rect 25148 36836 25176 36876
rect 25222 36864 25228 36916
rect 25280 36904 25286 36916
rect 26602 36904 26608 36916
rect 25280 36876 26608 36904
rect 25280 36864 25286 36876
rect 26602 36864 26608 36876
rect 26660 36864 26666 36916
rect 27157 36907 27215 36913
rect 27157 36873 27169 36907
rect 27203 36904 27215 36907
rect 27798 36904 27804 36916
rect 27203 36876 27804 36904
rect 27203 36873 27215 36876
rect 27157 36867 27215 36873
rect 27798 36864 27804 36876
rect 27856 36864 27862 36916
rect 27890 36864 27896 36916
rect 27948 36904 27954 36916
rect 27948 36876 30413 36904
rect 27948 36864 27954 36876
rect 25148 36808 27384 36836
rect 23293 36771 23351 36777
rect 23293 36737 23305 36771
rect 23339 36737 23351 36771
rect 25866 36768 25872 36780
rect 25827 36740 25872 36768
rect 23293 36731 23351 36737
rect 25866 36728 25872 36740
rect 25924 36728 25930 36780
rect 26326 36768 26332 36780
rect 26287 36740 26332 36768
rect 26326 36728 26332 36740
rect 26384 36728 26390 36780
rect 26602 36768 26608 36780
rect 26436 36740 26608 36768
rect 16224 36672 16712 36700
rect 12084 36604 12848 36632
rect 1581 36567 1639 36573
rect 1581 36533 1593 36567
rect 1627 36564 1639 36567
rect 1854 36564 1860 36576
rect 1627 36536 1860 36564
rect 1627 36533 1639 36536
rect 1581 36527 1639 36533
rect 1854 36524 1860 36536
rect 1912 36524 1918 36576
rect 2682 36564 2688 36576
rect 2643 36536 2688 36564
rect 2682 36524 2688 36536
rect 2740 36524 2746 36576
rect 4801 36567 4859 36573
rect 4801 36533 4813 36567
rect 4847 36564 4859 36567
rect 6454 36564 6460 36576
rect 4847 36536 6460 36564
rect 4847 36533 4859 36536
rect 4801 36527 4859 36533
rect 6454 36524 6460 36536
rect 6512 36524 6518 36576
rect 7742 36564 7748 36576
rect 7703 36536 7748 36564
rect 7742 36524 7748 36536
rect 7800 36524 7806 36576
rect 9122 36564 9128 36576
rect 9083 36536 9128 36564
rect 9122 36524 9128 36536
rect 9180 36524 9186 36576
rect 10318 36564 10324 36576
rect 10279 36536 10324 36564
rect 10318 36524 10324 36536
rect 10376 36524 10382 36576
rect 12820 36564 12848 36604
rect 14016 36564 14044 36672
rect 16758 36660 16764 36712
rect 16816 36700 16822 36712
rect 16853 36703 16911 36709
rect 16853 36700 16865 36703
rect 16816 36672 16865 36700
rect 16816 36660 16822 36672
rect 16853 36669 16865 36672
rect 16899 36669 16911 36703
rect 17129 36703 17187 36709
rect 17129 36700 17141 36703
rect 16853 36663 16911 36669
rect 16960 36672 17141 36700
rect 14461 36635 14519 36641
rect 14461 36601 14473 36635
rect 14507 36632 14519 36635
rect 16574 36632 16580 36644
rect 14507 36604 16580 36632
rect 14507 36601 14519 36604
rect 14461 36595 14519 36601
rect 16574 36592 16580 36604
rect 16632 36592 16638 36644
rect 16666 36592 16672 36644
rect 16724 36632 16730 36644
rect 16960 36632 16988 36672
rect 17129 36669 17141 36672
rect 17175 36669 17187 36703
rect 17129 36663 17187 36669
rect 17218 36660 17224 36712
rect 17276 36700 17282 36712
rect 19242 36700 19248 36712
rect 17276 36672 19248 36700
rect 17276 36660 17282 36672
rect 19242 36660 19248 36672
rect 19300 36660 19306 36712
rect 19521 36703 19579 36709
rect 19521 36669 19533 36703
rect 19567 36700 19579 36703
rect 20530 36700 20536 36712
rect 19567 36672 20536 36700
rect 19567 36669 19579 36672
rect 19521 36663 19579 36669
rect 20530 36660 20536 36672
rect 20588 36660 20594 36712
rect 23385 36703 23443 36709
rect 23385 36669 23397 36703
rect 23431 36700 23443 36703
rect 23934 36700 23940 36712
rect 23431 36672 23940 36700
rect 23431 36669 23443 36672
rect 23385 36663 23443 36669
rect 23934 36660 23940 36672
rect 23992 36660 23998 36712
rect 24026 36660 24032 36712
rect 24084 36700 24090 36712
rect 24084 36688 26280 36700
rect 26436 36688 26464 36740
rect 26602 36728 26608 36740
rect 26660 36768 26666 36780
rect 27246 36768 27252 36780
rect 26660 36740 27252 36768
rect 26660 36728 26666 36740
rect 27246 36728 27252 36740
rect 27304 36728 27310 36780
rect 27356 36777 27384 36808
rect 27430 36796 27436 36848
rect 27488 36836 27494 36848
rect 30282 36836 30288 36848
rect 27488 36808 30288 36836
rect 27488 36796 27494 36808
rect 30282 36796 30288 36808
rect 30340 36796 30346 36848
rect 30385 36845 30413 36876
rect 32214 36864 32220 36916
rect 32272 36904 32278 36916
rect 33229 36907 33287 36913
rect 33229 36904 33241 36907
rect 32272 36876 33241 36904
rect 32272 36864 32278 36876
rect 33229 36873 33241 36876
rect 33275 36873 33287 36907
rect 33229 36867 33287 36873
rect 30377 36839 30435 36845
rect 30377 36805 30389 36839
rect 30423 36805 30435 36839
rect 38102 36836 38108 36848
rect 38063 36808 38108 36836
rect 30377 36799 30435 36805
rect 38102 36796 38108 36808
rect 38160 36796 38166 36848
rect 27341 36771 27399 36777
rect 27341 36737 27353 36771
rect 27387 36737 27399 36771
rect 27341 36731 27399 36737
rect 32401 36771 32459 36777
rect 32401 36737 32413 36771
rect 32447 36737 32459 36771
rect 33042 36768 33048 36780
rect 33003 36740 33048 36768
rect 32401 36731 32459 36737
rect 27706 36700 27712 36712
rect 24084 36672 26464 36688
rect 24084 36660 24090 36672
rect 26252 36660 26464 36672
rect 26528 36672 27712 36700
rect 16724 36604 16988 36632
rect 16724 36592 16730 36604
rect 18138 36592 18144 36644
rect 18196 36632 18202 36644
rect 22094 36632 22100 36644
rect 18196 36604 22100 36632
rect 18196 36592 18202 36604
rect 22094 36592 22100 36604
rect 22152 36592 22158 36644
rect 22186 36592 22192 36644
rect 22244 36632 22250 36644
rect 25866 36632 25872 36644
rect 22244 36604 25872 36632
rect 22244 36592 22250 36604
rect 25866 36592 25872 36604
rect 25924 36592 25930 36644
rect 26528 36632 26556 36672
rect 27706 36660 27712 36672
rect 27764 36660 27770 36712
rect 27798 36660 27804 36712
rect 27856 36700 27862 36712
rect 27893 36703 27951 36709
rect 27893 36700 27905 36703
rect 27856 36672 27905 36700
rect 27856 36660 27862 36672
rect 27893 36669 27905 36672
rect 27939 36669 27951 36703
rect 28074 36700 28080 36712
rect 28035 36672 28080 36700
rect 27893 36663 27951 36669
rect 28074 36660 28080 36672
rect 28132 36660 28138 36712
rect 28994 36700 29000 36712
rect 28955 36672 29000 36700
rect 28994 36660 29000 36672
rect 29052 36660 29058 36712
rect 29086 36660 29092 36712
rect 29144 36700 29150 36712
rect 30285 36703 30343 36709
rect 30285 36700 30297 36703
rect 29144 36672 30297 36700
rect 29144 36660 29150 36672
rect 30285 36669 30297 36672
rect 30331 36669 30343 36703
rect 30285 36663 30343 36669
rect 30374 36660 30380 36712
rect 30432 36700 30438 36712
rect 30561 36703 30619 36709
rect 30561 36700 30573 36703
rect 30432 36672 30573 36700
rect 30432 36660 30438 36672
rect 30561 36669 30573 36672
rect 30607 36669 30619 36703
rect 30561 36663 30619 36669
rect 26252 36604 26556 36632
rect 15010 36564 15016 36576
rect 12820 36536 14044 36564
rect 14971 36536 15016 36564
rect 15010 36524 15016 36536
rect 15068 36524 15074 36576
rect 16117 36567 16175 36573
rect 16117 36533 16129 36567
rect 16163 36564 16175 36567
rect 16942 36564 16948 36576
rect 16163 36536 16948 36564
rect 16163 36533 16175 36536
rect 16117 36527 16175 36533
rect 16942 36524 16948 36536
rect 17000 36524 17006 36576
rect 17126 36524 17132 36576
rect 17184 36564 17190 36576
rect 17862 36564 17868 36576
rect 17184 36536 17868 36564
rect 17184 36524 17190 36536
rect 17862 36524 17868 36536
rect 17920 36564 17926 36576
rect 18601 36567 18659 36573
rect 18601 36564 18613 36567
rect 17920 36536 18613 36564
rect 17920 36524 17926 36536
rect 18601 36533 18613 36536
rect 18647 36533 18659 36567
rect 18601 36527 18659 36533
rect 20254 36524 20260 36576
rect 20312 36564 20318 36576
rect 21910 36564 21916 36576
rect 20312 36536 21916 36564
rect 20312 36524 20318 36536
rect 21910 36524 21916 36536
rect 21968 36524 21974 36576
rect 22002 36524 22008 36576
rect 22060 36564 22066 36576
rect 26252 36564 26280 36604
rect 26694 36592 26700 36644
rect 26752 36632 26758 36644
rect 32416 36632 32444 36731
rect 33042 36728 33048 36740
rect 33100 36728 33106 36780
rect 35434 36728 35440 36780
rect 35492 36768 35498 36780
rect 35713 36771 35771 36777
rect 35713 36768 35725 36771
rect 35492 36740 35725 36768
rect 35492 36728 35498 36740
rect 35713 36737 35725 36740
rect 35759 36737 35771 36771
rect 35713 36731 35771 36737
rect 36909 36771 36967 36777
rect 36909 36737 36921 36771
rect 36955 36768 36967 36771
rect 39298 36768 39304 36780
rect 36955 36740 39304 36768
rect 36955 36737 36967 36740
rect 36909 36731 36967 36737
rect 39298 36728 39304 36740
rect 39356 36728 39362 36780
rect 26752 36604 32444 36632
rect 26752 36592 26758 36604
rect 32674 36592 32680 36644
rect 32732 36632 32738 36644
rect 35529 36635 35587 36641
rect 35529 36632 35541 36635
rect 32732 36604 35541 36632
rect 32732 36592 32738 36604
rect 35529 36601 35541 36604
rect 35575 36601 35587 36635
rect 35529 36595 35587 36601
rect 26418 36564 26424 36576
rect 22060 36536 26280 36564
rect 26379 36536 26424 36564
rect 22060 36524 22066 36536
rect 26418 36524 26424 36536
rect 26476 36524 26482 36576
rect 27338 36524 27344 36576
rect 27396 36564 27402 36576
rect 28626 36564 28632 36576
rect 27396 36536 28632 36564
rect 27396 36524 27402 36536
rect 28626 36524 28632 36536
rect 28684 36524 28690 36576
rect 32490 36564 32496 36576
rect 32451 36536 32496 36564
rect 32490 36524 32496 36536
rect 32548 36524 32554 36576
rect 36722 36564 36728 36576
rect 36683 36536 36728 36564
rect 36722 36524 36728 36536
rect 36780 36524 36786 36576
rect 37274 36524 37280 36576
rect 37332 36564 37338 36576
rect 38197 36567 38255 36573
rect 38197 36564 38209 36567
rect 37332 36536 38209 36564
rect 37332 36524 37338 36536
rect 38197 36533 38209 36536
rect 38243 36533 38255 36567
rect 38197 36527 38255 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 2225 36363 2283 36369
rect 2225 36329 2237 36363
rect 2271 36360 2283 36363
rect 4706 36360 4712 36372
rect 2271 36332 4712 36360
rect 2271 36329 2283 36332
rect 2225 36323 2283 36329
rect 4706 36320 4712 36332
rect 4764 36320 4770 36372
rect 8481 36363 8539 36369
rect 8481 36329 8493 36363
rect 8527 36360 8539 36363
rect 8662 36360 8668 36372
rect 8527 36332 8668 36360
rect 8527 36329 8539 36332
rect 8481 36323 8539 36329
rect 8662 36320 8668 36332
rect 8720 36320 8726 36372
rect 13633 36363 13691 36369
rect 13633 36360 13645 36363
rect 8864 36332 13645 36360
rect 1581 36295 1639 36301
rect 1581 36261 1593 36295
rect 1627 36292 1639 36295
rect 7650 36292 7656 36304
rect 1627 36264 7656 36292
rect 1627 36261 1639 36264
rect 1581 36255 1639 36261
rect 7650 36252 7656 36264
rect 7708 36252 7714 36304
rect 8110 36252 8116 36304
rect 8168 36292 8174 36304
rect 8864 36292 8892 36332
rect 13633 36329 13645 36332
rect 13679 36329 13691 36363
rect 13633 36323 13691 36329
rect 13998 36320 14004 36372
rect 14056 36360 14062 36372
rect 18414 36360 18420 36372
rect 14056 36332 18420 36360
rect 14056 36320 14062 36332
rect 18414 36320 18420 36332
rect 18472 36320 18478 36372
rect 18782 36320 18788 36372
rect 18840 36360 18846 36372
rect 20530 36360 20536 36372
rect 18840 36332 20536 36360
rect 18840 36320 18846 36332
rect 20530 36320 20536 36332
rect 20588 36320 20594 36372
rect 20806 36320 20812 36372
rect 20864 36360 20870 36372
rect 21634 36360 21640 36372
rect 20864 36332 21640 36360
rect 20864 36320 20870 36332
rect 21634 36320 21640 36332
rect 21692 36320 21698 36372
rect 22646 36320 22652 36372
rect 22704 36360 22710 36372
rect 33042 36360 33048 36372
rect 22704 36332 33048 36360
rect 22704 36320 22710 36332
rect 33042 36320 33048 36332
rect 33100 36320 33106 36372
rect 37182 36320 37188 36372
rect 37240 36360 37246 36372
rect 37461 36363 37519 36369
rect 37461 36360 37473 36363
rect 37240 36332 37473 36360
rect 37240 36320 37246 36332
rect 37461 36329 37473 36332
rect 37507 36329 37519 36363
rect 37461 36323 37519 36329
rect 8168 36264 8892 36292
rect 8168 36252 8174 36264
rect 9122 36252 9128 36304
rect 9180 36292 9186 36304
rect 10781 36295 10839 36301
rect 10781 36292 10793 36295
rect 9180 36264 10793 36292
rect 9180 36252 9186 36264
rect 10781 36261 10793 36264
rect 10827 36261 10839 36295
rect 12894 36292 12900 36304
rect 10781 36255 10839 36261
rect 11624 36264 12900 36292
rect 6454 36224 6460 36236
rect 6415 36196 6460 36224
rect 6454 36184 6460 36196
rect 6512 36184 6518 36236
rect 9582 36224 9588 36236
rect 8404 36196 9588 36224
rect 14 36116 20 36168
rect 72 36156 78 36168
rect 1765 36159 1823 36165
rect 1765 36156 1777 36159
rect 72 36128 1777 36156
rect 72 36116 78 36128
rect 1765 36125 1777 36128
rect 1811 36125 1823 36159
rect 1765 36119 1823 36125
rect 2409 36159 2467 36165
rect 2409 36125 2421 36159
rect 2455 36156 2467 36159
rect 2866 36156 2872 36168
rect 2455 36128 2872 36156
rect 2455 36125 2467 36128
rect 2409 36119 2467 36125
rect 2866 36116 2872 36128
rect 2924 36116 2930 36168
rect 8404 36165 8432 36196
rect 9582 36184 9588 36196
rect 9640 36184 9646 36236
rect 9769 36227 9827 36233
rect 9769 36193 9781 36227
rect 9815 36224 9827 36227
rect 9876 36224 10088 36236
rect 10226 36224 10232 36236
rect 9815 36208 10232 36224
rect 9815 36196 9904 36208
rect 10060 36196 10232 36208
rect 9815 36193 9827 36196
rect 9769 36187 9827 36193
rect 10226 36184 10232 36196
rect 10284 36184 10290 36236
rect 10410 36224 10416 36236
rect 10371 36196 10416 36224
rect 10410 36184 10416 36196
rect 10468 36184 10474 36236
rect 8389 36159 8447 36165
rect 8389 36156 8401 36159
rect 7392 36128 8401 36156
rect 6546 36088 6552 36100
rect 6507 36060 6552 36088
rect 6546 36048 6552 36060
rect 6604 36048 6610 36100
rect 6822 36048 6828 36100
rect 6880 36088 6886 36100
rect 7392 36088 7420 36128
rect 8389 36125 8401 36128
rect 8435 36125 8447 36159
rect 8389 36119 8447 36125
rect 10597 36159 10655 36165
rect 10597 36125 10609 36159
rect 10643 36156 10655 36159
rect 10870 36156 10876 36168
rect 10643 36128 10876 36156
rect 10643 36125 10655 36128
rect 10597 36119 10655 36125
rect 10870 36116 10876 36128
rect 10928 36116 10934 36168
rect 11624 36156 11652 36264
rect 12894 36252 12900 36264
rect 12952 36252 12958 36304
rect 12986 36252 12992 36304
rect 13044 36292 13050 36304
rect 16390 36292 16396 36304
rect 13044 36264 16396 36292
rect 13044 36252 13050 36264
rect 16390 36252 16396 36264
rect 16448 36252 16454 36304
rect 18230 36252 18236 36304
rect 18288 36292 18294 36304
rect 18288 36264 21220 36292
rect 18288 36252 18294 36264
rect 11974 36184 11980 36236
rect 12032 36224 12038 36236
rect 12032 36196 14504 36224
rect 12032 36184 12038 36196
rect 11701 36159 11759 36165
rect 11701 36156 11713 36159
rect 11624 36128 11713 36156
rect 11701 36125 11713 36128
rect 11747 36125 11759 36159
rect 11701 36119 11759 36125
rect 6880 36060 7420 36088
rect 7469 36091 7527 36097
rect 6880 36048 6886 36060
rect 7469 36057 7481 36091
rect 7515 36057 7527 36091
rect 7469 36051 7527 36057
rect 7484 36020 7512 36051
rect 9122 36048 9128 36100
rect 9180 36088 9186 36100
rect 9309 36091 9367 36097
rect 9309 36088 9321 36091
rect 9180 36060 9321 36088
rect 9180 36048 9186 36060
rect 9309 36057 9321 36060
rect 9355 36057 9367 36091
rect 9309 36051 9367 36057
rect 9401 36091 9459 36097
rect 9401 36057 9413 36091
rect 9447 36088 9459 36091
rect 9766 36088 9772 36100
rect 9447 36060 9772 36088
rect 9447 36057 9459 36060
rect 9401 36051 9459 36057
rect 9766 36048 9772 36060
rect 9824 36048 9830 36100
rect 9950 36048 9956 36100
rect 10008 36088 10014 36100
rect 11716 36088 11744 36119
rect 11882 36116 11888 36168
rect 11940 36156 11946 36168
rect 12897 36159 12955 36165
rect 12897 36156 12909 36159
rect 11940 36128 12909 36156
rect 11940 36116 11946 36128
rect 12897 36125 12909 36128
rect 12943 36156 12955 36159
rect 13538 36156 13544 36168
rect 12943 36128 13544 36156
rect 12943 36125 12955 36128
rect 12897 36119 12955 36125
rect 13538 36116 13544 36128
rect 13596 36116 13602 36168
rect 14476 36158 14504 36196
rect 15562 36184 15568 36236
rect 15620 36224 15626 36236
rect 20254 36224 20260 36236
rect 15620 36196 20260 36224
rect 15620 36184 15626 36196
rect 20254 36184 20260 36196
rect 20312 36184 20318 36236
rect 20441 36227 20499 36233
rect 20441 36193 20453 36227
rect 20487 36224 20499 36227
rect 21082 36224 21088 36236
rect 20487 36196 21088 36224
rect 20487 36193 20499 36196
rect 20441 36187 20499 36193
rect 21082 36184 21088 36196
rect 21140 36184 21146 36236
rect 14553 36159 14611 36165
rect 14553 36158 14565 36159
rect 14476 36130 14565 36158
rect 14553 36125 14565 36130
rect 14599 36125 14611 36159
rect 16758 36156 16764 36168
rect 16719 36128 16764 36156
rect 14553 36119 14611 36125
rect 16758 36116 16764 36128
rect 16816 36116 16822 36168
rect 18138 36116 18144 36168
rect 18196 36116 18202 36168
rect 18322 36116 18328 36168
rect 18380 36156 18386 36168
rect 18380 36128 19656 36156
rect 18380 36116 18386 36128
rect 14642 36088 14648 36100
rect 10008 36060 11744 36088
rect 14603 36060 14648 36088
rect 10008 36048 10014 36060
rect 14642 36048 14648 36060
rect 14700 36048 14706 36100
rect 15562 36048 15568 36100
rect 15620 36088 15626 36100
rect 17037 36091 17095 36097
rect 17037 36088 17049 36091
rect 15620 36060 17049 36088
rect 15620 36048 15626 36060
rect 17037 36057 17049 36060
rect 17083 36057 17095 36091
rect 19426 36088 19432 36100
rect 17037 36051 17095 36057
rect 18432 36060 19432 36088
rect 11054 36020 11060 36032
rect 7484 35992 11060 36020
rect 11054 35980 11060 35992
rect 11112 35980 11118 36032
rect 11514 36020 11520 36032
rect 11475 35992 11520 36020
rect 11514 35980 11520 35992
rect 11572 35980 11578 36032
rect 11606 35980 11612 36032
rect 11664 36020 11670 36032
rect 12989 36023 13047 36029
rect 12989 36020 13001 36023
rect 11664 35992 13001 36020
rect 11664 35980 11670 35992
rect 12989 35989 13001 35992
rect 13035 35989 13047 36023
rect 12989 35983 13047 35989
rect 14274 35980 14280 36032
rect 14332 36020 14338 36032
rect 18432 36020 18460 36060
rect 19426 36048 19432 36060
rect 19484 36048 19490 36100
rect 19628 36088 19656 36128
rect 19702 36116 19708 36168
rect 19760 36156 19766 36168
rect 20070 36156 20076 36168
rect 19760 36128 20076 36156
rect 19760 36116 19766 36128
rect 20070 36116 20076 36128
rect 20128 36116 20134 36168
rect 20162 36088 20168 36100
rect 19628 36060 20168 36088
rect 20162 36048 20168 36060
rect 20220 36048 20226 36100
rect 20530 36048 20536 36100
rect 20588 36088 20594 36100
rect 20588 36060 20633 36088
rect 20588 36048 20594 36060
rect 20898 36048 20904 36100
rect 20956 36088 20962 36100
rect 21085 36091 21143 36097
rect 21085 36088 21097 36091
rect 20956 36060 21097 36088
rect 20956 36048 20962 36060
rect 21085 36057 21097 36060
rect 21131 36057 21143 36091
rect 21192 36088 21220 36264
rect 26694 36252 26700 36304
rect 26752 36292 26758 36304
rect 26973 36295 27031 36301
rect 26973 36292 26985 36295
rect 26752 36264 26985 36292
rect 26752 36252 26758 36264
rect 26973 36261 26985 36264
rect 27019 36261 27031 36295
rect 26973 36255 27031 36261
rect 27430 36252 27436 36304
rect 27488 36292 27494 36304
rect 31665 36295 31723 36301
rect 31665 36292 31677 36295
rect 27488 36264 31677 36292
rect 27488 36252 27494 36264
rect 31665 36261 31677 36264
rect 31711 36261 31723 36295
rect 31665 36255 31723 36261
rect 22189 36227 22247 36233
rect 22189 36193 22201 36227
rect 22235 36224 22247 36227
rect 22235 36196 23888 36224
rect 22235 36193 22247 36196
rect 22189 36187 22247 36193
rect 23382 36156 23388 36168
rect 23032 36128 23388 36156
rect 22281 36091 22339 36097
rect 21192 36060 22232 36088
rect 21085 36051 21143 36057
rect 14332 35992 18460 36020
rect 14332 35980 14338 35992
rect 18506 35980 18512 36032
rect 18564 36020 18570 36032
rect 18564 35992 18609 36020
rect 18564 35980 18570 35992
rect 18690 35980 18696 36032
rect 18748 36020 18754 36032
rect 19702 36020 19708 36032
rect 18748 35992 19708 36020
rect 18748 35980 18754 35992
rect 19702 35980 19708 35992
rect 19760 35980 19766 36032
rect 19797 36023 19855 36029
rect 19797 35989 19809 36023
rect 19843 36020 19855 36023
rect 22094 36020 22100 36032
rect 19843 35992 22100 36020
rect 19843 35989 19855 35992
rect 19797 35983 19855 35989
rect 22094 35980 22100 35992
rect 22152 35980 22158 36032
rect 22204 36020 22232 36060
rect 22281 36057 22293 36091
rect 22327 36088 22339 36091
rect 23032 36088 23060 36128
rect 23382 36116 23388 36128
rect 23440 36116 23446 36168
rect 23474 36116 23480 36168
rect 23532 36156 23538 36168
rect 23661 36159 23719 36165
rect 23661 36156 23673 36159
rect 23532 36128 23673 36156
rect 23532 36116 23538 36128
rect 23661 36125 23673 36128
rect 23707 36125 23719 36159
rect 23860 36156 23888 36196
rect 25130 36184 25136 36236
rect 25188 36224 25194 36236
rect 25188 36196 27200 36224
rect 25188 36184 25194 36196
rect 27172 36165 27200 36196
rect 27246 36184 27252 36236
rect 27304 36224 27310 36236
rect 28353 36227 28411 36233
rect 28353 36224 28365 36227
rect 27304 36196 28365 36224
rect 27304 36184 27310 36196
rect 28353 36193 28365 36196
rect 28399 36193 28411 36227
rect 28353 36187 28411 36193
rect 30193 36227 30251 36233
rect 30193 36193 30205 36227
rect 30239 36224 30251 36227
rect 32401 36227 32459 36233
rect 32401 36224 32413 36227
rect 30239 36196 32413 36224
rect 30239 36193 30251 36196
rect 30193 36187 30251 36193
rect 32401 36193 32413 36196
rect 32447 36193 32459 36227
rect 38654 36224 38660 36236
rect 32401 36187 32459 36193
rect 36832 36196 38660 36224
rect 27157 36159 27215 36165
rect 23860 36128 24532 36156
rect 23661 36119 23719 36125
rect 22327 36060 23060 36088
rect 23201 36091 23259 36097
rect 22327 36057 22339 36060
rect 22281 36051 22339 36057
rect 23201 36057 23213 36091
rect 23247 36088 23259 36091
rect 24026 36088 24032 36100
rect 23247 36060 24032 36088
rect 23247 36057 23259 36060
rect 23201 36051 23259 36057
rect 24026 36048 24032 36060
rect 24084 36048 24090 36100
rect 23753 36023 23811 36029
rect 23753 36020 23765 36023
rect 22204 35992 23765 36020
rect 23753 35989 23765 35992
rect 23799 35989 23811 36023
rect 24504 36020 24532 36128
rect 27157 36125 27169 36159
rect 27203 36125 27215 36159
rect 31846 36156 31852 36168
rect 31807 36128 31852 36156
rect 27157 36119 27215 36125
rect 31846 36116 31852 36128
rect 31904 36116 31910 36168
rect 32306 36156 32312 36168
rect 32267 36128 32312 36156
rect 32306 36116 32312 36128
rect 32364 36116 32370 36168
rect 36832 36165 36860 36196
rect 38654 36184 38660 36196
rect 38712 36184 38718 36236
rect 36817 36159 36875 36165
rect 36817 36125 36829 36159
rect 36863 36125 36875 36159
rect 36817 36119 36875 36125
rect 37277 36159 37335 36165
rect 37277 36125 37289 36159
rect 37323 36125 37335 36159
rect 37277 36119 37335 36125
rect 24670 36088 24676 36100
rect 24631 36060 24676 36088
rect 24670 36048 24676 36060
rect 24728 36048 24734 36100
rect 24762 36048 24768 36100
rect 24820 36088 24826 36100
rect 25317 36091 25375 36097
rect 24820 36060 24865 36088
rect 24820 36048 24826 36060
rect 25317 36057 25329 36091
rect 25363 36088 25375 36091
rect 25498 36088 25504 36100
rect 25363 36060 25504 36088
rect 25363 36057 25375 36060
rect 25317 36051 25375 36057
rect 25498 36048 25504 36060
rect 25556 36048 25562 36100
rect 25869 36091 25927 36097
rect 25869 36057 25881 36091
rect 25915 36057 25927 36091
rect 25869 36051 25927 36057
rect 25884 36020 25912 36051
rect 25958 36048 25964 36100
rect 26016 36088 26022 36100
rect 26016 36060 26061 36088
rect 26016 36048 26022 36060
rect 26234 36048 26240 36100
rect 26292 36088 26298 36100
rect 26513 36091 26571 36097
rect 26513 36088 26525 36091
rect 26292 36060 26525 36088
rect 26292 36048 26298 36060
rect 26513 36057 26525 36060
rect 26559 36088 26571 36091
rect 27062 36088 27068 36100
rect 26559 36060 27068 36088
rect 26559 36057 26571 36060
rect 26513 36051 26571 36057
rect 27062 36048 27068 36060
rect 27120 36048 27126 36100
rect 28074 36088 28080 36100
rect 28035 36060 28080 36088
rect 28074 36048 28080 36060
rect 28132 36048 28138 36100
rect 28169 36091 28227 36097
rect 28169 36057 28181 36091
rect 28215 36088 28227 36091
rect 28994 36088 29000 36100
rect 28215 36060 29000 36088
rect 28215 36057 28227 36060
rect 28169 36051 28227 36057
rect 28994 36048 29000 36060
rect 29052 36048 29058 36100
rect 30285 36091 30343 36097
rect 30285 36057 30297 36091
rect 30331 36088 30343 36091
rect 30834 36088 30840 36100
rect 30331 36060 30840 36088
rect 30331 36057 30343 36060
rect 30285 36051 30343 36057
rect 30834 36048 30840 36060
rect 30892 36048 30898 36100
rect 31018 36048 31024 36100
rect 31076 36088 31082 36100
rect 31205 36091 31263 36097
rect 31205 36088 31217 36091
rect 31076 36060 31217 36088
rect 31076 36048 31082 36060
rect 31205 36057 31217 36060
rect 31251 36057 31263 36091
rect 37292 36088 37320 36119
rect 37366 36116 37372 36168
rect 37424 36156 37430 36168
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 37424 36128 38025 36156
rect 37424 36116 37430 36128
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 38378 36088 38384 36100
rect 37292 36060 38384 36088
rect 31205 36051 31263 36057
rect 38378 36048 38384 36060
rect 38436 36048 38442 36100
rect 30374 36020 30380 36032
rect 24504 35992 30380 36020
rect 23753 35983 23811 35989
rect 30374 35980 30380 35992
rect 30432 35980 30438 36032
rect 34514 35980 34520 36032
rect 34572 36020 34578 36032
rect 36633 36023 36691 36029
rect 36633 36020 36645 36023
rect 34572 35992 36645 36020
rect 34572 35980 34578 35992
rect 36633 35989 36645 35992
rect 36679 35989 36691 36023
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 36633 35983 36691 35989
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 10870 35816 10876 35828
rect 10831 35788 10876 35816
rect 10870 35776 10876 35788
rect 10928 35776 10934 35828
rect 16942 35816 16948 35828
rect 12406 35788 16948 35816
rect 9306 35748 9312 35760
rect 9267 35720 9312 35748
rect 9306 35708 9312 35720
rect 9364 35708 9370 35760
rect 12406 35748 12434 35788
rect 16942 35776 16948 35788
rect 17000 35776 17006 35828
rect 20165 35819 20223 35825
rect 20165 35816 20177 35819
rect 17052 35788 20177 35816
rect 17052 35748 17080 35788
rect 20165 35785 20177 35788
rect 20211 35785 20223 35819
rect 20165 35779 20223 35785
rect 20714 35776 20720 35828
rect 20772 35816 20778 35828
rect 20809 35819 20867 35825
rect 20809 35816 20821 35819
rect 20772 35788 20821 35816
rect 20772 35776 20778 35788
rect 20809 35785 20821 35788
rect 20855 35785 20867 35819
rect 20809 35779 20867 35785
rect 20898 35776 20904 35828
rect 20956 35816 20962 35828
rect 21174 35816 21180 35828
rect 20956 35788 21180 35816
rect 20956 35776 20962 35788
rect 21174 35776 21180 35788
rect 21232 35776 21238 35828
rect 22094 35776 22100 35828
rect 22152 35816 22158 35828
rect 23201 35819 23259 35825
rect 23201 35816 23213 35819
rect 22152 35788 23213 35816
rect 22152 35776 22158 35788
rect 23201 35785 23213 35788
rect 23247 35785 23259 35819
rect 23201 35779 23259 35785
rect 24670 35776 24676 35828
rect 24728 35816 24734 35828
rect 25593 35819 25651 35825
rect 25593 35816 25605 35819
rect 24728 35788 25605 35816
rect 24728 35776 24734 35788
rect 25593 35785 25605 35788
rect 25639 35785 25651 35819
rect 25593 35779 25651 35785
rect 25958 35776 25964 35828
rect 26016 35816 26022 35828
rect 26237 35819 26295 35825
rect 26237 35816 26249 35819
rect 26016 35788 26249 35816
rect 26016 35776 26022 35788
rect 26237 35785 26249 35788
rect 26283 35785 26295 35819
rect 26237 35779 26295 35785
rect 27614 35776 27620 35828
rect 27672 35816 27678 35828
rect 27672 35788 30420 35816
rect 27672 35776 27678 35788
rect 21542 35748 21548 35760
rect 9416 35720 12434 35748
rect 13938 35720 17080 35748
rect 18354 35720 21548 35748
rect 1670 35680 1676 35692
rect 1631 35652 1676 35680
rect 1670 35640 1676 35652
rect 1728 35640 1734 35692
rect 2593 35683 2651 35689
rect 2593 35649 2605 35683
rect 2639 35680 2651 35683
rect 3418 35680 3424 35692
rect 2639 35652 3424 35680
rect 2639 35649 2651 35652
rect 2593 35643 2651 35649
rect 3418 35640 3424 35652
rect 3476 35640 3482 35692
rect 3602 35640 3608 35692
rect 3660 35680 3666 35692
rect 9033 35683 9091 35689
rect 9033 35680 9045 35683
rect 3660 35652 9045 35680
rect 3660 35640 3666 35652
rect 9033 35649 9045 35652
rect 9079 35649 9091 35683
rect 9033 35643 9091 35649
rect 4062 35572 4068 35624
rect 4120 35612 4126 35624
rect 9416 35612 9444 35720
rect 21542 35708 21548 35720
rect 21600 35708 21606 35760
rect 22278 35748 22284 35760
rect 22066 35720 22284 35748
rect 11057 35683 11115 35689
rect 11057 35649 11069 35683
rect 11103 35680 11115 35683
rect 11514 35680 11520 35692
rect 11103 35652 11520 35680
rect 11103 35649 11115 35652
rect 11057 35643 11115 35649
rect 11514 35640 11520 35652
rect 11572 35640 11578 35692
rect 19429 35683 19487 35689
rect 19429 35649 19441 35683
rect 19475 35649 19487 35683
rect 19429 35643 19487 35649
rect 4120 35584 9444 35612
rect 4120 35572 4126 35584
rect 12434 35572 12440 35624
rect 12492 35612 12498 35624
rect 12713 35615 12771 35621
rect 12492 35584 12537 35612
rect 12492 35572 12498 35584
rect 12713 35581 12725 35615
rect 12759 35612 12771 35615
rect 12802 35612 12808 35624
rect 12759 35584 12808 35612
rect 12759 35581 12771 35584
rect 12713 35575 12771 35581
rect 12802 35572 12808 35584
rect 12860 35572 12866 35624
rect 14642 35572 14648 35624
rect 14700 35612 14706 35624
rect 16853 35615 16911 35621
rect 16853 35612 16865 35615
rect 14700 35584 16865 35612
rect 14700 35572 14706 35584
rect 16853 35581 16865 35584
rect 16899 35581 16911 35615
rect 16853 35575 16911 35581
rect 17129 35615 17187 35621
rect 17129 35581 17141 35615
rect 17175 35612 17187 35615
rect 17218 35612 17224 35624
rect 17175 35584 17224 35612
rect 17175 35581 17187 35584
rect 17129 35575 17187 35581
rect 17218 35572 17224 35584
rect 17276 35572 17282 35624
rect 17862 35572 17868 35624
rect 17920 35612 17926 35624
rect 19444 35612 19472 35643
rect 19978 35640 19984 35692
rect 20036 35680 20042 35692
rect 20073 35683 20131 35689
rect 20073 35680 20085 35683
rect 20036 35652 20085 35680
rect 20036 35640 20042 35652
rect 20073 35649 20085 35652
rect 20119 35680 20131 35683
rect 20346 35680 20352 35692
rect 20119 35652 20352 35680
rect 20119 35649 20131 35652
rect 20073 35643 20131 35649
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 20714 35680 20720 35692
rect 20675 35652 20720 35680
rect 20714 35640 20720 35652
rect 20772 35640 20778 35692
rect 22066 35680 22094 35720
rect 22278 35708 22284 35720
rect 22336 35708 22342 35760
rect 22462 35708 22468 35760
rect 22520 35748 22526 35760
rect 26418 35748 26424 35760
rect 22520 35720 24348 35748
rect 22520 35708 22526 35720
rect 21192 35652 22094 35680
rect 17920 35584 19472 35612
rect 17920 35572 17926 35584
rect 20162 35572 20168 35624
rect 20220 35612 20226 35624
rect 21192 35612 21220 35652
rect 22186 35640 22192 35692
rect 22244 35680 22250 35692
rect 22244 35652 22289 35680
rect 22244 35640 22250 35652
rect 22370 35640 22376 35692
rect 22428 35680 22434 35692
rect 23109 35683 23167 35689
rect 23109 35680 23121 35683
rect 22428 35652 23121 35680
rect 22428 35640 22434 35652
rect 23109 35649 23121 35652
rect 23155 35649 23167 35683
rect 23109 35643 23167 35649
rect 23474 35640 23480 35692
rect 23532 35680 23538 35692
rect 23753 35683 23811 35689
rect 23753 35680 23765 35683
rect 23532 35652 23765 35680
rect 23532 35640 23538 35652
rect 23753 35649 23765 35652
rect 23799 35649 23811 35683
rect 23753 35643 23811 35649
rect 20220 35584 21220 35612
rect 20220 35572 20226 35584
rect 21266 35572 21272 35624
rect 21324 35612 21330 35624
rect 22005 35615 22063 35621
rect 22005 35612 22017 35615
rect 21324 35584 22017 35612
rect 21324 35572 21330 35584
rect 22005 35581 22017 35584
rect 22051 35581 22063 35615
rect 22005 35575 22063 35581
rect 22094 35572 22100 35624
rect 22152 35612 22158 35624
rect 23845 35615 23903 35621
rect 23845 35612 23857 35615
rect 22152 35584 23857 35612
rect 22152 35572 22158 35584
rect 23845 35581 23857 35584
rect 23891 35581 23903 35615
rect 24320 35612 24348 35720
rect 24412 35720 26424 35748
rect 24412 35689 24440 35720
rect 26418 35708 26424 35720
rect 26476 35708 26482 35760
rect 27706 35748 27712 35760
rect 27080 35720 27712 35748
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35649 24455 35683
rect 24578 35680 24584 35692
rect 24539 35652 24584 35680
rect 24397 35643 24455 35649
rect 24578 35640 24584 35652
rect 24636 35640 24642 35692
rect 25406 35640 25412 35692
rect 25464 35680 25470 35692
rect 25501 35683 25559 35689
rect 25501 35680 25513 35683
rect 25464 35652 25513 35680
rect 25464 35640 25470 35652
rect 25501 35649 25513 35652
rect 25547 35649 25559 35683
rect 25501 35643 25559 35649
rect 25682 35640 25688 35692
rect 25740 35680 25746 35692
rect 26145 35683 26203 35689
rect 26145 35680 26157 35683
rect 25740 35652 26157 35680
rect 25740 35640 25746 35652
rect 26145 35649 26157 35652
rect 26191 35680 26203 35683
rect 27080 35680 27108 35720
rect 27706 35708 27712 35720
rect 27764 35708 27770 35760
rect 27982 35748 27988 35760
rect 27943 35720 27988 35748
rect 27982 35708 27988 35720
rect 28040 35708 28046 35760
rect 29181 35751 29239 35757
rect 29181 35717 29193 35751
rect 29227 35748 29239 35751
rect 29822 35748 29828 35760
rect 29227 35720 29828 35748
rect 29227 35717 29239 35720
rect 29181 35711 29239 35717
rect 29822 35708 29828 35720
rect 29880 35708 29886 35760
rect 26191 35652 27108 35680
rect 26191 35649 26203 35652
rect 26145 35643 26203 35649
rect 27154 35640 27160 35692
rect 27212 35680 27218 35692
rect 30392 35689 30420 35788
rect 30834 35776 30840 35828
rect 30892 35816 30898 35828
rect 30929 35819 30987 35825
rect 30929 35816 30941 35819
rect 30892 35788 30941 35816
rect 30892 35776 30898 35788
rect 30929 35785 30941 35788
rect 30975 35785 30987 35819
rect 30929 35779 30987 35785
rect 30377 35683 30435 35689
rect 27212 35652 27257 35680
rect 27212 35640 27218 35652
rect 30377 35649 30389 35683
rect 30423 35649 30435 35683
rect 30377 35643 30435 35649
rect 30558 35640 30564 35692
rect 30616 35680 30622 35692
rect 30837 35683 30895 35689
rect 30837 35680 30849 35683
rect 30616 35652 30849 35680
rect 30616 35640 30622 35652
rect 30837 35649 30849 35652
rect 30883 35649 30895 35683
rect 30837 35643 30895 35649
rect 32493 35683 32551 35689
rect 32493 35649 32505 35683
rect 32539 35649 32551 35683
rect 32493 35643 32551 35649
rect 26878 35612 26884 35624
rect 24320 35584 26884 35612
rect 23845 35575 23903 35581
rect 26878 35572 26884 35584
rect 26936 35572 26942 35624
rect 27893 35615 27951 35621
rect 27893 35612 27905 35615
rect 26988 35584 27905 35612
rect 14108 35516 16988 35544
rect 1486 35436 1492 35488
rect 1544 35476 1550 35488
rect 1765 35479 1823 35485
rect 1765 35476 1777 35479
rect 1544 35448 1777 35476
rect 1544 35436 1550 35448
rect 1765 35445 1777 35448
rect 1811 35445 1823 35479
rect 1765 35439 1823 35445
rect 2590 35436 2596 35488
rect 2648 35476 2654 35488
rect 2685 35479 2743 35485
rect 2685 35476 2697 35479
rect 2648 35448 2697 35476
rect 2648 35436 2654 35448
rect 2685 35445 2697 35448
rect 2731 35445 2743 35479
rect 2685 35439 2743 35445
rect 3513 35479 3571 35485
rect 3513 35445 3525 35479
rect 3559 35476 3571 35479
rect 3970 35476 3976 35488
rect 3559 35448 3976 35476
rect 3559 35445 3571 35448
rect 3513 35439 3571 35445
rect 3970 35436 3976 35448
rect 4028 35436 4034 35488
rect 7834 35436 7840 35488
rect 7892 35476 7898 35488
rect 12250 35476 12256 35488
rect 7892 35448 12256 35476
rect 7892 35436 7898 35448
rect 12250 35436 12256 35448
rect 12308 35436 12314 35488
rect 12526 35436 12532 35488
rect 12584 35476 12590 35488
rect 14108 35476 14136 35516
rect 12584 35448 14136 35476
rect 12584 35436 12590 35448
rect 14182 35436 14188 35488
rect 14240 35476 14246 35488
rect 16960 35476 16988 35516
rect 18414 35504 18420 35556
rect 18472 35544 18478 35556
rect 18601 35547 18659 35553
rect 18601 35544 18613 35547
rect 18472 35516 18613 35544
rect 18472 35504 18478 35516
rect 18601 35513 18613 35516
rect 18647 35544 18659 35547
rect 19521 35547 19579 35553
rect 18647 35516 19334 35544
rect 18647 35513 18659 35516
rect 18601 35507 18659 35513
rect 18506 35476 18512 35488
rect 14240 35448 14285 35476
rect 16960 35448 18512 35476
rect 14240 35436 14246 35448
rect 18506 35436 18512 35448
rect 18564 35436 18570 35488
rect 19306 35476 19334 35516
rect 19521 35513 19533 35547
rect 19567 35544 19579 35547
rect 20530 35544 20536 35556
rect 19567 35516 20536 35544
rect 19567 35513 19579 35516
rect 19521 35507 19579 35513
rect 20530 35504 20536 35516
rect 20588 35504 20594 35556
rect 22462 35544 22468 35556
rect 22066 35516 22468 35544
rect 20990 35476 20996 35488
rect 19306 35448 20996 35476
rect 20990 35436 20996 35448
rect 21048 35436 21054 35488
rect 21174 35436 21180 35488
rect 21232 35476 21238 35488
rect 22066 35476 22094 35516
rect 22462 35504 22468 35516
rect 22520 35504 22526 35556
rect 22649 35547 22707 35553
rect 22649 35513 22661 35547
rect 22695 35544 22707 35547
rect 25041 35547 25099 35553
rect 25041 35544 25053 35547
rect 22695 35516 25053 35544
rect 22695 35513 22707 35516
rect 22649 35507 22707 35513
rect 25041 35513 25053 35516
rect 25087 35544 25099 35547
rect 26988 35544 27016 35584
rect 27893 35581 27905 35584
rect 27939 35581 27951 35615
rect 28166 35612 28172 35624
rect 28127 35584 28172 35612
rect 27893 35575 27951 35581
rect 28166 35572 28172 35584
rect 28224 35572 28230 35624
rect 28258 35572 28264 35624
rect 28316 35572 28322 35624
rect 29089 35615 29147 35621
rect 29089 35581 29101 35615
rect 29135 35612 29147 35615
rect 31481 35615 31539 35621
rect 31481 35612 31493 35615
rect 29135 35584 31493 35612
rect 29135 35581 29147 35584
rect 29089 35575 29147 35581
rect 31481 35581 31493 35584
rect 31527 35581 31539 35615
rect 32508 35612 32536 35643
rect 37458 35612 37464 35624
rect 31481 35575 31539 35581
rect 31956 35584 32536 35612
rect 37419 35584 37464 35612
rect 25087 35516 27016 35544
rect 25087 35513 25099 35516
rect 25041 35507 25099 35513
rect 27430 35504 27436 35556
rect 27488 35544 27494 35556
rect 28276 35544 28304 35572
rect 29641 35547 29699 35553
rect 29641 35544 29653 35547
rect 27488 35516 28028 35544
rect 28276 35516 29653 35544
rect 27488 35504 27494 35516
rect 21232 35448 22094 35476
rect 21232 35436 21238 35448
rect 22278 35436 22284 35488
rect 22336 35476 22342 35488
rect 27154 35476 27160 35488
rect 22336 35448 27160 35476
rect 22336 35436 22342 35448
rect 27154 35436 27160 35448
rect 27212 35436 27218 35488
rect 27249 35479 27307 35485
rect 27249 35445 27261 35479
rect 27295 35476 27307 35479
rect 27890 35476 27896 35488
rect 27295 35448 27896 35476
rect 27295 35445 27307 35448
rect 27249 35439 27307 35445
rect 27890 35436 27896 35448
rect 27948 35436 27954 35488
rect 28000 35476 28028 35516
rect 29641 35513 29653 35516
rect 29687 35544 29699 35547
rect 30006 35544 30012 35556
rect 29687 35516 30012 35544
rect 29687 35513 29699 35516
rect 29641 35507 29699 35513
rect 30006 35504 30012 35516
rect 30064 35504 30070 35556
rect 30193 35547 30251 35553
rect 30193 35513 30205 35547
rect 30239 35544 30251 35547
rect 31846 35544 31852 35556
rect 30239 35516 31852 35544
rect 30239 35513 30251 35516
rect 30193 35507 30251 35513
rect 31846 35504 31852 35516
rect 31904 35504 31910 35556
rect 29086 35476 29092 35488
rect 28000 35448 29092 35476
rect 29086 35436 29092 35448
rect 29144 35436 29150 35488
rect 29730 35436 29736 35488
rect 29788 35476 29794 35488
rect 31956 35476 31984 35584
rect 37458 35572 37464 35584
rect 37516 35572 37522 35624
rect 37734 35612 37740 35624
rect 37695 35584 37740 35612
rect 37734 35572 37740 35584
rect 37792 35572 37798 35624
rect 29788 35448 31984 35476
rect 29788 35436 29794 35448
rect 32030 35436 32036 35488
rect 32088 35476 32094 35488
rect 32309 35479 32367 35485
rect 32309 35476 32321 35479
rect 32088 35448 32321 35476
rect 32088 35436 32094 35448
rect 32309 35445 32321 35448
rect 32355 35445 32367 35479
rect 32309 35439 32367 35445
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 3142 35232 3148 35284
rect 3200 35272 3206 35284
rect 3329 35275 3387 35281
rect 3329 35272 3341 35275
rect 3200 35244 3341 35272
rect 3200 35232 3206 35244
rect 3329 35241 3341 35244
rect 3375 35272 3387 35275
rect 3602 35272 3608 35284
rect 3375 35244 3608 35272
rect 3375 35241 3387 35244
rect 3329 35235 3387 35241
rect 3602 35232 3608 35244
rect 3660 35232 3666 35284
rect 4062 35272 4068 35284
rect 4023 35244 4068 35272
rect 4062 35232 4068 35244
rect 4120 35232 4126 35284
rect 4890 35232 4896 35284
rect 4948 35272 4954 35284
rect 9582 35272 9588 35284
rect 4948 35244 9588 35272
rect 4948 35232 4954 35244
rect 9582 35232 9588 35244
rect 9640 35232 9646 35284
rect 9766 35232 9772 35284
rect 9824 35272 9830 35284
rect 10321 35275 10379 35281
rect 10321 35272 10333 35275
rect 9824 35244 10333 35272
rect 9824 35232 9830 35244
rect 10321 35241 10333 35244
rect 10367 35241 10379 35275
rect 10321 35235 10379 35241
rect 11228 35275 11286 35281
rect 11228 35241 11240 35275
rect 11274 35272 11286 35275
rect 12526 35272 12532 35284
rect 11274 35244 12532 35272
rect 11274 35241 11286 35244
rect 11228 35235 11286 35241
rect 12526 35232 12532 35244
rect 12584 35232 12590 35284
rect 12713 35275 12771 35281
rect 12713 35241 12725 35275
rect 12759 35272 12771 35275
rect 23753 35275 23811 35281
rect 12759 35244 22094 35272
rect 12759 35241 12771 35244
rect 12713 35235 12771 35241
rect 12250 35164 12256 35216
rect 12308 35204 12314 35216
rect 12728 35204 12756 35235
rect 16390 35204 16396 35216
rect 12308 35176 12756 35204
rect 16351 35176 16396 35204
rect 12308 35164 12314 35176
rect 16390 35164 16396 35176
rect 16448 35164 16454 35216
rect 19334 35204 19340 35216
rect 18156 35176 19340 35204
rect 1857 35139 1915 35145
rect 1857 35105 1869 35139
rect 1903 35136 1915 35139
rect 5350 35136 5356 35148
rect 1903 35108 5356 35136
rect 1903 35105 1915 35108
rect 1857 35099 1915 35105
rect 5350 35096 5356 35108
rect 5408 35096 5414 35148
rect 6273 35139 6331 35145
rect 6273 35105 6285 35139
rect 6319 35136 6331 35139
rect 8202 35136 8208 35148
rect 6319 35108 8208 35136
rect 6319 35105 6331 35108
rect 6273 35099 6331 35105
rect 8202 35096 8208 35108
rect 8260 35096 8266 35148
rect 10965 35139 11023 35145
rect 10965 35105 10977 35139
rect 11011 35136 11023 35139
rect 12434 35136 12440 35148
rect 11011 35108 12440 35136
rect 11011 35105 11023 35108
rect 10965 35099 11023 35105
rect 12434 35096 12440 35108
rect 12492 35136 12498 35148
rect 13170 35136 13176 35148
rect 12492 35108 13176 35136
rect 12492 35096 12498 35108
rect 13170 35096 13176 35108
rect 13228 35096 13234 35148
rect 13354 35136 13360 35148
rect 13315 35108 13360 35136
rect 13354 35096 13360 35108
rect 13412 35096 13418 35148
rect 14642 35136 14648 35148
rect 14603 35108 14648 35136
rect 14642 35096 14648 35108
rect 14700 35096 14706 35148
rect 14921 35139 14979 35145
rect 14921 35105 14933 35139
rect 14967 35136 14979 35139
rect 16482 35136 16488 35148
rect 14967 35108 16488 35136
rect 14967 35105 14979 35108
rect 14921 35099 14979 35105
rect 16482 35096 16488 35108
rect 16540 35096 16546 35148
rect 17126 35136 17132 35148
rect 17087 35108 17132 35136
rect 17126 35096 17132 35108
rect 17184 35096 17190 35148
rect 17494 35096 17500 35148
rect 17552 35136 17558 35148
rect 18156 35136 18184 35176
rect 19334 35164 19340 35176
rect 19392 35164 19398 35216
rect 19978 35164 19984 35216
rect 20036 35204 20042 35216
rect 21818 35204 21824 35216
rect 20036 35176 21824 35204
rect 20036 35164 20042 35176
rect 21818 35164 21824 35176
rect 21876 35164 21882 35216
rect 22066 35204 22094 35244
rect 23753 35241 23765 35275
rect 23799 35272 23811 35275
rect 24762 35272 24768 35284
rect 23799 35244 24768 35272
rect 23799 35241 23811 35244
rect 23753 35235 23811 35241
rect 24762 35232 24768 35244
rect 24820 35232 24826 35284
rect 26510 35232 26516 35284
rect 26568 35272 26574 35284
rect 29914 35272 29920 35284
rect 26568 35244 29920 35272
rect 26568 35232 26574 35244
rect 29914 35232 29920 35244
rect 29972 35232 29978 35284
rect 30466 35272 30472 35284
rect 30427 35244 30472 35272
rect 30466 35232 30472 35244
rect 30524 35232 30530 35284
rect 31021 35275 31079 35281
rect 31021 35241 31033 35275
rect 31067 35272 31079 35275
rect 32306 35272 32312 35284
rect 31067 35244 32312 35272
rect 31067 35241 31079 35244
rect 31021 35235 31079 35241
rect 32306 35232 32312 35244
rect 32364 35232 32370 35284
rect 28074 35204 28080 35216
rect 22066 35176 28080 35204
rect 28074 35164 28080 35176
rect 28132 35164 28138 35216
rect 28350 35164 28356 35216
rect 28408 35164 28414 35216
rect 30006 35164 30012 35216
rect 30064 35204 30070 35216
rect 30064 35176 31754 35204
rect 30064 35164 30070 35176
rect 24673 35139 24731 35145
rect 24673 35136 24685 35139
rect 17552 35108 18184 35136
rect 18248 35108 24685 35136
rect 17552 35096 17558 35108
rect 1581 35071 1639 35077
rect 1581 35037 1593 35071
rect 1627 35037 1639 35071
rect 1581 35031 1639 35037
rect 1596 34932 1624 35031
rect 3326 35028 3332 35080
rect 3384 35068 3390 35080
rect 3973 35071 4031 35077
rect 3973 35068 3985 35071
rect 3384 35040 3985 35068
rect 3384 35028 3390 35040
rect 3973 35037 3985 35040
rect 4019 35037 4031 35071
rect 3973 35031 4031 35037
rect 5997 35071 6055 35077
rect 5997 35037 6009 35071
rect 6043 35037 6055 35071
rect 10502 35068 10508 35080
rect 10463 35040 10508 35068
rect 5997 35031 6055 35037
rect 2590 34960 2596 35012
rect 2648 34960 2654 35012
rect 6012 35000 6040 35031
rect 10502 35028 10508 35040
rect 10560 35028 10566 35080
rect 13262 35068 13268 35080
rect 13223 35040 13268 35068
rect 13262 35028 13268 35040
rect 13320 35028 13326 35080
rect 16850 35068 16856 35080
rect 16811 35040 16856 35068
rect 16850 35028 16856 35040
rect 16908 35028 16914 35080
rect 18248 35054 18276 35108
rect 24673 35105 24685 35108
rect 24719 35105 24731 35139
rect 26234 35136 26240 35148
rect 26147 35108 26240 35136
rect 24673 35099 24731 35105
rect 26234 35096 26240 35108
rect 26292 35136 26298 35148
rect 27430 35136 27436 35148
rect 26292 35108 27436 35136
rect 26292 35096 26298 35108
rect 27430 35096 27436 35108
rect 27488 35096 27494 35148
rect 27801 35139 27859 35145
rect 27801 35136 27813 35139
rect 27540 35108 27813 35136
rect 19426 35068 19432 35080
rect 19387 35040 19432 35068
rect 19426 35028 19432 35040
rect 19484 35028 19490 35080
rect 20162 35068 20168 35080
rect 20123 35040 20168 35068
rect 20162 35028 20168 35040
rect 20220 35028 20226 35080
rect 20254 35028 20260 35080
rect 20312 35068 20318 35080
rect 20714 35068 20720 35080
rect 20312 35040 20720 35068
rect 20312 35028 20318 35040
rect 20714 35028 20720 35040
rect 20772 35068 20778 35080
rect 20809 35071 20867 35077
rect 20809 35068 20821 35071
rect 20772 35040 20821 35068
rect 20772 35028 20778 35040
rect 20809 35037 20821 35040
rect 20855 35037 20867 35071
rect 21450 35068 21456 35080
rect 21411 35040 21456 35068
rect 20809 35031 20867 35037
rect 21450 35028 21456 35040
rect 21508 35028 21514 35080
rect 22121 35071 22179 35077
rect 22121 35037 22133 35071
rect 22167 35068 22179 35071
rect 22370 35068 22376 35080
rect 22167 35040 22376 35068
rect 22167 35037 22179 35040
rect 22121 35031 22179 35037
rect 22370 35028 22376 35040
rect 22428 35028 22434 35080
rect 22741 35071 22799 35077
rect 22741 35037 22753 35071
rect 22787 35068 22799 35071
rect 23474 35068 23480 35080
rect 22787 35040 23480 35068
rect 22787 35037 22799 35040
rect 22741 35031 22799 35037
rect 14826 35000 14832 35012
rect 3252 34972 6040 35000
rect 6380 34972 6762 35000
rect 12466 34972 14832 35000
rect 2682 34932 2688 34944
rect 1596 34904 2688 34932
rect 2682 34892 2688 34904
rect 2740 34932 2746 34944
rect 3252 34932 3280 34972
rect 2740 34904 3280 34932
rect 2740 34892 2746 34904
rect 4614 34892 4620 34944
rect 4672 34932 4678 34944
rect 6380 34932 6408 34972
rect 14826 34960 14832 34972
rect 14884 34960 14890 35012
rect 16146 34972 17080 35000
rect 7742 34932 7748 34944
rect 4672 34904 6408 34932
rect 7655 34904 7748 34932
rect 4672 34892 4678 34904
rect 7742 34892 7748 34904
rect 7800 34932 7806 34944
rect 12618 34932 12624 34944
rect 7800 34904 12624 34932
rect 7800 34892 7806 34904
rect 12618 34892 12624 34904
rect 12676 34892 12682 34944
rect 12710 34892 12716 34944
rect 12768 34932 12774 34944
rect 16942 34932 16948 34944
rect 12768 34904 16948 34932
rect 12768 34892 12774 34904
rect 16942 34892 16948 34904
rect 17000 34892 17006 34944
rect 17052 34932 17080 34972
rect 18432 34972 21680 35000
rect 18432 34932 18460 34972
rect 18598 34932 18604 34944
rect 17052 34904 18460 34932
rect 18559 34904 18604 34932
rect 18598 34892 18604 34904
rect 18656 34892 18662 34944
rect 19521 34935 19579 34941
rect 19521 34901 19533 34935
rect 19567 34932 19579 34935
rect 20162 34932 20168 34944
rect 19567 34904 20168 34932
rect 19567 34901 19579 34904
rect 19521 34895 19579 34901
rect 20162 34892 20168 34904
rect 20220 34892 20226 34944
rect 20257 34935 20315 34941
rect 20257 34901 20269 34935
rect 20303 34932 20315 34935
rect 20438 34932 20444 34944
rect 20303 34904 20444 34932
rect 20303 34901 20315 34904
rect 20257 34895 20315 34901
rect 20438 34892 20444 34904
rect 20496 34892 20502 34944
rect 20714 34892 20720 34944
rect 20772 34932 20778 34944
rect 20901 34935 20959 34941
rect 20901 34932 20913 34935
rect 20772 34904 20913 34932
rect 20772 34892 20778 34904
rect 20901 34901 20913 34904
rect 20947 34901 20959 34935
rect 20901 34895 20959 34901
rect 20990 34892 20996 34944
rect 21048 34932 21054 34944
rect 21545 34935 21603 34941
rect 21545 34932 21557 34935
rect 21048 34904 21557 34932
rect 21048 34892 21054 34904
rect 21545 34901 21557 34904
rect 21591 34901 21603 34935
rect 21652 34932 21680 34972
rect 21818 34960 21824 35012
rect 21876 35000 21882 35012
rect 22756 35000 22784 35031
rect 23474 35028 23480 35040
rect 23532 35028 23538 35080
rect 23658 35068 23664 35080
rect 23619 35040 23664 35068
rect 23658 35028 23664 35040
rect 23716 35028 23722 35080
rect 24581 35071 24639 35077
rect 24581 35037 24593 35071
rect 24627 35068 24639 35071
rect 25225 35071 25283 35077
rect 25225 35068 25237 35071
rect 24627 35040 25237 35068
rect 24627 35037 24639 35040
rect 24581 35031 24639 35037
rect 25225 35037 25237 35040
rect 25271 35068 25283 35071
rect 25590 35068 25596 35080
rect 25271 35040 25596 35068
rect 25271 35037 25283 35040
rect 25225 35031 25283 35037
rect 21876 34972 22784 35000
rect 23492 35000 23520 35028
rect 24596 35000 24624 35031
rect 25590 35028 25596 35040
rect 25648 35028 25654 35080
rect 27540 35068 27568 35108
rect 27801 35105 27813 35108
rect 27847 35105 27859 35139
rect 28166 35136 28172 35148
rect 28127 35108 28172 35136
rect 27801 35099 27859 35105
rect 28166 35096 28172 35108
rect 28224 35096 28230 35148
rect 28368 35136 28396 35164
rect 31726 35136 31754 35176
rect 28368 35108 31248 35136
rect 31726 35108 35894 35136
rect 28902 35068 28908 35080
rect 27080 35040 27568 35068
rect 28863 35040 28908 35068
rect 23492 34972 24624 35000
rect 26329 35003 26387 35009
rect 21876 34960 21882 34972
rect 26329 34969 26341 35003
rect 26375 34969 26387 35003
rect 26329 34963 26387 34969
rect 22189 34935 22247 34941
rect 22189 34932 22201 34935
rect 21652 34904 22201 34932
rect 21545 34895 21603 34901
rect 22189 34901 22201 34904
rect 22235 34901 22247 34935
rect 22830 34932 22836 34944
rect 22791 34904 22836 34932
rect 22189 34895 22247 34901
rect 22830 34892 22836 34904
rect 22888 34892 22894 34944
rect 22922 34892 22928 34944
rect 22980 34932 22986 34944
rect 25317 34935 25375 34941
rect 25317 34932 25329 34935
rect 22980 34904 25329 34932
rect 22980 34892 22986 34904
rect 25317 34901 25329 34904
rect 25363 34901 25375 34935
rect 26344 34932 26372 34963
rect 26878 34960 26884 35012
rect 26936 35000 26942 35012
rect 27080 35000 27108 35040
rect 28902 35028 28908 35040
rect 28960 35028 28966 35080
rect 29914 35068 29920 35080
rect 29875 35040 29920 35068
rect 29914 35028 29920 35040
rect 29972 35028 29978 35080
rect 30006 35028 30012 35080
rect 30064 35068 30070 35080
rect 31220 35077 31248 35108
rect 30377 35071 30435 35077
rect 30377 35068 30389 35071
rect 30064 35040 30389 35068
rect 30064 35028 30070 35040
rect 30377 35037 30389 35040
rect 30423 35037 30435 35071
rect 30377 35031 30435 35037
rect 31205 35071 31263 35077
rect 31205 35037 31217 35071
rect 31251 35037 31263 35071
rect 35866 35068 35894 35108
rect 37829 35071 37887 35077
rect 37829 35068 37841 35071
rect 35866 35040 37841 35068
rect 31205 35031 31263 35037
rect 37829 35037 37841 35040
rect 37875 35037 37887 35071
rect 37829 35031 37887 35037
rect 26936 34972 27108 35000
rect 26936 34960 26942 34972
rect 27154 34960 27160 35012
rect 27212 35000 27218 35012
rect 27249 35003 27307 35009
rect 27249 35000 27261 35003
rect 27212 34972 27261 35000
rect 27212 34960 27218 34972
rect 27249 34969 27261 34972
rect 27295 35000 27307 35003
rect 27522 35000 27528 35012
rect 27295 34972 27528 35000
rect 27295 34969 27307 34972
rect 27249 34963 27307 34969
rect 27522 34960 27528 34972
rect 27580 34960 27586 35012
rect 27890 35000 27896 35012
rect 27851 34972 27896 35000
rect 27890 34960 27896 34972
rect 27948 34960 27954 35012
rect 27982 34960 27988 35012
rect 28040 35000 28046 35012
rect 31018 35000 31024 35012
rect 28040 34972 31024 35000
rect 28040 34960 28046 34972
rect 31018 34960 31024 34972
rect 31076 34960 31082 35012
rect 28534 34932 28540 34944
rect 26344 34904 28540 34932
rect 25317 34895 25375 34901
rect 28534 34892 28540 34904
rect 28592 34892 28598 34944
rect 28994 34932 29000 34944
rect 28955 34904 29000 34932
rect 28994 34892 29000 34904
rect 29052 34892 29058 34944
rect 29270 34892 29276 34944
rect 29328 34932 29334 34944
rect 29733 34935 29791 34941
rect 29733 34932 29745 34935
rect 29328 34904 29745 34932
rect 29328 34892 29334 34904
rect 29733 34901 29745 34904
rect 29779 34901 29791 34935
rect 38010 34932 38016 34944
rect 37971 34904 38016 34932
rect 29733 34895 29791 34901
rect 38010 34892 38016 34904
rect 38068 34892 38074 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 3326 34728 3332 34740
rect 1627 34700 3332 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 3326 34688 3332 34700
rect 3384 34688 3390 34740
rect 5350 34728 5356 34740
rect 3896 34700 5212 34728
rect 5263 34700 5356 34728
rect 3896 34660 3924 34700
rect 2240 34632 3924 34660
rect 1762 34592 1768 34604
rect 1723 34564 1768 34592
rect 1762 34552 1768 34564
rect 1820 34552 1826 34604
rect 2240 34601 2268 34632
rect 3970 34620 3976 34672
rect 4028 34660 4034 34672
rect 4028 34632 4370 34660
rect 4028 34620 4034 34632
rect 2225 34595 2283 34601
rect 2225 34561 2237 34595
rect 2271 34561 2283 34595
rect 2225 34555 2283 34561
rect 2317 34595 2375 34601
rect 2317 34561 2329 34595
rect 2363 34592 2375 34595
rect 2866 34592 2872 34604
rect 2363 34564 2872 34592
rect 2363 34561 2375 34564
rect 2317 34555 2375 34561
rect 2866 34552 2872 34564
rect 2924 34552 2930 34604
rect 5184 34592 5212 34700
rect 5350 34688 5356 34700
rect 5408 34688 5414 34740
rect 6546 34688 6552 34740
rect 6604 34728 6610 34740
rect 6641 34731 6699 34737
rect 6641 34728 6653 34731
rect 6604 34700 6653 34728
rect 6604 34688 6610 34700
rect 6641 34697 6653 34700
rect 6687 34697 6699 34731
rect 6641 34691 6699 34697
rect 10502 34688 10508 34740
rect 10560 34728 10566 34740
rect 11701 34731 11759 34737
rect 11701 34728 11713 34731
rect 10560 34700 11713 34728
rect 10560 34688 10566 34700
rect 11701 34697 11713 34700
rect 11747 34697 11759 34731
rect 15562 34728 15568 34740
rect 11701 34691 11759 34697
rect 11808 34700 15424 34728
rect 15523 34700 15568 34728
rect 5368 34660 5396 34688
rect 11808 34660 11836 34700
rect 13262 34660 13268 34672
rect 5368 34632 11836 34660
rect 11900 34632 13268 34660
rect 5718 34592 5724 34604
rect 5184 34564 5724 34592
rect 5718 34552 5724 34564
rect 5776 34592 5782 34604
rect 6270 34592 6276 34604
rect 5776 34564 6276 34592
rect 5776 34552 5782 34564
rect 6270 34552 6276 34564
rect 6328 34552 6334 34604
rect 6549 34595 6607 34601
rect 6549 34561 6561 34595
rect 6595 34592 6607 34595
rect 7742 34592 7748 34604
rect 6595 34564 7748 34592
rect 6595 34561 6607 34564
rect 6549 34555 6607 34561
rect 2682 34484 2688 34536
rect 2740 34524 2746 34536
rect 3605 34527 3663 34533
rect 3605 34524 3617 34527
rect 2740 34496 3617 34524
rect 2740 34484 2746 34496
rect 3605 34493 3617 34496
rect 3651 34493 3663 34527
rect 3605 34487 3663 34493
rect 3881 34527 3939 34533
rect 3881 34493 3893 34527
rect 3927 34524 3939 34527
rect 6564 34524 6592 34555
rect 7742 34552 7748 34564
rect 7800 34552 7806 34604
rect 8113 34595 8171 34601
rect 8113 34561 8125 34595
rect 8159 34561 8171 34595
rect 8113 34555 8171 34561
rect 8128 34524 8156 34555
rect 9582 34552 9588 34604
rect 9640 34592 9646 34604
rect 11900 34601 11928 34632
rect 13262 34620 13268 34632
rect 13320 34620 13326 34672
rect 14366 34620 14372 34672
rect 14424 34660 14430 34672
rect 15396 34660 15424 34700
rect 15562 34688 15568 34700
rect 15620 34688 15626 34740
rect 16666 34688 16672 34740
rect 16724 34728 16730 34740
rect 17862 34728 17868 34740
rect 16724 34700 17868 34728
rect 16724 34688 16730 34700
rect 17862 34688 17868 34700
rect 17920 34688 17926 34740
rect 17954 34688 17960 34740
rect 18012 34728 18018 34740
rect 19978 34728 19984 34740
rect 18012 34700 19984 34728
rect 18012 34688 18018 34700
rect 19978 34688 19984 34700
rect 20036 34688 20042 34740
rect 22094 34728 22100 34740
rect 20180 34700 22100 34728
rect 17402 34660 17408 34672
rect 14424 34632 14582 34660
rect 15396 34632 17408 34660
rect 14424 34620 14430 34632
rect 17402 34620 17408 34632
rect 17460 34620 17466 34672
rect 20180 34660 20208 34700
rect 22094 34688 22100 34700
rect 22152 34688 22158 34740
rect 23934 34688 23940 34740
rect 23992 34728 23998 34740
rect 25038 34728 25044 34740
rect 23992 34700 25044 34728
rect 23992 34688 23998 34700
rect 25038 34688 25044 34700
rect 25096 34688 25102 34740
rect 28534 34728 28540 34740
rect 26344 34700 28028 34728
rect 28495 34700 28540 34728
rect 18354 34632 20208 34660
rect 20530 34620 20536 34672
rect 20588 34660 20594 34672
rect 20901 34663 20959 34669
rect 20901 34660 20913 34663
rect 20588 34632 20913 34660
rect 20588 34620 20594 34632
rect 20901 34629 20913 34632
rect 20947 34629 20959 34663
rect 22462 34660 22468 34672
rect 22423 34632 22468 34660
rect 20901 34623 20959 34629
rect 22462 34620 22468 34632
rect 22520 34620 22526 34672
rect 25685 34663 25743 34669
rect 25685 34660 25697 34663
rect 22940 34632 25697 34660
rect 11885 34595 11943 34601
rect 11885 34592 11897 34595
rect 9640 34564 11897 34592
rect 9640 34552 9646 34564
rect 11885 34561 11897 34564
rect 11931 34561 11943 34595
rect 12434 34592 12440 34604
rect 11885 34555 11943 34561
rect 12406 34552 12440 34592
rect 12492 34552 12498 34604
rect 12618 34592 12624 34604
rect 12579 34564 12624 34592
rect 12618 34552 12624 34564
rect 12676 34552 12682 34604
rect 12710 34552 12716 34604
rect 12768 34592 12774 34604
rect 22370 34592 22376 34604
rect 12768 34564 12813 34592
rect 22331 34564 22376 34592
rect 12768 34552 12774 34564
rect 22370 34552 22376 34564
rect 22428 34552 22434 34604
rect 3927 34496 6592 34524
rect 6656 34496 8156 34524
rect 8205 34527 8263 34533
rect 3927 34493 3939 34496
rect 3881 34487 3939 34493
rect 6270 34416 6276 34468
rect 6328 34456 6334 34468
rect 6656 34456 6684 34496
rect 8205 34493 8217 34527
rect 8251 34524 8263 34527
rect 12406 34524 12434 34552
rect 8251 34496 12434 34524
rect 13817 34527 13875 34533
rect 8251 34493 8263 34496
rect 8205 34487 8263 34493
rect 13817 34493 13829 34527
rect 13863 34493 13875 34527
rect 13817 34487 13875 34493
rect 14093 34527 14151 34533
rect 14093 34493 14105 34527
rect 14139 34524 14151 34527
rect 16850 34524 16856 34536
rect 14139 34496 15148 34524
rect 16811 34496 16856 34524
rect 14139 34493 14151 34496
rect 14093 34487 14151 34493
rect 6328 34428 6684 34456
rect 6328 34416 6334 34428
rect 13170 34348 13176 34400
rect 13228 34388 13234 34400
rect 13832 34388 13860 34487
rect 15120 34456 15148 34496
rect 16850 34484 16856 34496
rect 16908 34484 16914 34536
rect 17218 34484 17224 34536
rect 17276 34524 17282 34536
rect 18601 34527 18659 34533
rect 18601 34524 18613 34527
rect 17276 34496 18613 34524
rect 17276 34484 17282 34496
rect 18601 34493 18613 34496
rect 18647 34524 18659 34527
rect 18647 34496 19334 34524
rect 18647 34493 18659 34496
rect 18601 34487 18659 34493
rect 16298 34456 16304 34468
rect 15120 34428 16304 34456
rect 16298 34416 16304 34428
rect 16356 34416 16362 34468
rect 16482 34416 16488 34468
rect 16540 34456 16546 34468
rect 16540 34428 16988 34456
rect 16540 34416 16546 34428
rect 16960 34400 16988 34428
rect 18138 34416 18144 34468
rect 18196 34456 18202 34468
rect 19306 34456 19334 34496
rect 20806 34484 20812 34536
rect 20864 34524 20870 34536
rect 21174 34524 21180 34536
rect 20864 34496 20909 34524
rect 21135 34496 21180 34524
rect 20864 34484 20870 34496
rect 21174 34484 21180 34496
rect 21232 34484 21238 34536
rect 21542 34484 21548 34536
rect 21600 34524 21606 34536
rect 22940 34524 22968 34632
rect 25685 34629 25697 34632
rect 25731 34629 25743 34663
rect 25685 34623 25743 34629
rect 23014 34552 23020 34604
rect 23072 34592 23078 34604
rect 23382 34592 23388 34604
rect 23072 34564 23388 34592
rect 23072 34552 23078 34564
rect 23382 34552 23388 34564
rect 23440 34552 23446 34604
rect 23661 34595 23719 34601
rect 23661 34592 23673 34595
rect 23492 34564 23673 34592
rect 23492 34536 23520 34564
rect 23661 34561 23673 34564
rect 23707 34561 23719 34595
rect 23661 34555 23719 34561
rect 23842 34552 23848 34604
rect 23900 34592 23906 34604
rect 24305 34595 24363 34601
rect 24305 34592 24317 34595
rect 23900 34564 24317 34592
rect 23900 34552 23906 34564
rect 24305 34561 24317 34564
rect 24351 34561 24363 34595
rect 24305 34555 24363 34561
rect 24949 34595 25007 34601
rect 24949 34561 24961 34595
rect 24995 34561 25007 34595
rect 25590 34592 25596 34604
rect 25551 34564 25596 34592
rect 24949 34555 25007 34561
rect 23106 34524 23112 34536
rect 21600 34496 22968 34524
rect 23067 34496 23112 34524
rect 21600 34484 21606 34496
rect 23106 34484 23112 34496
rect 23164 34484 23170 34536
rect 23474 34484 23480 34536
rect 23532 34484 23538 34536
rect 23750 34524 23756 34536
rect 23711 34496 23756 34524
rect 23750 34484 23756 34496
rect 23808 34484 23814 34536
rect 24964 34524 24992 34555
rect 25590 34552 25596 34564
rect 25648 34552 25654 34604
rect 26237 34595 26295 34601
rect 26237 34561 26249 34595
rect 26283 34590 26295 34595
rect 26344 34590 26372 34700
rect 27893 34663 27951 34669
rect 27893 34660 27905 34663
rect 27264 34632 27905 34660
rect 26283 34562 26372 34590
rect 26283 34561 26295 34562
rect 26237 34555 26295 34561
rect 26418 34552 26424 34604
rect 26476 34592 26482 34604
rect 27157 34595 27215 34601
rect 27157 34592 27169 34595
rect 26476 34564 27169 34592
rect 26476 34552 26482 34564
rect 27157 34561 27169 34564
rect 27203 34561 27215 34595
rect 27157 34555 27215 34561
rect 23860 34496 24992 34524
rect 25041 34527 25099 34533
rect 22278 34456 22284 34468
rect 18196 34428 18644 34456
rect 19306 34428 22284 34456
rect 18196 34416 18202 34428
rect 14642 34388 14648 34400
rect 13228 34360 14648 34388
rect 13228 34348 13234 34360
rect 14642 34348 14648 34360
rect 14700 34348 14706 34400
rect 15838 34348 15844 34400
rect 15896 34388 15902 34400
rect 16666 34388 16672 34400
rect 15896 34360 16672 34388
rect 15896 34348 15902 34360
rect 16666 34348 16672 34360
rect 16724 34348 16730 34400
rect 16942 34348 16948 34400
rect 17000 34348 17006 34400
rect 17116 34391 17174 34397
rect 17116 34357 17128 34391
rect 17162 34388 17174 34391
rect 18506 34388 18512 34400
rect 17162 34360 18512 34388
rect 17162 34357 17174 34360
rect 17116 34351 17174 34357
rect 18506 34348 18512 34360
rect 18564 34348 18570 34400
rect 18616 34388 18644 34428
rect 22278 34416 22284 34428
rect 22336 34416 22342 34468
rect 23198 34456 23204 34468
rect 22388 34428 23204 34456
rect 22388 34388 22416 34428
rect 23198 34416 23204 34428
rect 23256 34416 23262 34468
rect 23566 34416 23572 34468
rect 23624 34456 23630 34468
rect 23860 34456 23888 34496
rect 25041 34493 25053 34527
rect 25087 34524 25099 34527
rect 25222 34524 25228 34536
rect 25087 34496 25228 34524
rect 25087 34493 25099 34496
rect 25041 34487 25099 34493
rect 25222 34484 25228 34496
rect 25280 34484 25286 34536
rect 25314 34484 25320 34536
rect 25372 34524 25378 34536
rect 26329 34527 26387 34533
rect 26329 34524 26341 34527
rect 25372 34496 26341 34524
rect 25372 34484 25378 34496
rect 26329 34493 26341 34496
rect 26375 34493 26387 34527
rect 26329 34487 26387 34493
rect 26878 34484 26884 34536
rect 26936 34524 26942 34536
rect 27264 34524 27292 34632
rect 27893 34629 27905 34632
rect 27939 34629 27951 34663
rect 27893 34623 27951 34629
rect 27798 34592 27804 34604
rect 27759 34564 27804 34592
rect 27798 34552 27804 34564
rect 27856 34552 27862 34604
rect 28000 34592 28028 34700
rect 28534 34688 28540 34700
rect 28592 34688 28598 34740
rect 29822 34728 29828 34740
rect 29783 34700 29828 34728
rect 29822 34688 29828 34700
rect 29880 34688 29886 34740
rect 30374 34688 30380 34740
rect 30432 34728 30438 34740
rect 30469 34731 30527 34737
rect 30469 34728 30481 34731
rect 30432 34700 30481 34728
rect 30432 34688 30438 34700
rect 30469 34697 30481 34700
rect 30515 34697 30527 34731
rect 30469 34691 30527 34697
rect 28074 34620 28080 34672
rect 28132 34660 28138 34672
rect 28132 34632 29132 34660
rect 28132 34620 28138 34632
rect 28442 34592 28448 34604
rect 28000 34564 28448 34592
rect 28442 34552 28448 34564
rect 28500 34552 28506 34604
rect 29104 34601 29132 34632
rect 29089 34595 29147 34601
rect 29089 34561 29101 34595
rect 29135 34561 29147 34595
rect 29733 34595 29791 34601
rect 29733 34592 29745 34595
rect 29089 34555 29147 34561
rect 29288 34564 29745 34592
rect 26936 34496 27292 34524
rect 26936 34484 26942 34496
rect 27430 34484 27436 34536
rect 27488 34524 27494 34536
rect 29181 34527 29239 34533
rect 29181 34524 29193 34527
rect 27488 34496 29193 34524
rect 27488 34484 27494 34496
rect 29181 34493 29193 34496
rect 29227 34493 29239 34527
rect 29181 34487 29239 34493
rect 29288 34456 29316 34564
rect 29733 34561 29745 34564
rect 29779 34561 29791 34595
rect 29733 34555 29791 34561
rect 30377 34595 30435 34601
rect 30377 34561 30389 34595
rect 30423 34592 30435 34595
rect 36722 34592 36728 34604
rect 30423 34564 36728 34592
rect 30423 34561 30435 34564
rect 30377 34555 30435 34561
rect 36722 34552 36728 34564
rect 36780 34552 36786 34604
rect 37826 34552 37832 34604
rect 37884 34592 37890 34604
rect 38013 34595 38071 34601
rect 38013 34592 38025 34595
rect 37884 34564 38025 34592
rect 37884 34552 37890 34564
rect 38013 34561 38025 34564
rect 38059 34561 38071 34595
rect 38013 34555 38071 34561
rect 30006 34524 30012 34536
rect 23624 34428 23888 34456
rect 23952 34428 29316 34456
rect 29380 34496 30012 34524
rect 23624 34416 23630 34428
rect 18616 34360 22416 34388
rect 22554 34348 22560 34400
rect 22612 34388 22618 34400
rect 23952 34388 23980 34428
rect 24394 34388 24400 34400
rect 22612 34360 23980 34388
rect 24355 34360 24400 34388
rect 22612 34348 22618 34360
rect 24394 34348 24400 34360
rect 24452 34348 24458 34400
rect 26694 34348 26700 34400
rect 26752 34388 26758 34400
rect 27249 34391 27307 34397
rect 27249 34388 27261 34391
rect 26752 34360 27261 34388
rect 26752 34348 26758 34360
rect 27249 34357 27261 34360
rect 27295 34357 27307 34391
rect 27249 34351 27307 34357
rect 27522 34348 27528 34400
rect 27580 34388 27586 34400
rect 29380 34388 29408 34496
rect 30006 34484 30012 34496
rect 30064 34484 30070 34536
rect 38194 34388 38200 34400
rect 27580 34360 29408 34388
rect 38155 34360 38200 34388
rect 27580 34348 27586 34360
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 4065 34187 4123 34193
rect 4065 34153 4077 34187
rect 4111 34184 4123 34187
rect 4614 34184 4620 34196
rect 4111 34156 4620 34184
rect 4111 34153 4123 34156
rect 4065 34147 4123 34153
rect 4614 34144 4620 34156
rect 4672 34144 4678 34196
rect 8202 34144 8208 34196
rect 8260 34184 8266 34196
rect 8481 34187 8539 34193
rect 8481 34184 8493 34187
rect 8260 34156 8493 34184
rect 8260 34144 8266 34156
rect 8481 34153 8493 34156
rect 8527 34153 8539 34187
rect 8481 34147 8539 34153
rect 13722 34144 13728 34196
rect 13780 34184 13786 34196
rect 22189 34187 22247 34193
rect 22189 34184 22201 34187
rect 13780 34156 22201 34184
rect 13780 34144 13786 34156
rect 22189 34153 22201 34156
rect 22235 34153 22247 34187
rect 27246 34184 27252 34196
rect 22189 34147 22247 34153
rect 23400 34156 27252 34184
rect 15838 34116 15844 34128
rect 13740 34088 15844 34116
rect 6733 34051 6791 34057
rect 6733 34017 6745 34051
rect 6779 34048 6791 34051
rect 8938 34048 8944 34060
rect 6779 34020 8944 34048
rect 6779 34017 6791 34020
rect 6733 34011 6791 34017
rect 8938 34008 8944 34020
rect 8996 34008 9002 34060
rect 11054 34048 11060 34060
rect 11015 34020 11060 34048
rect 11054 34008 11060 34020
rect 11112 34008 11118 34060
rect 11977 34051 12035 34057
rect 11977 34017 11989 34051
rect 12023 34048 12035 34051
rect 13262 34048 13268 34060
rect 12023 34020 13268 34048
rect 12023 34017 12035 34020
rect 11977 34011 12035 34017
rect 13262 34008 13268 34020
rect 13320 34008 13326 34060
rect 13740 34057 13768 34088
rect 15838 34076 15844 34088
rect 15896 34076 15902 34128
rect 18506 34116 18512 34128
rect 17328 34088 18512 34116
rect 13725 34051 13783 34057
rect 13725 34017 13737 34051
rect 13771 34017 13783 34051
rect 13725 34011 13783 34017
rect 14642 34008 14648 34060
rect 14700 34048 14706 34060
rect 15013 34051 15071 34057
rect 15013 34048 15025 34051
rect 14700 34020 15025 34048
rect 14700 34008 14706 34020
rect 15013 34017 15025 34020
rect 15059 34017 15071 34051
rect 15013 34011 15071 34017
rect 15933 34051 15991 34057
rect 15933 34017 15945 34051
rect 15979 34048 15991 34051
rect 16850 34048 16856 34060
rect 15979 34020 16856 34048
rect 15979 34017 15991 34020
rect 15933 34011 15991 34017
rect 16850 34008 16856 34020
rect 16908 34008 16914 34060
rect 16942 34008 16948 34060
rect 17000 34048 17006 34060
rect 17328 34048 17356 34088
rect 18506 34076 18512 34088
rect 18564 34076 18570 34128
rect 18598 34076 18604 34128
rect 18656 34116 18662 34128
rect 23400 34116 23428 34156
rect 27246 34144 27252 34156
rect 27304 34144 27310 34196
rect 28997 34187 29055 34193
rect 27356 34156 28396 34184
rect 23566 34116 23572 34128
rect 18656 34088 23428 34116
rect 23527 34088 23572 34116
rect 18656 34076 18662 34088
rect 23566 34076 23572 34088
rect 23624 34116 23630 34128
rect 23624 34088 24716 34116
rect 23624 34076 23630 34088
rect 17000 34020 17356 34048
rect 17000 34008 17006 34020
rect 17402 34008 17408 34060
rect 17460 34048 17466 34060
rect 18414 34048 18420 34060
rect 17460 34020 18420 34048
rect 17460 34008 17466 34020
rect 18414 34008 18420 34020
rect 18472 34008 18478 34060
rect 23201 34051 23259 34057
rect 23201 34017 23213 34051
rect 23247 34048 23259 34051
rect 23934 34048 23940 34060
rect 23247 34020 23940 34048
rect 23247 34017 23259 34020
rect 23201 34011 23259 34017
rect 23934 34008 23940 34020
rect 23992 34008 23998 34060
rect 24688 34057 24716 34088
rect 25498 34076 25504 34128
rect 25556 34116 25562 34128
rect 27356 34116 27384 34156
rect 28166 34116 28172 34128
rect 25556 34088 27384 34116
rect 27540 34088 28172 34116
rect 25556 34076 25562 34088
rect 24673 34051 24731 34057
rect 24673 34017 24685 34051
rect 24719 34017 24731 34051
rect 24946 34048 24952 34060
rect 24907 34020 24952 34048
rect 24673 34011 24731 34017
rect 24946 34008 24952 34020
rect 25004 34008 25010 34060
rect 25406 34008 25412 34060
rect 25464 34048 25470 34060
rect 27430 34048 27436 34060
rect 25464 34020 27436 34048
rect 25464 34008 25470 34020
rect 27430 34008 27436 34020
rect 27488 34008 27494 34060
rect 3418 33940 3424 33992
rect 3476 33980 3482 33992
rect 3973 33983 4031 33989
rect 3973 33980 3985 33983
rect 3476 33952 3985 33980
rect 3476 33940 3482 33952
rect 3973 33949 3985 33952
rect 4019 33949 4031 33983
rect 3973 33943 4031 33949
rect 8110 33940 8116 33992
rect 8168 33940 8174 33992
rect 14277 33983 14335 33989
rect 14277 33949 14289 33983
rect 14323 33980 14335 33983
rect 15378 33980 15384 33992
rect 14323 33952 15384 33980
rect 14323 33949 14335 33952
rect 14277 33943 14335 33949
rect 15378 33940 15384 33952
rect 15436 33940 15442 33992
rect 19150 33980 19156 33992
rect 17342 33952 19156 33980
rect 19150 33940 19156 33952
rect 19208 33940 19214 33992
rect 20254 33940 20260 33992
rect 20312 33980 20318 33992
rect 22097 33983 22155 33989
rect 22097 33980 22109 33983
rect 20312 33952 22109 33980
rect 20312 33940 20318 33952
rect 22097 33949 22109 33952
rect 22143 33980 22155 33983
rect 22370 33980 22376 33992
rect 22143 33952 22376 33980
rect 22143 33949 22155 33952
rect 22097 33943 22155 33949
rect 22370 33940 22376 33952
rect 22428 33940 22434 33992
rect 23385 33983 23443 33989
rect 23385 33949 23397 33983
rect 23431 33980 23443 33983
rect 24486 33980 24492 33992
rect 23431 33952 24492 33980
rect 23431 33949 23443 33952
rect 23385 33943 23443 33949
rect 24486 33940 24492 33952
rect 24544 33940 24550 33992
rect 25590 33940 25596 33992
rect 25648 33980 25654 33992
rect 25777 33983 25835 33989
rect 25777 33980 25789 33983
rect 25648 33952 25789 33980
rect 25648 33940 25654 33952
rect 25777 33949 25789 33952
rect 25823 33949 25835 33983
rect 25777 33943 25835 33949
rect 27249 33983 27307 33989
rect 27249 33949 27261 33983
rect 27295 33980 27307 33983
rect 27540 33980 27568 34088
rect 28166 34076 28172 34088
rect 28224 34076 28230 34128
rect 28368 34125 28396 34156
rect 28997 34153 29009 34187
rect 29043 34184 29055 34187
rect 29086 34184 29092 34196
rect 29043 34156 29092 34184
rect 29043 34153 29055 34156
rect 28997 34147 29055 34153
rect 29086 34144 29092 34156
rect 29144 34144 29150 34196
rect 37826 34184 37832 34196
rect 37787 34156 37832 34184
rect 37826 34144 37832 34156
rect 37884 34144 37890 34196
rect 28353 34119 28411 34125
rect 28353 34085 28365 34119
rect 28399 34116 28411 34119
rect 29178 34116 29184 34128
rect 28399 34088 29184 34116
rect 28399 34085 28411 34088
rect 28353 34079 28411 34085
rect 29178 34076 29184 34088
rect 29236 34076 29242 34128
rect 27801 34051 27859 34057
rect 27801 34017 27813 34051
rect 27847 34048 27859 34051
rect 28994 34048 29000 34060
rect 27847 34020 29000 34048
rect 27847 34017 27859 34020
rect 27801 34011 27859 34017
rect 28994 34008 29000 34020
rect 29052 34008 29058 34060
rect 27295 33952 27568 33980
rect 27295 33949 27307 33952
rect 27249 33943 27307 33949
rect 28534 33940 28540 33992
rect 28592 33980 28598 33992
rect 28905 33983 28963 33989
rect 28905 33980 28917 33983
rect 28592 33952 28917 33980
rect 28592 33940 28598 33952
rect 28905 33949 28917 33952
rect 28951 33949 28963 33983
rect 28905 33943 28963 33949
rect 30377 33983 30435 33989
rect 30377 33949 30389 33983
rect 30423 33980 30435 33983
rect 33042 33980 33048 33992
rect 30423 33952 33048 33980
rect 30423 33949 30435 33952
rect 30377 33943 30435 33949
rect 33042 33940 33048 33952
rect 33100 33940 33106 33992
rect 38010 33980 38016 33992
rect 37971 33952 38016 33980
rect 38010 33940 38016 33952
rect 38068 33940 38074 33992
rect 7009 33915 7067 33921
rect 7009 33881 7021 33915
rect 7055 33881 7067 33915
rect 7009 33875 7067 33881
rect 7024 33844 7052 33875
rect 10318 33872 10324 33924
rect 10376 33912 10382 33924
rect 10505 33915 10563 33921
rect 10505 33912 10517 33915
rect 10376 33884 10517 33912
rect 10376 33872 10382 33884
rect 10505 33881 10517 33884
rect 10551 33881 10563 33915
rect 10505 33875 10563 33881
rect 10594 33872 10600 33924
rect 10652 33912 10658 33924
rect 12253 33915 12311 33921
rect 10652 33884 10697 33912
rect 10652 33872 10658 33884
rect 12253 33881 12265 33915
rect 12299 33912 12311 33915
rect 12526 33912 12532 33924
rect 12299 33884 12532 33912
rect 12299 33881 12311 33884
rect 12253 33875 12311 33881
rect 12526 33872 12532 33884
rect 12584 33872 12590 33924
rect 13478 33884 16160 33912
rect 11422 33844 11428 33856
rect 7024 33816 11428 33844
rect 11422 33804 11428 33816
rect 11480 33804 11486 33856
rect 11698 33804 11704 33856
rect 11756 33844 11762 33856
rect 16022 33844 16028 33856
rect 11756 33816 16028 33844
rect 11756 33804 11762 33816
rect 16022 33804 16028 33816
rect 16080 33804 16086 33856
rect 16132 33844 16160 33884
rect 16206 33872 16212 33924
rect 16264 33912 16270 33924
rect 22830 33912 22836 33924
rect 16264 33884 16309 33912
rect 17512 33884 22836 33912
rect 16264 33872 16270 33884
rect 17512 33844 17540 33884
rect 22830 33872 22836 33884
rect 22888 33872 22894 33924
rect 24765 33915 24823 33921
rect 24765 33881 24777 33915
rect 24811 33881 24823 33915
rect 24765 33875 24823 33881
rect 26605 33915 26663 33921
rect 26605 33881 26617 33915
rect 26651 33881 26663 33915
rect 26605 33875 26663 33881
rect 17678 33844 17684 33856
rect 16132 33816 17540 33844
rect 17639 33816 17684 33844
rect 17678 33804 17684 33816
rect 17736 33804 17742 33856
rect 17862 33804 17868 33856
rect 17920 33844 17926 33856
rect 21174 33844 21180 33856
rect 17920 33816 21180 33844
rect 17920 33804 17926 33816
rect 21174 33804 21180 33816
rect 21232 33804 21238 33856
rect 24773 33844 24801 33875
rect 25406 33844 25412 33856
rect 24773 33816 25412 33844
rect 25406 33804 25412 33816
rect 25464 33804 25470 33856
rect 25866 33844 25872 33856
rect 25827 33816 25872 33844
rect 25866 33804 25872 33816
rect 25924 33804 25930 33856
rect 26620 33844 26648 33875
rect 26694 33872 26700 33924
rect 26752 33912 26758 33924
rect 26752 33884 26797 33912
rect 26752 33872 26758 33884
rect 27798 33872 27804 33924
rect 27856 33912 27862 33924
rect 27893 33915 27951 33921
rect 27893 33912 27905 33915
rect 27856 33884 27905 33912
rect 27856 33872 27862 33884
rect 27893 33881 27905 33884
rect 27939 33881 27951 33915
rect 27893 33875 27951 33881
rect 27982 33844 27988 33856
rect 26620 33816 27988 33844
rect 27982 33804 27988 33816
rect 28040 33804 28046 33856
rect 29730 33844 29736 33856
rect 29691 33816 29736 33844
rect 29730 33804 29736 33816
rect 29788 33804 29794 33856
rect 29822 33804 29828 33856
rect 29880 33844 29886 33856
rect 30469 33847 30527 33853
rect 30469 33844 30481 33847
rect 29880 33816 30481 33844
rect 29880 33804 29886 33816
rect 30469 33813 30481 33816
rect 30515 33813 30527 33847
rect 30469 33807 30527 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 4798 33640 4804 33652
rect 1596 33612 4804 33640
rect 1596 33513 1624 33612
rect 4798 33600 4804 33612
rect 4856 33600 4862 33652
rect 10594 33600 10600 33652
rect 10652 33640 10658 33652
rect 11793 33643 11851 33649
rect 11793 33640 11805 33643
rect 10652 33612 11805 33640
rect 10652 33600 10658 33612
rect 11793 33609 11805 33612
rect 11839 33609 11851 33643
rect 11793 33603 11851 33609
rect 14921 33643 14979 33649
rect 14921 33609 14933 33643
rect 14967 33640 14979 33643
rect 15838 33640 15844 33652
rect 14967 33612 15844 33640
rect 14967 33609 14979 33612
rect 14921 33603 14979 33609
rect 15838 33600 15844 33612
rect 15896 33640 15902 33652
rect 16206 33640 16212 33652
rect 15896 33612 16212 33640
rect 15896 33600 15902 33612
rect 16206 33600 16212 33612
rect 16264 33600 16270 33652
rect 17402 33600 17408 33652
rect 17460 33600 17466 33652
rect 17494 33600 17500 33652
rect 17552 33640 17558 33652
rect 20898 33640 20904 33652
rect 17552 33612 20904 33640
rect 17552 33600 17558 33612
rect 20898 33600 20904 33612
rect 20956 33600 20962 33652
rect 21082 33640 21088 33652
rect 21043 33612 21088 33640
rect 21082 33600 21088 33612
rect 21140 33600 21146 33652
rect 21174 33600 21180 33652
rect 21232 33640 21238 33652
rect 23477 33643 23535 33649
rect 23477 33640 23489 33643
rect 21232 33612 23489 33640
rect 21232 33600 21238 33612
rect 23477 33609 23489 33612
rect 23523 33609 23535 33643
rect 23477 33603 23535 33609
rect 24486 33600 24492 33652
rect 24544 33640 24550 33652
rect 26421 33643 26479 33649
rect 26421 33640 26433 33643
rect 24544 33612 26433 33640
rect 24544 33600 24550 33612
rect 26421 33609 26433 33612
rect 26467 33609 26479 33643
rect 29730 33640 29736 33652
rect 26421 33603 26479 33609
rect 28920 33612 29736 33640
rect 2682 33572 2688 33584
rect 2516 33544 2688 33572
rect 2516 33513 2544 33544
rect 2682 33532 2688 33544
rect 2740 33532 2746 33584
rect 2774 33532 2780 33584
rect 2832 33572 2838 33584
rect 7745 33575 7803 33581
rect 2832 33544 3266 33572
rect 2832 33532 2838 33544
rect 7745 33541 7757 33575
rect 7791 33572 7803 33575
rect 7834 33572 7840 33584
rect 7791 33544 7840 33572
rect 7791 33541 7803 33544
rect 7745 33535 7803 33541
rect 7834 33532 7840 33544
rect 7892 33532 7898 33584
rect 13722 33572 13728 33584
rect 8970 33544 13728 33572
rect 13722 33532 13728 33544
rect 13780 33532 13786 33584
rect 17126 33572 17132 33584
rect 14674 33544 17132 33572
rect 17126 33532 17132 33544
rect 17184 33532 17190 33584
rect 17221 33575 17279 33581
rect 17221 33541 17233 33575
rect 17267 33572 17279 33575
rect 17420 33572 17448 33600
rect 17267 33544 17448 33572
rect 22572 33544 23152 33572
rect 17267 33541 17279 33544
rect 17221 33535 17279 33541
rect 1581 33507 1639 33513
rect 1581 33473 1593 33507
rect 1627 33473 1639 33507
rect 1581 33467 1639 33473
rect 2501 33507 2559 33513
rect 2501 33473 2513 33507
rect 2547 33473 2559 33507
rect 2501 33467 2559 33473
rect 4985 33507 5043 33513
rect 4985 33473 4997 33507
rect 5031 33504 5043 33507
rect 6178 33504 6184 33516
rect 5031 33476 6184 33504
rect 5031 33473 5043 33476
rect 4985 33467 5043 33473
rect 6178 33464 6184 33476
rect 6236 33464 6242 33516
rect 11698 33504 11704 33516
rect 9324 33476 11704 33504
rect 2777 33439 2835 33445
rect 2777 33405 2789 33439
rect 2823 33436 2835 33439
rect 3142 33436 3148 33448
rect 2823 33408 3148 33436
rect 2823 33405 2835 33408
rect 2777 33399 2835 33405
rect 3142 33396 3148 33408
rect 3200 33396 3206 33448
rect 5534 33396 5540 33448
rect 5592 33436 5598 33448
rect 5629 33439 5687 33445
rect 5629 33436 5641 33439
rect 5592 33408 5641 33436
rect 5592 33396 5598 33408
rect 5629 33405 5641 33408
rect 5675 33405 5687 33439
rect 7466 33436 7472 33448
rect 7427 33408 7472 33436
rect 5629 33399 5687 33405
rect 7466 33396 7472 33408
rect 7524 33396 7530 33448
rect 8202 33396 8208 33448
rect 8260 33436 8266 33448
rect 9324 33436 9352 33476
rect 11698 33464 11704 33476
rect 11756 33464 11762 33516
rect 13170 33504 13176 33516
rect 13131 33476 13176 33504
rect 13170 33464 13176 33476
rect 13228 33464 13234 33516
rect 20990 33504 20996 33516
rect 8260 33408 9352 33436
rect 8260 33396 8266 33408
rect 9398 33396 9404 33448
rect 9456 33436 9462 33448
rect 9493 33439 9551 33445
rect 9493 33436 9505 33439
rect 9456 33408 9505 33436
rect 9456 33396 9462 33408
rect 9493 33405 9505 33408
rect 9539 33405 9551 33439
rect 9493 33399 9551 33405
rect 13449 33439 13507 33445
rect 13449 33405 13461 33439
rect 13495 33436 13507 33439
rect 13998 33436 14004 33448
rect 13495 33408 14004 33436
rect 13495 33405 13507 33408
rect 13449 33399 13507 33405
rect 13998 33396 14004 33408
rect 14056 33396 14062 33448
rect 16850 33396 16856 33448
rect 16908 33436 16914 33448
rect 16945 33439 17003 33445
rect 16945 33436 16957 33439
rect 16908 33408 16957 33436
rect 16908 33396 16914 33408
rect 16945 33405 16957 33408
rect 16991 33405 17003 33439
rect 17862 33436 17868 33448
rect 16945 33399 17003 33405
rect 17052 33408 17868 33436
rect 1762 33368 1768 33380
rect 1723 33340 1768 33368
rect 1762 33328 1768 33340
rect 1820 33328 1826 33380
rect 15102 33328 15108 33380
rect 15160 33368 15166 33380
rect 17052 33368 17080 33408
rect 17862 33396 17868 33408
rect 17920 33396 17926 33448
rect 18340 33436 18368 33490
rect 20951 33476 20996 33504
rect 20990 33464 20996 33476
rect 21048 33464 21054 33516
rect 22005 33507 22063 33513
rect 22005 33473 22017 33507
rect 22051 33504 22063 33507
rect 22572 33504 22600 33544
rect 23124 33516 23152 33544
rect 23934 33532 23940 33584
rect 23992 33572 23998 33584
rect 24302 33572 24308 33584
rect 23992 33544 24308 33572
rect 23992 33532 23998 33544
rect 24302 33532 24308 33544
rect 24360 33532 24366 33584
rect 24394 33532 24400 33584
rect 24452 33572 24458 33584
rect 28920 33581 28948 33612
rect 29730 33600 29736 33612
rect 29788 33600 29794 33652
rect 25041 33575 25099 33581
rect 25041 33572 25053 33575
rect 24452 33544 25053 33572
rect 24452 33532 24458 33544
rect 25041 33541 25053 33544
rect 25087 33541 25099 33575
rect 25041 33535 25099 33541
rect 28905 33575 28963 33581
rect 28905 33541 28917 33575
rect 28951 33541 28963 33575
rect 28905 33535 28963 33541
rect 28994 33532 29000 33584
rect 29052 33572 29058 33584
rect 29052 33544 29097 33572
rect 29052 33532 29058 33544
rect 22051 33476 22600 33504
rect 22649 33507 22707 33513
rect 22051 33473 22063 33476
rect 22005 33467 22063 33473
rect 22649 33473 22661 33507
rect 22695 33504 22707 33507
rect 22738 33504 22744 33516
rect 22695 33476 22744 33504
rect 22695 33473 22707 33476
rect 22649 33467 22707 33473
rect 22738 33464 22744 33476
rect 22796 33464 22802 33516
rect 23106 33464 23112 33516
rect 23164 33504 23170 33516
rect 23385 33507 23443 33513
rect 23385 33504 23397 33507
rect 23164 33476 23397 33504
rect 23164 33464 23170 33476
rect 23385 33473 23397 33476
rect 23431 33504 23443 33507
rect 23474 33504 23480 33516
rect 23431 33476 23480 33504
rect 23431 33473 23443 33476
rect 23385 33467 23443 33473
rect 23474 33464 23480 33476
rect 23532 33464 23538 33516
rect 24026 33504 24032 33516
rect 23987 33476 24032 33504
rect 24026 33464 24032 33476
rect 24084 33464 24090 33516
rect 26605 33507 26663 33513
rect 26605 33473 26617 33507
rect 26651 33473 26663 33507
rect 26605 33467 26663 33473
rect 22922 33436 22928 33448
rect 18340 33408 22928 33436
rect 22922 33396 22928 33408
rect 22980 33396 22986 33448
rect 24950 33427 25008 33433
rect 24950 33393 24962 33427
rect 24996 33424 25008 33427
rect 25038 33424 25044 33448
rect 24996 33396 25044 33424
rect 25096 33396 25102 33448
rect 25958 33436 25964 33448
rect 25919 33408 25964 33436
rect 25958 33396 25964 33408
rect 26016 33396 26022 33448
rect 26620 33436 26648 33467
rect 26786 33464 26792 33516
rect 26844 33504 26850 33516
rect 27157 33507 27215 33513
rect 27157 33504 27169 33507
rect 26844 33476 27169 33504
rect 26844 33464 26850 33476
rect 27157 33473 27169 33476
rect 27203 33473 27215 33507
rect 27157 33467 27215 33473
rect 27246 33464 27252 33516
rect 27304 33504 27310 33516
rect 27801 33507 27859 33513
rect 27801 33504 27813 33507
rect 27304 33476 27813 33504
rect 27304 33464 27310 33476
rect 27801 33473 27813 33476
rect 27847 33473 27859 33507
rect 27801 33467 27859 33473
rect 27890 33436 27896 33448
rect 26620 33408 27896 33436
rect 27890 33396 27896 33408
rect 27948 33396 27954 33448
rect 29178 33436 29184 33448
rect 29139 33408 29184 33436
rect 29178 33396 29184 33408
rect 29236 33396 29242 33448
rect 24996 33393 25008 33396
rect 24950 33387 25008 33393
rect 22097 33371 22155 33377
rect 22097 33368 22109 33371
rect 15160 33340 17080 33368
rect 18340 33340 22109 33368
rect 15160 33328 15166 33340
rect 4249 33303 4307 33309
rect 4249 33269 4261 33303
rect 4295 33300 4307 33303
rect 4614 33300 4620 33312
rect 4295 33272 4620 33300
rect 4295 33269 4307 33272
rect 4249 33263 4307 33269
rect 4614 33260 4620 33272
rect 4672 33260 4678 33312
rect 4706 33260 4712 33312
rect 4764 33300 4770 33312
rect 5077 33303 5135 33309
rect 5077 33300 5089 33303
rect 4764 33272 5089 33300
rect 4764 33260 4770 33272
rect 5077 33269 5089 33272
rect 5123 33269 5135 33303
rect 5077 33263 5135 33269
rect 15654 33260 15660 33312
rect 15712 33300 15718 33312
rect 18340 33300 18368 33340
rect 22097 33337 22109 33340
rect 22143 33337 22155 33371
rect 22097 33331 22155 33337
rect 27249 33371 27307 33377
rect 27249 33337 27261 33371
rect 27295 33368 27307 33371
rect 28074 33368 28080 33380
rect 27295 33340 28080 33368
rect 27295 33337 27307 33340
rect 27249 33331 27307 33337
rect 28074 33328 28080 33340
rect 28132 33328 28138 33380
rect 15712 33272 18368 33300
rect 15712 33260 15718 33272
rect 18506 33260 18512 33312
rect 18564 33300 18570 33312
rect 18693 33303 18751 33309
rect 18693 33300 18705 33303
rect 18564 33272 18705 33300
rect 18564 33260 18570 33272
rect 18693 33269 18705 33272
rect 18739 33300 18751 33303
rect 22554 33300 22560 33312
rect 18739 33272 22560 33300
rect 18739 33269 18751 33272
rect 18693 33263 18751 33269
rect 22554 33260 22560 33272
rect 22612 33260 22618 33312
rect 22646 33260 22652 33312
rect 22704 33300 22710 33312
rect 22741 33303 22799 33309
rect 22741 33300 22753 33303
rect 22704 33272 22753 33300
rect 22704 33260 22710 33272
rect 22741 33269 22753 33272
rect 22787 33269 22799 33303
rect 22741 33263 22799 33269
rect 24121 33303 24179 33309
rect 24121 33269 24133 33303
rect 24167 33300 24179 33303
rect 24854 33300 24860 33312
rect 24167 33272 24860 33300
rect 24167 33269 24179 33272
rect 24121 33263 24179 33269
rect 24854 33260 24860 33272
rect 24912 33260 24918 33312
rect 27614 33260 27620 33312
rect 27672 33300 27678 33312
rect 27893 33303 27951 33309
rect 27893 33300 27905 33303
rect 27672 33272 27905 33300
rect 27672 33260 27678 33272
rect 27893 33269 27905 33272
rect 27939 33269 27951 33303
rect 27893 33263 27951 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1844 33099 1902 33105
rect 1844 33065 1856 33099
rect 1890 33096 1902 33099
rect 4525 33099 4583 33105
rect 1890 33068 4476 33096
rect 1890 33065 1902 33068
rect 1844 33059 1902 33065
rect 4448 33028 4476 33068
rect 4525 33065 4537 33099
rect 4571 33096 4583 33099
rect 4798 33096 4804 33108
rect 4571 33068 4804 33096
rect 4571 33065 4583 33068
rect 4525 33059 4583 33065
rect 4798 33056 4804 33068
rect 4856 33056 4862 33108
rect 14366 33096 14372 33108
rect 14327 33068 14372 33096
rect 14366 33056 14372 33068
rect 14424 33056 14430 33108
rect 18966 33096 18972 33108
rect 14476 33068 18972 33096
rect 6822 33028 6828 33040
rect 4448 33000 6828 33028
rect 6822 32988 6828 33000
rect 6880 32988 6886 33040
rect 13998 32988 14004 33040
rect 14056 33028 14062 33040
rect 14476 33028 14504 33068
rect 18966 33056 18972 33068
rect 19024 33056 19030 33108
rect 19150 33056 19156 33108
rect 19208 33096 19214 33108
rect 20441 33099 20499 33105
rect 20441 33096 20453 33099
rect 19208 33068 20453 33096
rect 19208 33056 19214 33068
rect 20441 33065 20453 33068
rect 20487 33065 20499 33099
rect 23934 33096 23940 33108
rect 23895 33068 23940 33096
rect 20441 33059 20499 33065
rect 23934 33056 23940 33068
rect 23992 33056 23998 33108
rect 27430 33096 27436 33108
rect 24044 33068 27436 33096
rect 14056 33000 14504 33028
rect 14568 33000 16988 33028
rect 14056 32988 14062 33000
rect 1581 32963 1639 32969
rect 1581 32929 1593 32963
rect 1627 32960 1639 32963
rect 2590 32960 2596 32972
rect 1627 32932 2596 32960
rect 1627 32929 1639 32932
rect 1581 32923 1639 32929
rect 2590 32920 2596 32932
rect 2648 32920 2654 32972
rect 5534 32960 5540 32972
rect 5495 32932 5540 32960
rect 5534 32920 5540 32932
rect 5592 32920 5598 32972
rect 9953 32963 10011 32969
rect 9953 32929 9965 32963
rect 9999 32960 10011 32963
rect 14182 32960 14188 32972
rect 9999 32932 14188 32960
rect 9999 32929 10011 32932
rect 9953 32923 10011 32929
rect 14182 32920 14188 32932
rect 14240 32920 14246 32972
rect 14568 32960 14596 33000
rect 16758 32960 16764 32972
rect 14292 32932 14596 32960
rect 14660 32932 16764 32960
rect 4706 32892 4712 32904
rect 4667 32864 4712 32892
rect 4706 32852 4712 32864
rect 4764 32852 4770 32904
rect 6178 32852 6184 32904
rect 6236 32892 6242 32904
rect 6822 32892 6828 32904
rect 6236 32864 6281 32892
rect 6783 32864 6828 32892
rect 6236 32852 6242 32864
rect 6822 32852 6828 32864
rect 6880 32852 6886 32904
rect 7285 32895 7343 32901
rect 7285 32861 7297 32895
rect 7331 32861 7343 32895
rect 7285 32855 7343 32861
rect 2866 32784 2872 32836
rect 2924 32784 2930 32836
rect 5629 32827 5687 32833
rect 5629 32793 5641 32827
rect 5675 32793 5687 32827
rect 7300 32824 7328 32855
rect 8938 32852 8944 32904
rect 8996 32892 9002 32904
rect 9677 32895 9735 32901
rect 9677 32892 9689 32895
rect 8996 32864 9689 32892
rect 8996 32852 9002 32864
rect 9677 32861 9689 32864
rect 9723 32861 9735 32895
rect 9677 32855 9735 32861
rect 11422 32852 11428 32904
rect 11480 32892 11486 32904
rect 14292 32901 14320 32932
rect 11701 32895 11759 32901
rect 11701 32892 11713 32895
rect 11480 32864 11713 32892
rect 11480 32852 11486 32864
rect 11701 32861 11713 32864
rect 11747 32861 11759 32895
rect 11701 32855 11759 32861
rect 14277 32895 14335 32901
rect 14277 32861 14289 32895
rect 14323 32861 14335 32895
rect 14277 32855 14335 32861
rect 10226 32824 10232 32836
rect 7300 32796 10232 32824
rect 5629 32787 5687 32793
rect 3329 32759 3387 32765
rect 3329 32725 3341 32759
rect 3375 32756 3387 32759
rect 4890 32756 4896 32768
rect 3375 32728 4896 32756
rect 3375 32725 3387 32728
rect 3329 32719 3387 32725
rect 4890 32716 4896 32728
rect 4948 32716 4954 32768
rect 5644 32756 5672 32787
rect 10226 32784 10232 32796
rect 10284 32784 10290 32836
rect 11606 32824 11612 32836
rect 11178 32796 11612 32824
rect 11606 32784 11612 32796
rect 11664 32784 11670 32836
rect 14660 32824 14688 32932
rect 16758 32920 16764 32932
rect 16816 32920 16822 32972
rect 16960 32960 16988 33000
rect 18874 32988 18880 33040
rect 18932 33028 18938 33040
rect 19426 33028 19432 33040
rect 18932 33000 19432 33028
rect 18932 32988 18938 33000
rect 19426 32988 19432 33000
rect 19484 32988 19490 33040
rect 20622 32988 20628 33040
rect 20680 33028 20686 33040
rect 21542 33028 21548 33040
rect 20680 33000 21548 33028
rect 20680 32988 20686 33000
rect 21542 32988 21548 33000
rect 21600 33028 21606 33040
rect 23198 33028 23204 33040
rect 21600 33000 23204 33028
rect 21600 32988 21606 33000
rect 23198 32988 23204 33000
rect 23256 32988 23262 33040
rect 24044 33028 24072 33068
rect 27430 33056 27436 33068
rect 27488 33056 27494 33108
rect 23860 33000 24072 33028
rect 16960 32932 18828 32960
rect 16850 32892 16856 32904
rect 15948 32864 16856 32892
rect 15948 32836 15976 32864
rect 16850 32852 16856 32864
rect 16908 32852 16914 32904
rect 18690 32892 18696 32904
rect 18262 32864 18696 32892
rect 18690 32852 18696 32864
rect 18748 32852 18754 32904
rect 12406 32796 14688 32824
rect 15197 32827 15255 32833
rect 6641 32759 6699 32765
rect 6641 32756 6653 32759
rect 5644 32728 6653 32756
rect 6641 32725 6653 32728
rect 6687 32725 6699 32759
rect 6641 32719 6699 32725
rect 6914 32716 6920 32768
rect 6972 32756 6978 32768
rect 7377 32759 7435 32765
rect 7377 32756 7389 32759
rect 6972 32728 7389 32756
rect 6972 32716 6978 32728
rect 7377 32725 7389 32728
rect 7423 32725 7435 32759
rect 7377 32719 7435 32725
rect 7558 32716 7564 32768
rect 7616 32756 7622 32768
rect 12406 32756 12434 32796
rect 15197 32793 15209 32827
rect 15243 32824 15255 32827
rect 15378 32824 15384 32836
rect 15243 32796 15384 32824
rect 15243 32793 15255 32796
rect 15197 32787 15255 32793
rect 15378 32784 15384 32796
rect 15436 32784 15442 32836
rect 15930 32824 15936 32836
rect 15891 32796 15936 32824
rect 15930 32784 15936 32796
rect 15988 32784 15994 32836
rect 16574 32784 16580 32836
rect 16632 32824 16638 32836
rect 17034 32824 17040 32836
rect 16632 32796 17040 32824
rect 16632 32784 16638 32796
rect 17034 32784 17040 32796
rect 17092 32784 17098 32836
rect 17129 32827 17187 32833
rect 17129 32793 17141 32827
rect 17175 32793 17187 32827
rect 18800 32824 18828 32932
rect 19610 32920 19616 32972
rect 19668 32960 19674 32972
rect 23293 32963 23351 32969
rect 23293 32960 23305 32963
rect 19668 32932 23305 32960
rect 19668 32920 19674 32932
rect 23293 32929 23305 32932
rect 23339 32929 23351 32963
rect 23293 32923 23351 32929
rect 18874 32852 18880 32904
rect 18932 32892 18938 32904
rect 19426 32892 19432 32904
rect 18932 32864 19432 32892
rect 18932 32852 18938 32864
rect 19426 32852 19432 32864
rect 19484 32852 19490 32904
rect 20349 32895 20407 32901
rect 20349 32861 20361 32895
rect 20395 32892 20407 32895
rect 20530 32892 20536 32904
rect 20395 32864 20536 32892
rect 20395 32861 20407 32864
rect 20349 32855 20407 32861
rect 20530 32852 20536 32864
rect 20588 32852 20594 32904
rect 22370 32852 22376 32904
rect 22428 32892 22434 32904
rect 22557 32895 22615 32901
rect 22557 32892 22569 32895
rect 22428 32864 22569 32892
rect 22428 32852 22434 32864
rect 22557 32861 22569 32864
rect 22603 32861 22615 32895
rect 22557 32855 22615 32861
rect 22922 32852 22928 32904
rect 22980 32892 22986 32904
rect 23106 32892 23112 32904
rect 22980 32864 23112 32892
rect 22980 32852 22986 32864
rect 23106 32852 23112 32864
rect 23164 32892 23170 32904
rect 23860 32901 23888 33000
rect 24118 32988 24124 33040
rect 24176 33028 24182 33040
rect 24176 33000 28856 33028
rect 24176 32988 24182 33000
rect 24302 32920 24308 32972
rect 24360 32960 24366 32972
rect 24673 32963 24731 32969
rect 24673 32960 24685 32963
rect 24360 32932 24685 32960
rect 24360 32920 24366 32932
rect 24673 32929 24685 32932
rect 24719 32929 24731 32963
rect 25130 32960 25136 32972
rect 25091 32932 25136 32960
rect 24673 32923 24731 32929
rect 25130 32920 25136 32932
rect 25188 32920 25194 32972
rect 26789 32963 26847 32969
rect 26789 32929 26801 32963
rect 26835 32960 26847 32963
rect 26970 32960 26976 32972
rect 26835 32932 26976 32960
rect 26835 32929 26847 32932
rect 26789 32923 26847 32929
rect 26970 32920 26976 32932
rect 27028 32920 27034 32972
rect 27709 32963 27767 32969
rect 27709 32929 27721 32963
rect 27755 32960 27767 32963
rect 27755 32932 28764 32960
rect 27755 32929 27767 32932
rect 27709 32923 27767 32929
rect 23201 32895 23259 32901
rect 23201 32892 23213 32895
rect 23164 32864 23213 32892
rect 23164 32852 23170 32864
rect 23201 32861 23213 32864
rect 23247 32861 23259 32895
rect 23201 32855 23259 32861
rect 23845 32895 23903 32901
rect 23845 32861 23857 32895
rect 23891 32861 23903 32895
rect 23845 32855 23903 32861
rect 20254 32824 20260 32836
rect 18800 32796 20260 32824
rect 17129 32787 17187 32793
rect 7616 32728 12434 32756
rect 7616 32716 7622 32728
rect 13078 32716 13084 32768
rect 13136 32756 13142 32768
rect 15102 32756 15108 32768
rect 13136 32728 15108 32756
rect 13136 32716 13142 32728
rect 15102 32716 15108 32728
rect 15160 32716 15166 32768
rect 15286 32716 15292 32768
rect 15344 32756 15350 32768
rect 17144 32756 17172 32787
rect 20254 32784 20260 32796
rect 20312 32784 20318 32836
rect 21082 32824 21088 32836
rect 21043 32796 21088 32824
rect 21082 32784 21088 32796
rect 21140 32784 21146 32836
rect 21174 32784 21180 32836
rect 21232 32824 21238 32836
rect 22094 32824 22100 32836
rect 21232 32796 21277 32824
rect 22055 32796 22100 32824
rect 21232 32784 21238 32796
rect 22094 32784 22100 32796
rect 22152 32784 22158 32836
rect 22649 32827 22707 32833
rect 22649 32793 22661 32827
rect 22695 32824 22707 32827
rect 24765 32827 24823 32833
rect 22695 32796 24624 32824
rect 22695 32793 22707 32796
rect 22649 32787 22707 32793
rect 22002 32756 22008 32768
rect 15344 32728 22008 32756
rect 15344 32716 15350 32728
rect 22002 32716 22008 32728
rect 22060 32716 22066 32768
rect 22186 32716 22192 32768
rect 22244 32756 22250 32768
rect 23658 32756 23664 32768
rect 22244 32728 23664 32756
rect 22244 32716 22250 32728
rect 23658 32716 23664 32728
rect 23716 32756 23722 32768
rect 24486 32756 24492 32768
rect 23716 32728 24492 32756
rect 23716 32716 23722 32728
rect 24486 32716 24492 32728
rect 24544 32716 24550 32768
rect 24596 32756 24624 32796
rect 24765 32793 24777 32827
rect 24811 32793 24823 32827
rect 24765 32787 24823 32793
rect 24780 32756 24808 32787
rect 25406 32784 25412 32836
rect 25464 32824 25470 32836
rect 26145 32827 26203 32833
rect 26145 32824 26157 32827
rect 25464 32796 26157 32824
rect 25464 32784 25470 32796
rect 26145 32793 26157 32796
rect 26191 32793 26203 32827
rect 26145 32787 26203 32793
rect 26237 32827 26295 32833
rect 26237 32793 26249 32827
rect 26283 32793 26295 32827
rect 26237 32787 26295 32793
rect 27801 32827 27859 32833
rect 27801 32793 27813 32827
rect 27847 32793 27859 32827
rect 28350 32824 28356 32836
rect 28311 32796 28356 32824
rect 27801 32787 27859 32793
rect 24596 32728 24808 32756
rect 24946 32716 24952 32768
rect 25004 32756 25010 32768
rect 25498 32756 25504 32768
rect 25004 32728 25504 32756
rect 25004 32716 25010 32728
rect 25498 32716 25504 32728
rect 25556 32716 25562 32768
rect 26252 32756 26280 32787
rect 27614 32756 27620 32768
rect 26252 32728 27620 32756
rect 27614 32716 27620 32728
rect 27672 32716 27678 32768
rect 27816 32756 27844 32787
rect 28350 32784 28356 32796
rect 28408 32784 28414 32836
rect 28736 32824 28764 32932
rect 28828 32901 28856 33000
rect 28813 32895 28871 32901
rect 28813 32861 28825 32895
rect 28859 32861 28871 32895
rect 28813 32855 28871 32861
rect 29822 32824 29828 32836
rect 28736 32796 29828 32824
rect 29822 32784 29828 32796
rect 29880 32784 29886 32836
rect 38102 32824 38108 32836
rect 38063 32796 38108 32824
rect 38102 32784 38108 32796
rect 38160 32784 38166 32836
rect 28905 32759 28963 32765
rect 28905 32756 28917 32759
rect 27816 32728 28917 32756
rect 28905 32725 28917 32728
rect 28951 32725 28963 32759
rect 28905 32719 28963 32725
rect 37826 32716 37832 32768
rect 37884 32756 37890 32768
rect 38197 32759 38255 32765
rect 38197 32756 38209 32759
rect 37884 32728 38209 32756
rect 37884 32716 37890 32728
rect 38197 32725 38209 32728
rect 38243 32725 38255 32759
rect 38197 32719 38255 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 5721 32555 5779 32561
rect 5721 32521 5733 32555
rect 5767 32552 5779 32555
rect 7558 32552 7564 32564
rect 5767 32524 7564 32552
rect 5767 32521 5779 32524
rect 5721 32515 5779 32521
rect 7558 32512 7564 32524
rect 7616 32512 7622 32564
rect 15930 32552 15936 32564
rect 13280 32524 15936 32552
rect 7466 32484 7472 32496
rect 7427 32456 7472 32484
rect 7466 32444 7472 32456
rect 7524 32444 7530 32496
rect 13078 32484 13084 32496
rect 10442 32456 13084 32484
rect 13078 32444 13084 32456
rect 13136 32444 13142 32496
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32385 1639 32419
rect 1581 32379 1639 32385
rect 1596 32348 1624 32379
rect 2038 32376 2044 32428
rect 2096 32416 2102 32428
rect 2317 32419 2375 32425
rect 2317 32416 2329 32419
rect 2096 32388 2329 32416
rect 2096 32376 2102 32388
rect 2317 32385 2329 32388
rect 2363 32416 2375 32419
rect 5629 32419 5687 32425
rect 5629 32416 5641 32419
rect 2363 32388 5641 32416
rect 2363 32385 2375 32388
rect 2317 32379 2375 32385
rect 5629 32385 5641 32388
rect 5675 32385 5687 32419
rect 5629 32379 5687 32385
rect 6641 32419 6699 32425
rect 6641 32385 6653 32419
rect 6687 32385 6699 32419
rect 6641 32379 6699 32385
rect 6546 32348 6552 32360
rect 1596 32320 6552 32348
rect 6546 32308 6552 32320
rect 6604 32308 6610 32360
rect 1762 32212 1768 32224
rect 1723 32184 1768 32212
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 2409 32215 2467 32221
rect 2409 32181 2421 32215
rect 2455 32212 2467 32215
rect 5626 32212 5632 32224
rect 2455 32184 5632 32212
rect 2455 32181 2467 32184
rect 2409 32175 2467 32181
rect 5626 32172 5632 32184
rect 5684 32172 5690 32224
rect 6656 32212 6684 32379
rect 8294 32376 8300 32428
rect 8352 32416 8358 32428
rect 8938 32416 8944 32428
rect 8352 32388 8944 32416
rect 8352 32376 8358 32388
rect 8938 32376 8944 32388
rect 8996 32376 9002 32428
rect 13280 32425 13308 32524
rect 15930 32512 15936 32524
rect 15988 32512 15994 32564
rect 18874 32552 18880 32564
rect 17144 32524 18880 32552
rect 13538 32484 13544 32496
rect 13499 32456 13544 32484
rect 13538 32444 13544 32456
rect 13596 32444 13602 32496
rect 15286 32484 15292 32496
rect 15247 32456 15292 32484
rect 15286 32444 15292 32456
rect 15344 32444 15350 32496
rect 13265 32419 13323 32425
rect 13265 32385 13277 32419
rect 13311 32385 13323 32419
rect 15654 32416 15660 32428
rect 14674 32388 15660 32416
rect 13265 32379 13323 32385
rect 15654 32376 15660 32388
rect 15712 32376 15718 32428
rect 15948 32416 15976 32512
rect 17144 32493 17172 32524
rect 18874 32512 18880 32524
rect 18932 32512 18938 32564
rect 18966 32512 18972 32564
rect 19024 32552 19030 32564
rect 26326 32552 26332 32564
rect 19024 32524 20668 32552
rect 26287 32524 26332 32552
rect 19024 32512 19030 32524
rect 17129 32487 17187 32493
rect 17129 32453 17141 32487
rect 17175 32453 17187 32487
rect 19242 32484 19248 32496
rect 18354 32456 19248 32484
rect 17129 32447 17187 32453
rect 19242 32444 19248 32456
rect 19300 32444 19306 32496
rect 19978 32444 19984 32496
rect 20036 32484 20042 32496
rect 20640 32484 20668 32524
rect 26326 32512 26332 32524
rect 26384 32512 26390 32564
rect 27249 32555 27307 32561
rect 27249 32521 27261 32555
rect 27295 32552 27307 32555
rect 27798 32552 27804 32564
rect 27295 32524 27804 32552
rect 27295 32521 27307 32524
rect 27249 32515 27307 32521
rect 27798 32512 27804 32524
rect 27856 32512 27862 32564
rect 27893 32555 27951 32561
rect 27893 32521 27905 32555
rect 27939 32552 27951 32555
rect 28994 32552 29000 32564
rect 27939 32524 29000 32552
rect 27939 32521 27951 32524
rect 27893 32515 27951 32521
rect 28994 32512 29000 32524
rect 29052 32512 29058 32564
rect 33042 32512 33048 32564
rect 33100 32552 33106 32564
rect 38105 32555 38163 32561
rect 38105 32552 38117 32555
rect 33100 32524 38117 32552
rect 33100 32512 33106 32524
rect 38105 32521 38117 32524
rect 38151 32521 38163 32555
rect 38105 32515 38163 32521
rect 22738 32484 22744 32496
rect 20036 32456 20576 32484
rect 20640 32456 22744 32484
rect 20036 32444 20042 32456
rect 20548 32428 20576 32456
rect 22738 32444 22744 32456
rect 22796 32444 22802 32496
rect 23290 32484 23296 32496
rect 23251 32456 23296 32484
rect 23290 32444 23296 32456
rect 23348 32444 23354 32496
rect 24854 32493 24860 32496
rect 24850 32447 24860 32493
rect 24912 32484 24918 32496
rect 24912 32456 24950 32484
rect 24854 32444 24860 32447
rect 24912 32444 24918 32456
rect 16758 32416 16764 32428
rect 15948 32388 16764 32416
rect 16758 32376 16764 32388
rect 16816 32416 16822 32428
rect 16853 32419 16911 32425
rect 16853 32416 16865 32419
rect 16816 32388 16865 32416
rect 16816 32376 16822 32388
rect 16853 32385 16865 32388
rect 16899 32385 16911 32419
rect 16853 32379 16911 32385
rect 18506 32376 18512 32428
rect 18564 32416 18570 32428
rect 19705 32419 19763 32425
rect 18564 32388 18828 32416
rect 18564 32376 18570 32388
rect 9217 32351 9275 32357
rect 9217 32317 9229 32351
rect 9263 32348 9275 32351
rect 9263 32320 18644 32348
rect 9263 32317 9275 32320
rect 9217 32311 9275 32317
rect 18616 32289 18644 32320
rect 18601 32283 18659 32289
rect 18601 32249 18613 32283
rect 18647 32280 18659 32283
rect 18690 32280 18696 32292
rect 18647 32252 18696 32280
rect 18647 32249 18659 32252
rect 18601 32243 18659 32249
rect 18690 32240 18696 32252
rect 18748 32240 18754 32292
rect 18800 32280 18828 32388
rect 19705 32385 19717 32419
rect 19751 32385 19763 32419
rect 19705 32379 19763 32385
rect 18966 32308 18972 32360
rect 19024 32348 19030 32360
rect 19720 32348 19748 32379
rect 20254 32376 20260 32428
rect 20312 32416 20318 32428
rect 20349 32419 20407 32425
rect 20349 32416 20361 32419
rect 20312 32388 20361 32416
rect 20312 32376 20318 32388
rect 20349 32385 20361 32388
rect 20395 32385 20407 32419
rect 20349 32379 20407 32385
rect 20530 32376 20536 32428
rect 20588 32416 20594 32428
rect 20993 32419 21051 32425
rect 20993 32416 21005 32419
rect 20588 32388 21005 32416
rect 20588 32376 20594 32388
rect 20993 32385 21005 32388
rect 21039 32416 21051 32419
rect 21450 32416 21456 32428
rect 21039 32388 21456 32416
rect 21039 32385 21051 32388
rect 20993 32379 21051 32385
rect 21450 32376 21456 32388
rect 21508 32376 21514 32428
rect 21726 32376 21732 32428
rect 21784 32416 21790 32428
rect 21910 32416 21916 32428
rect 21784 32388 21916 32416
rect 21784 32376 21790 32388
rect 21910 32376 21916 32388
rect 21968 32416 21974 32428
rect 22005 32419 22063 32425
rect 22005 32416 22017 32419
rect 21968 32388 22017 32416
rect 21968 32376 21974 32388
rect 22005 32385 22017 32388
rect 22051 32385 22063 32419
rect 22005 32379 22063 32385
rect 22462 32376 22468 32428
rect 22520 32416 22526 32428
rect 22922 32416 22928 32428
rect 22520 32388 22928 32416
rect 22520 32376 22526 32388
rect 22922 32376 22928 32388
rect 22980 32376 22986 32428
rect 26237 32419 26295 32425
rect 26237 32385 26249 32419
rect 26283 32385 26295 32419
rect 26237 32379 26295 32385
rect 19024 32320 19748 32348
rect 19797 32351 19855 32357
rect 19024 32308 19030 32320
rect 19797 32317 19809 32351
rect 19843 32348 19855 32351
rect 22554 32348 22560 32360
rect 19843 32320 22560 32348
rect 19843 32317 19855 32320
rect 19797 32311 19855 32317
rect 22554 32308 22560 32320
rect 22612 32308 22618 32360
rect 23198 32348 23204 32360
rect 23159 32320 23204 32348
rect 23198 32308 23204 32320
rect 23256 32308 23262 32360
rect 24213 32351 24271 32357
rect 24213 32317 24225 32351
rect 24259 32317 24271 32351
rect 24213 32311 24271 32317
rect 24765 32351 24823 32357
rect 24765 32317 24777 32351
rect 24811 32348 24823 32351
rect 24946 32348 24952 32360
rect 24811 32320 24952 32348
rect 24811 32317 24823 32320
rect 24765 32311 24823 32317
rect 24118 32280 24124 32292
rect 18800 32252 24124 32280
rect 24118 32240 24124 32252
rect 24176 32240 24182 32292
rect 24228 32280 24256 32311
rect 24946 32308 24952 32320
rect 25004 32308 25010 32360
rect 25041 32351 25099 32357
rect 25041 32317 25053 32351
rect 25087 32317 25099 32351
rect 26252 32348 26280 32379
rect 26970 32376 26976 32428
rect 27028 32416 27034 32428
rect 27157 32419 27215 32425
rect 27157 32416 27169 32419
rect 27028 32388 27169 32416
rect 27028 32376 27034 32388
rect 27157 32385 27169 32388
rect 27203 32385 27215 32419
rect 27157 32379 27215 32385
rect 27614 32376 27620 32428
rect 27672 32416 27678 32428
rect 27801 32419 27859 32425
rect 27801 32416 27813 32419
rect 27672 32388 27813 32416
rect 27672 32376 27678 32388
rect 27801 32385 27813 32388
rect 27847 32385 27859 32419
rect 38286 32416 38292 32428
rect 38247 32388 38292 32416
rect 27801 32379 27859 32385
rect 38286 32376 38292 32388
rect 38344 32376 38350 32428
rect 27522 32348 27528 32360
rect 26252 32320 27528 32348
rect 25041 32311 25099 32317
rect 24854 32280 24860 32292
rect 24228 32252 24860 32280
rect 24854 32240 24860 32252
rect 24912 32240 24918 32292
rect 10226 32212 10232 32224
rect 6656 32184 10232 32212
rect 10226 32172 10232 32184
rect 10284 32172 10290 32224
rect 10686 32212 10692 32224
rect 10599 32184 10692 32212
rect 10686 32172 10692 32184
rect 10744 32212 10750 32224
rect 18966 32212 18972 32224
rect 10744 32184 18972 32212
rect 10744 32172 10750 32184
rect 18966 32172 18972 32184
rect 19024 32172 19030 32224
rect 19334 32172 19340 32224
rect 19392 32212 19398 32224
rect 20441 32215 20499 32221
rect 20441 32212 20453 32215
rect 19392 32184 20453 32212
rect 19392 32172 19398 32184
rect 20441 32181 20453 32184
rect 20487 32181 20499 32215
rect 21082 32212 21088 32224
rect 21043 32184 21088 32212
rect 20441 32175 20499 32181
rect 21082 32172 21088 32184
rect 21140 32172 21146 32224
rect 22094 32172 22100 32224
rect 22152 32212 22158 32224
rect 22152 32184 22197 32212
rect 22152 32172 22158 32184
rect 23106 32172 23112 32224
rect 23164 32212 23170 32224
rect 25056 32212 25084 32311
rect 27522 32308 27528 32320
rect 27580 32308 27586 32360
rect 23164 32184 25084 32212
rect 23164 32172 23170 32184
rect 25498 32172 25504 32224
rect 25556 32212 25562 32224
rect 28534 32212 28540 32224
rect 25556 32184 28540 32212
rect 25556 32172 25562 32184
rect 28534 32172 28540 32184
rect 28592 32172 28598 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 2958 32008 2964 32020
rect 2919 31980 2964 32008
rect 2958 31968 2964 31980
rect 3016 31968 3022 32020
rect 4065 32011 4123 32017
rect 4065 31977 4077 32011
rect 4111 32008 4123 32011
rect 4111 31980 6776 32008
rect 4111 31977 4123 31980
rect 4065 31971 4123 31977
rect 6748 31940 6776 31980
rect 6822 31968 6828 32020
rect 6880 32008 6886 32020
rect 7561 32011 7619 32017
rect 7561 32008 7573 32011
rect 6880 31980 7573 32008
rect 6880 31968 6886 31980
rect 7561 31977 7573 31980
rect 7607 31977 7619 32011
rect 7561 31971 7619 31977
rect 12056 32011 12114 32017
rect 12056 31977 12068 32011
rect 12102 32008 12114 32011
rect 12710 32008 12716 32020
rect 12102 31980 12716 32008
rect 12102 31977 12114 31980
rect 12056 31971 12114 31977
rect 12710 31968 12716 31980
rect 12768 31968 12774 32020
rect 15930 31968 15936 32020
rect 15988 32008 15994 32020
rect 22094 32008 22100 32020
rect 15988 31980 22100 32008
rect 15988 31968 15994 31980
rect 22094 31968 22100 31980
rect 22152 31968 22158 32020
rect 23290 31968 23296 32020
rect 23348 32008 23354 32020
rect 24673 32011 24731 32017
rect 24673 32008 24685 32011
rect 23348 31980 24685 32008
rect 23348 31968 23354 31980
rect 24673 31977 24685 31980
rect 24719 31977 24731 32011
rect 24673 31971 24731 31977
rect 10318 31940 10324 31952
rect 6748 31912 10324 31940
rect 10318 31900 10324 31912
rect 10376 31900 10382 31952
rect 15378 31940 15384 31952
rect 13188 31912 15384 31940
rect 2682 31832 2688 31884
rect 2740 31872 2746 31884
rect 4154 31872 4160 31884
rect 2740 31844 4160 31872
rect 2740 31832 2746 31844
rect 4154 31832 4160 31844
rect 4212 31872 4218 31884
rect 5077 31875 5135 31881
rect 5077 31872 5089 31875
rect 4212 31844 5089 31872
rect 4212 31832 4218 31844
rect 5077 31841 5089 31844
rect 5123 31872 5135 31875
rect 7466 31872 7472 31884
rect 5123 31844 7472 31872
rect 5123 31841 5135 31844
rect 5077 31835 5135 31841
rect 7466 31832 7472 31844
rect 7524 31832 7530 31884
rect 10226 31832 10232 31884
rect 10284 31872 10290 31884
rect 13188 31872 13216 31912
rect 15378 31900 15384 31912
rect 15436 31900 15442 31952
rect 20622 31940 20628 31952
rect 18708 31912 20628 31940
rect 10284 31844 13216 31872
rect 13541 31875 13599 31881
rect 10284 31832 10290 31844
rect 13541 31841 13553 31875
rect 13587 31841 13599 31875
rect 16758 31872 16764 31884
rect 16719 31844 16764 31872
rect 13541 31835 13599 31841
rect 1854 31804 1860 31816
rect 1815 31776 1860 31804
rect 1854 31764 1860 31776
rect 1912 31764 1918 31816
rect 1949 31807 2007 31813
rect 1949 31773 1961 31807
rect 1995 31804 2007 31807
rect 2406 31804 2412 31816
rect 1995 31776 2412 31804
rect 1995 31773 2007 31776
rect 1949 31767 2007 31773
rect 2406 31764 2412 31776
rect 2464 31764 2470 31816
rect 3142 31804 3148 31816
rect 3055 31776 3148 31804
rect 3142 31764 3148 31776
rect 3200 31804 3206 31816
rect 3973 31807 4031 31813
rect 3973 31804 3985 31807
rect 3200 31776 3985 31804
rect 3200 31764 3206 31776
rect 3973 31773 3985 31776
rect 4019 31773 4031 31807
rect 3973 31767 4031 31773
rect 6454 31764 6460 31816
rect 6512 31764 6518 31816
rect 7098 31804 7104 31816
rect 7059 31776 7104 31804
rect 7098 31764 7104 31776
rect 7156 31764 7162 31816
rect 7745 31807 7803 31813
rect 7745 31773 7757 31807
rect 7791 31804 7803 31807
rect 7834 31804 7840 31816
rect 7791 31776 7840 31804
rect 7791 31773 7803 31776
rect 7745 31767 7803 31773
rect 7834 31764 7840 31776
rect 7892 31764 7898 31816
rect 8938 31764 8944 31816
rect 8996 31804 9002 31816
rect 11790 31804 11796 31816
rect 8996 31776 10456 31804
rect 11751 31776 11796 31804
rect 8996 31764 9002 31776
rect 5353 31739 5411 31745
rect 5353 31705 5365 31739
rect 5399 31736 5411 31739
rect 10321 31739 10379 31745
rect 5399 31708 5764 31736
rect 5399 31705 5411 31708
rect 5353 31699 5411 31705
rect 5736 31668 5764 31708
rect 10321 31705 10333 31739
rect 10367 31705 10379 31739
rect 10428 31736 10456 31776
rect 11790 31764 11796 31776
rect 11848 31764 11854 31816
rect 13556 31804 13584 31835
rect 16758 31832 16764 31844
rect 16816 31832 16822 31884
rect 18506 31872 18512 31884
rect 18467 31844 18512 31872
rect 18506 31832 18512 31844
rect 18564 31832 18570 31884
rect 18708 31804 18736 31912
rect 20622 31900 20628 31912
rect 20680 31900 20686 31952
rect 20732 31912 23336 31940
rect 20732 31881 20760 31912
rect 20717 31875 20775 31881
rect 20717 31841 20729 31875
rect 20763 31841 20775 31875
rect 20717 31835 20775 31841
rect 21729 31875 21787 31881
rect 21729 31841 21741 31875
rect 21775 31872 21787 31875
rect 22002 31872 22008 31884
rect 21775 31844 22008 31872
rect 21775 31841 21787 31844
rect 21729 31835 21787 31841
rect 22002 31832 22008 31844
rect 22060 31832 22066 31884
rect 22186 31832 22192 31884
rect 22244 31872 22250 31884
rect 22465 31875 22523 31881
rect 22465 31872 22477 31875
rect 22244 31844 22477 31872
rect 22244 31832 22250 31844
rect 22465 31841 22477 31844
rect 22511 31841 22523 31875
rect 22465 31835 22523 31841
rect 22830 31832 22836 31884
rect 22888 31872 22894 31884
rect 23106 31872 23112 31884
rect 22888 31844 23112 31872
rect 22888 31832 22894 31844
rect 23106 31832 23112 31844
rect 23164 31832 23170 31884
rect 23308 31872 23336 31912
rect 23382 31900 23388 31952
rect 23440 31940 23446 31952
rect 25961 31943 26019 31949
rect 25961 31940 25973 31943
rect 23440 31912 25973 31940
rect 23440 31900 23446 31912
rect 25961 31909 25973 31912
rect 26007 31909 26019 31943
rect 27614 31940 27620 31952
rect 25961 31903 26019 31909
rect 26804 31912 27620 31940
rect 26804 31881 26832 31912
rect 27614 31900 27620 31912
rect 27672 31900 27678 31952
rect 26789 31875 26847 31881
rect 26789 31872 26801 31875
rect 23308 31844 26801 31872
rect 26789 31841 26801 31844
rect 26835 31841 26847 31875
rect 26789 31835 26847 31841
rect 27433 31875 27491 31881
rect 27433 31841 27445 31875
rect 27479 31872 27491 31875
rect 28350 31872 28356 31884
rect 27479 31844 28356 31872
rect 27479 31841 27491 31844
rect 27433 31835 27491 31841
rect 13556 31776 16804 31804
rect 18170 31776 18736 31804
rect 11146 31736 11152 31748
rect 10428 31708 11152 31736
rect 10321 31699 10379 31705
rect 5994 31668 6000 31680
rect 5736 31640 6000 31668
rect 5994 31628 6000 31640
rect 6052 31628 6058 31680
rect 10226 31628 10232 31680
rect 10284 31668 10290 31680
rect 10336 31668 10364 31699
rect 11146 31696 11152 31708
rect 11204 31696 11210 31748
rect 15930 31736 15936 31748
rect 13294 31708 15936 31736
rect 15930 31696 15936 31708
rect 15988 31696 15994 31748
rect 16776 31736 16804 31776
rect 18782 31764 18788 31816
rect 18840 31804 18846 31816
rect 24581 31807 24639 31813
rect 18840 31776 20576 31804
rect 18840 31764 18846 31776
rect 16942 31736 16948 31748
rect 16776 31708 16948 31736
rect 16942 31696 16948 31708
rect 17000 31696 17006 31748
rect 17037 31739 17095 31745
rect 17037 31705 17049 31739
rect 17083 31736 17095 31739
rect 17126 31736 17132 31748
rect 17083 31708 17132 31736
rect 17083 31705 17095 31708
rect 17037 31699 17095 31705
rect 17126 31696 17132 31708
rect 17184 31696 17190 31748
rect 20548 31736 20576 31776
rect 24581 31773 24593 31807
rect 24627 31804 24639 31807
rect 24762 31804 24768 31816
rect 24627 31776 24768 31804
rect 24627 31773 24639 31776
rect 24581 31767 24639 31773
rect 24762 31764 24768 31776
rect 24820 31764 24826 31816
rect 25225 31807 25283 31813
rect 25225 31804 25237 31807
rect 24872 31776 25237 31804
rect 20809 31739 20867 31745
rect 20809 31736 20821 31739
rect 20548 31708 20821 31736
rect 20809 31705 20821 31708
rect 20855 31705 20867 31739
rect 22554 31736 22560 31748
rect 22515 31708 22560 31736
rect 20809 31699 20867 31705
rect 22554 31696 22560 31708
rect 22612 31696 22618 31748
rect 23382 31696 23388 31748
rect 23440 31736 23446 31748
rect 24872 31736 24900 31776
rect 25225 31773 25237 31776
rect 25271 31773 25283 31807
rect 25225 31767 25283 31773
rect 25314 31764 25320 31816
rect 25372 31804 25378 31816
rect 25372 31776 25417 31804
rect 25372 31764 25378 31776
rect 25774 31764 25780 31816
rect 25832 31804 25838 31816
rect 25869 31807 25927 31813
rect 25869 31804 25881 31807
rect 25832 31776 25881 31804
rect 25832 31764 25838 31776
rect 25869 31773 25881 31776
rect 25915 31773 25927 31807
rect 25869 31767 25927 31773
rect 26878 31736 26884 31748
rect 23440 31708 24900 31736
rect 26839 31708 26884 31736
rect 23440 31696 23446 31708
rect 26878 31696 26884 31708
rect 26936 31696 26942 31748
rect 26970 31696 26976 31748
rect 27028 31736 27034 31748
rect 27246 31736 27252 31748
rect 27028 31708 27252 31736
rect 27028 31696 27034 31708
rect 27246 31696 27252 31708
rect 27304 31696 27310 31748
rect 27816 31736 27844 31844
rect 28350 31832 28356 31844
rect 28408 31872 28414 31884
rect 28408 31844 28856 31872
rect 28408 31832 28414 31844
rect 28828 31804 28856 31844
rect 28902 31832 28908 31884
rect 28960 31872 28966 31884
rect 32122 31872 32128 31884
rect 28960 31844 32128 31872
rect 28960 31832 28966 31844
rect 32122 31832 32128 31844
rect 32180 31832 32186 31884
rect 30374 31804 30380 31816
rect 28828 31776 30380 31804
rect 30374 31764 30380 31776
rect 30432 31764 30438 31816
rect 27985 31739 28043 31745
rect 27985 31736 27997 31739
rect 27816 31708 27997 31736
rect 27985 31705 27997 31708
rect 28031 31705 28043 31739
rect 27985 31699 28043 31705
rect 28074 31696 28080 31748
rect 28132 31736 28138 31748
rect 28132 31708 28177 31736
rect 28132 31696 28138 31708
rect 10962 31668 10968 31680
rect 10284 31640 10968 31668
rect 10284 31628 10290 31640
rect 10962 31628 10968 31640
rect 11020 31628 11026 31680
rect 11238 31628 11244 31680
rect 11296 31668 11302 31680
rect 22370 31668 22376 31680
rect 11296 31640 22376 31668
rect 11296 31628 11302 31640
rect 22370 31628 22376 31640
rect 22428 31668 22434 31680
rect 22922 31668 22928 31680
rect 22428 31640 22928 31668
rect 22428 31628 22434 31640
rect 22922 31628 22928 31640
rect 22980 31628 22986 31680
rect 23106 31628 23112 31680
rect 23164 31668 23170 31680
rect 25866 31668 25872 31680
rect 23164 31640 25872 31668
rect 23164 31628 23170 31640
rect 25866 31628 25872 31640
rect 25924 31628 25930 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1581 31467 1639 31473
rect 1581 31433 1593 31467
rect 1627 31464 1639 31467
rect 3142 31464 3148 31476
rect 1627 31436 3148 31464
rect 1627 31433 1639 31436
rect 1581 31427 1639 31433
rect 3142 31424 3148 31436
rect 3200 31424 3206 31476
rect 4062 31464 4068 31476
rect 3988 31436 4068 31464
rect 1762 31328 1768 31340
rect 1723 31300 1768 31328
rect 1762 31288 1768 31300
rect 1820 31288 1826 31340
rect 3329 31331 3387 31337
rect 3329 31297 3341 31331
rect 3375 31328 3387 31331
rect 3418 31328 3424 31340
rect 3375 31300 3424 31328
rect 3375 31297 3387 31300
rect 3329 31291 3387 31297
rect 3418 31288 3424 31300
rect 3476 31288 3482 31340
rect 3988 31337 4016 31436
rect 4062 31424 4068 31436
rect 4120 31424 4126 31476
rect 6546 31424 6552 31476
rect 6604 31464 6610 31476
rect 6733 31467 6791 31473
rect 6733 31464 6745 31467
rect 6604 31436 6745 31464
rect 6604 31424 6610 31436
rect 6733 31433 6745 31436
rect 6779 31433 6791 31467
rect 23106 31464 23112 31476
rect 6733 31427 6791 31433
rect 10980 31436 23112 31464
rect 8294 31396 8300 31408
rect 8128 31368 8300 31396
rect 3973 31331 4031 31337
rect 3973 31297 3985 31331
rect 4019 31297 4031 31331
rect 3973 31291 4031 31297
rect 5350 31288 5356 31340
rect 5408 31288 5414 31340
rect 6914 31328 6920 31340
rect 6875 31300 6920 31328
rect 6914 31288 6920 31300
rect 6972 31288 6978 31340
rect 8128 31337 8156 31368
rect 8294 31356 8300 31368
rect 8352 31356 8358 31408
rect 10980 31396 11008 31436
rect 23106 31424 23112 31436
rect 23164 31424 23170 31476
rect 23201 31467 23259 31473
rect 23201 31433 23213 31467
rect 23247 31464 23259 31467
rect 23566 31464 23572 31476
rect 23247 31436 23572 31464
rect 23247 31433 23259 31436
rect 23201 31427 23259 31433
rect 23566 31424 23572 31436
rect 23624 31424 23630 31476
rect 24394 31424 24400 31476
rect 24452 31464 24458 31476
rect 27249 31467 27307 31473
rect 27249 31464 27261 31467
rect 24452 31436 27261 31464
rect 24452 31424 24458 31436
rect 27249 31433 27261 31436
rect 27295 31433 27307 31467
rect 27249 31427 27307 31433
rect 27801 31467 27859 31473
rect 27801 31433 27813 31467
rect 27847 31464 27859 31467
rect 27890 31464 27896 31476
rect 27847 31436 27896 31464
rect 27847 31433 27859 31436
rect 27801 31427 27859 31433
rect 27890 31424 27896 31436
rect 27948 31424 27954 31476
rect 12342 31396 12348 31408
rect 9614 31368 11008 31396
rect 12303 31368 12348 31396
rect 12342 31356 12348 31368
rect 12400 31356 12406 31408
rect 12434 31356 12440 31408
rect 12492 31396 12498 31408
rect 16117 31399 16175 31405
rect 16117 31396 16129 31399
rect 12492 31368 12834 31396
rect 14016 31368 16129 31396
rect 12492 31356 12498 31368
rect 8113 31331 8171 31337
rect 8113 31297 8125 31331
rect 8159 31297 8171 31331
rect 8113 31291 8171 31297
rect 11790 31288 11796 31340
rect 11848 31328 11854 31340
rect 12069 31331 12127 31337
rect 12069 31328 12081 31331
rect 11848 31300 12081 31328
rect 11848 31288 11854 31300
rect 12069 31297 12081 31300
rect 12115 31297 12127 31331
rect 12069 31291 12127 31297
rect 4249 31263 4307 31269
rect 4249 31229 4261 31263
rect 4295 31260 4307 31263
rect 4890 31260 4896 31272
rect 4295 31232 4896 31260
rect 4295 31229 4307 31232
rect 4249 31223 4307 31229
rect 4890 31220 4896 31232
rect 4948 31220 4954 31272
rect 5994 31260 6000 31272
rect 5907 31232 6000 31260
rect 5994 31220 6000 31232
rect 6052 31220 6058 31272
rect 8389 31263 8447 31269
rect 8389 31229 8401 31263
rect 8435 31260 8447 31263
rect 10686 31260 10692 31272
rect 8435 31232 10692 31260
rect 8435 31229 8447 31232
rect 8389 31223 8447 31229
rect 10686 31220 10692 31232
rect 10744 31220 10750 31272
rect 12084 31260 12112 31291
rect 14016 31260 14044 31368
rect 16117 31365 16129 31368
rect 16163 31365 16175 31399
rect 16117 31359 16175 31365
rect 17129 31399 17187 31405
rect 17129 31365 17141 31399
rect 17175 31396 17187 31399
rect 17402 31396 17408 31408
rect 17175 31368 17408 31396
rect 17175 31365 17187 31368
rect 17129 31359 17187 31365
rect 15378 31328 15384 31340
rect 15291 31300 15384 31328
rect 15378 31288 15384 31300
rect 15436 31288 15442 31340
rect 16132 31328 16160 31359
rect 17402 31356 17408 31368
rect 17460 31356 17466 31408
rect 21177 31399 21235 31405
rect 21177 31396 21189 31399
rect 18354 31368 21189 31396
rect 21177 31365 21189 31368
rect 21223 31365 21235 31399
rect 21177 31359 21235 31365
rect 22922 31356 22928 31408
rect 22980 31396 22986 31408
rect 25685 31399 25743 31405
rect 22980 31368 24348 31396
rect 22980 31356 22986 31368
rect 16850 31328 16856 31340
rect 16132 31300 16856 31328
rect 16850 31288 16856 31300
rect 16908 31288 16914 31340
rect 20346 31288 20352 31340
rect 20404 31328 20410 31340
rect 20441 31331 20499 31337
rect 20441 31328 20453 31331
rect 20404 31300 20453 31328
rect 20404 31288 20410 31300
rect 20441 31297 20453 31300
rect 20487 31297 20499 31331
rect 20441 31291 20499 31297
rect 20806 31288 20812 31340
rect 20864 31328 20870 31340
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 20864 31300 21097 31328
rect 20864 31288 20870 31300
rect 21085 31297 21097 31300
rect 21131 31328 21143 31331
rect 21818 31328 21824 31340
rect 21131 31300 21824 31328
rect 21131 31297 21143 31300
rect 21085 31291 21143 31297
rect 21818 31288 21824 31300
rect 21876 31288 21882 31340
rect 22741 31331 22799 31337
rect 22741 31297 22753 31331
rect 22787 31328 22799 31331
rect 23474 31328 23480 31340
rect 22787 31300 23480 31328
rect 22787 31297 22799 31300
rect 22741 31291 22799 31297
rect 23474 31288 23480 31300
rect 23532 31288 23538 31340
rect 23658 31328 23664 31340
rect 23619 31300 23664 31328
rect 23658 31288 23664 31300
rect 23716 31288 23722 31340
rect 24320 31337 24348 31368
rect 25685 31365 25697 31399
rect 25731 31396 25743 31399
rect 26050 31396 26056 31408
rect 25731 31368 26056 31396
rect 25731 31365 25743 31368
rect 25685 31359 25743 31365
rect 26050 31356 26056 31368
rect 26108 31356 26114 31408
rect 27614 31356 27620 31408
rect 27672 31396 27678 31408
rect 30009 31399 30067 31405
rect 30009 31396 30021 31399
rect 27672 31368 30021 31396
rect 27672 31356 27678 31368
rect 30009 31365 30021 31368
rect 30055 31365 30067 31399
rect 30009 31359 30067 31365
rect 24305 31331 24363 31337
rect 24305 31297 24317 31331
rect 24351 31297 24363 31331
rect 24305 31291 24363 31297
rect 24946 31288 24952 31340
rect 25004 31328 25010 31340
rect 25133 31331 25191 31337
rect 25133 31328 25145 31331
rect 25004 31300 25145 31328
rect 25004 31288 25010 31300
rect 25133 31297 25145 31300
rect 25179 31297 25191 31331
rect 25133 31291 25191 31297
rect 25498 31288 25504 31340
rect 25556 31328 25562 31340
rect 25593 31331 25651 31337
rect 25593 31328 25605 31331
rect 25556 31300 25605 31328
rect 25556 31288 25562 31300
rect 25593 31297 25605 31300
rect 25639 31297 25651 31331
rect 26421 31331 26479 31337
rect 26421 31328 26433 31331
rect 25593 31291 25651 31297
rect 25700 31300 26433 31328
rect 12084 31232 14044 31260
rect 14093 31263 14151 31269
rect 14093 31229 14105 31263
rect 14139 31229 14151 31263
rect 14093 31223 14151 31229
rect 3421 31127 3479 31133
rect 3421 31093 3433 31127
rect 3467 31124 3479 31127
rect 3878 31124 3884 31136
rect 3467 31096 3884 31124
rect 3467 31093 3479 31096
rect 3421 31087 3479 31093
rect 3878 31084 3884 31096
rect 3936 31084 3942 31136
rect 6012 31124 6040 31220
rect 11238 31192 11244 31204
rect 9416 31164 11244 31192
rect 9416 31124 9444 31164
rect 11238 31152 11244 31164
rect 11296 31152 11302 31204
rect 13906 31152 13912 31204
rect 13964 31192 13970 31204
rect 14108 31192 14136 31223
rect 13964 31164 14136 31192
rect 13964 31152 13970 31164
rect 9858 31124 9864 31136
rect 6012 31096 9444 31124
rect 9819 31096 9864 31124
rect 9858 31084 9864 31096
rect 9916 31124 9922 31136
rect 10134 31124 10140 31136
rect 9916 31096 10140 31124
rect 9916 31084 9922 31096
rect 10134 31084 10140 31096
rect 10192 31084 10198 31136
rect 15396 31124 15424 31288
rect 16666 31220 16672 31272
rect 16724 31260 16730 31272
rect 20533 31263 20591 31269
rect 20533 31260 20545 31263
rect 16724 31232 20545 31260
rect 16724 31220 16730 31232
rect 20533 31229 20545 31232
rect 20579 31229 20591 31263
rect 20533 31223 20591 31229
rect 22186 31220 22192 31272
rect 22244 31260 22250 31272
rect 22557 31263 22615 31269
rect 22557 31260 22569 31263
rect 22244 31232 22569 31260
rect 22244 31220 22250 31232
rect 22557 31229 22569 31232
rect 22603 31260 22615 31263
rect 22646 31260 22652 31272
rect 22603 31232 22652 31260
rect 22603 31229 22615 31232
rect 22557 31223 22615 31229
rect 22646 31220 22652 31232
rect 22704 31220 22710 31272
rect 23566 31220 23572 31272
rect 23624 31260 23630 31272
rect 23842 31260 23848 31272
rect 23624 31232 23848 31260
rect 23624 31220 23630 31232
rect 23842 31220 23848 31232
rect 23900 31220 23906 31272
rect 22278 31192 22284 31204
rect 18432 31164 22284 31192
rect 17494 31124 17500 31136
rect 15396 31096 17500 31124
rect 17494 31084 17500 31096
rect 17552 31084 17558 31136
rect 17586 31084 17592 31136
rect 17644 31124 17650 31136
rect 18432 31124 18460 31164
rect 22278 31152 22284 31164
rect 22336 31152 22342 31204
rect 24397 31195 24455 31201
rect 24397 31161 24409 31195
rect 24443 31192 24455 31195
rect 25590 31192 25596 31204
rect 24443 31164 25596 31192
rect 24443 31161 24455 31164
rect 24397 31155 24455 31161
rect 25590 31152 25596 31164
rect 25648 31152 25654 31204
rect 18598 31124 18604 31136
rect 17644 31096 18460 31124
rect 18559 31096 18604 31124
rect 17644 31084 17650 31096
rect 18598 31084 18604 31096
rect 18656 31124 18662 31136
rect 23566 31124 23572 31136
rect 18656 31096 23572 31124
rect 18656 31084 18662 31096
rect 23566 31084 23572 31096
rect 23624 31084 23630 31136
rect 23753 31127 23811 31133
rect 23753 31093 23765 31127
rect 23799 31124 23811 31127
rect 24762 31124 24768 31136
rect 23799 31096 24768 31124
rect 23799 31093 23811 31096
rect 23753 31087 23811 31093
rect 24762 31084 24768 31096
rect 24820 31084 24826 31136
rect 24949 31127 25007 31133
rect 24949 31093 24961 31127
rect 24995 31124 25007 31127
rect 25700 31124 25728 31300
rect 26421 31297 26433 31300
rect 26467 31297 26479 31331
rect 27154 31328 27160 31340
rect 27115 31300 27160 31328
rect 26421 31291 26479 31297
rect 27154 31288 27160 31300
rect 27212 31288 27218 31340
rect 27985 31331 28043 31337
rect 27985 31297 27997 31331
rect 28031 31297 28043 31331
rect 29086 31328 29092 31340
rect 29047 31300 29092 31328
rect 27985 31291 28043 31297
rect 25774 31220 25780 31272
rect 25832 31260 25838 31272
rect 28000 31260 28028 31291
rect 29086 31288 29092 31300
rect 29144 31288 29150 31340
rect 29917 31331 29975 31337
rect 29917 31297 29929 31331
rect 29963 31328 29975 31331
rect 31754 31328 31760 31340
rect 29963 31300 31760 31328
rect 29963 31297 29975 31300
rect 29917 31291 29975 31297
rect 31754 31288 31760 31300
rect 31812 31328 31818 31340
rect 32582 31328 32588 31340
rect 31812 31300 32588 31328
rect 31812 31288 31818 31300
rect 32582 31288 32588 31300
rect 32640 31288 32646 31340
rect 28442 31260 28448 31272
rect 25832 31232 28028 31260
rect 28403 31232 28448 31260
rect 25832 31220 25838 31232
rect 28442 31220 28448 31232
rect 28500 31220 28506 31272
rect 26237 31195 26295 31201
rect 26237 31161 26249 31195
rect 26283 31192 26295 31195
rect 27798 31192 27804 31204
rect 26283 31164 27804 31192
rect 26283 31161 26295 31164
rect 26237 31155 26295 31161
rect 27798 31152 27804 31164
rect 27856 31152 27862 31204
rect 24995 31096 25728 31124
rect 24995 31093 25007 31096
rect 24949 31087 25007 31093
rect 26510 31084 26516 31136
rect 26568 31124 26574 31136
rect 26694 31124 26700 31136
rect 26568 31096 26700 31124
rect 26568 31084 26574 31096
rect 26694 31084 26700 31096
rect 26752 31084 26758 31136
rect 29178 31124 29184 31136
rect 29139 31096 29184 31124
rect 29178 31084 29184 31096
rect 29236 31084 29242 31136
rect 30098 31084 30104 31136
rect 30156 31124 30162 31136
rect 32674 31124 32680 31136
rect 30156 31096 32680 31124
rect 30156 31084 30162 31096
rect 32674 31084 32680 31096
rect 32732 31084 32738 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 16025 30923 16083 30929
rect 16025 30889 16037 30923
rect 16071 30920 16083 30923
rect 17586 30920 17592 30932
rect 16071 30892 17592 30920
rect 16071 30889 16083 30892
rect 16025 30883 16083 30889
rect 17586 30880 17592 30892
rect 17644 30880 17650 30932
rect 24946 30920 24952 30932
rect 17696 30892 24952 30920
rect 15746 30812 15752 30864
rect 15804 30852 15810 30864
rect 17696 30852 17724 30892
rect 24946 30880 24952 30892
rect 25004 30880 25010 30932
rect 25498 30880 25504 30932
rect 25556 30920 25562 30932
rect 25556 30892 26740 30920
rect 25556 30880 25562 30892
rect 15804 30824 17724 30852
rect 15804 30812 15810 30824
rect 17770 30812 17776 30864
rect 17828 30852 17834 30864
rect 24026 30852 24032 30864
rect 17828 30824 24032 30852
rect 17828 30812 17834 30824
rect 24026 30812 24032 30824
rect 24084 30812 24090 30864
rect 24964 30852 24992 30880
rect 24964 30824 26648 30852
rect 11146 30744 11152 30796
rect 11204 30784 11210 30796
rect 14277 30787 14335 30793
rect 14277 30784 14289 30787
rect 11204 30756 14289 30784
rect 11204 30744 11210 30756
rect 14277 30753 14289 30756
rect 14323 30753 14335 30787
rect 14277 30747 14335 30753
rect 14553 30787 14611 30793
rect 14553 30753 14565 30787
rect 14599 30784 14611 30787
rect 18414 30784 18420 30796
rect 14599 30756 18420 30784
rect 14599 30753 14611 30756
rect 14553 30747 14611 30753
rect 18414 30744 18420 30756
rect 18472 30744 18478 30796
rect 20162 30744 20168 30796
rect 20220 30784 20226 30796
rect 20438 30784 20444 30796
rect 20220 30756 20444 30784
rect 20220 30744 20226 30756
rect 20438 30744 20444 30756
rect 20496 30744 20502 30796
rect 25777 30787 25835 30793
rect 25777 30784 25789 30787
rect 21560 30756 22094 30784
rect 16206 30676 16212 30728
rect 16264 30716 16270 30728
rect 19242 30716 19248 30728
rect 16264 30688 19248 30716
rect 16264 30676 16270 30688
rect 19242 30676 19248 30688
rect 19300 30676 19306 30728
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30716 19763 30719
rect 19978 30716 19984 30728
rect 19751 30688 19984 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 19978 30676 19984 30688
rect 20036 30716 20042 30728
rect 20254 30716 20260 30728
rect 20036 30688 20260 30716
rect 20036 30676 20042 30688
rect 20254 30676 20260 30688
rect 20312 30676 20318 30728
rect 21450 30676 21456 30728
rect 21508 30716 21514 30728
rect 21560 30725 21588 30756
rect 21545 30719 21603 30725
rect 21545 30716 21557 30719
rect 21508 30688 21557 30716
rect 21508 30676 21514 30688
rect 21545 30685 21557 30688
rect 21591 30685 21603 30719
rect 22066 30716 22094 30756
rect 22940 30756 25789 30784
rect 22741 30719 22799 30725
rect 22741 30716 22753 30719
rect 21545 30679 21603 30685
rect 21652 30688 21956 30716
rect 22066 30688 22753 30716
rect 19334 30648 19340 30660
rect 15778 30620 19340 30648
rect 19334 30608 19340 30620
rect 19392 30608 19398 30660
rect 20530 30608 20536 30660
rect 20588 30648 20594 30660
rect 21082 30648 21088 30660
rect 20588 30620 20633 30648
rect 21043 30620 21088 30648
rect 20588 30608 20594 30620
rect 21082 30608 21088 30620
rect 21140 30648 21146 30660
rect 21652 30648 21680 30688
rect 21818 30648 21824 30660
rect 21140 30620 21680 30648
rect 21779 30620 21824 30648
rect 21140 30608 21146 30620
rect 21818 30608 21824 30620
rect 21876 30608 21882 30660
rect 21928 30648 21956 30688
rect 22741 30685 22753 30688
rect 22787 30685 22799 30719
rect 22741 30679 22799 30685
rect 22940 30648 22968 30756
rect 25777 30753 25789 30756
rect 25823 30753 25835 30787
rect 25777 30747 25835 30753
rect 23661 30719 23719 30725
rect 23661 30716 23673 30719
rect 23124 30688 23673 30716
rect 23124 30660 23152 30688
rect 23661 30685 23673 30688
rect 23707 30685 23719 30719
rect 23661 30679 23719 30685
rect 23750 30676 23756 30728
rect 23808 30716 23814 30728
rect 26620 30725 26648 30824
rect 24581 30719 24639 30725
rect 24581 30716 24593 30719
rect 23808 30688 24593 30716
rect 23808 30676 23814 30688
rect 24581 30685 24593 30688
rect 24627 30685 24639 30719
rect 24581 30679 24639 30685
rect 26605 30719 26663 30725
rect 26605 30685 26617 30719
rect 26651 30685 26663 30719
rect 26712 30716 26740 30892
rect 27154 30880 27160 30932
rect 27212 30920 27218 30932
rect 27212 30892 37780 30920
rect 27212 30880 27218 30892
rect 30098 30852 30104 30864
rect 28552 30824 30104 30852
rect 28552 30725 28580 30824
rect 30098 30812 30104 30824
rect 30156 30812 30162 30864
rect 30374 30852 30380 30864
rect 30335 30824 30380 30852
rect 30374 30812 30380 30824
rect 30432 30812 30438 30864
rect 34885 30855 34943 30861
rect 34885 30821 34897 30855
rect 34931 30852 34943 30855
rect 37366 30852 37372 30864
rect 34931 30824 37372 30852
rect 34931 30821 34943 30824
rect 34885 30815 34943 30821
rect 37366 30812 37372 30824
rect 37424 30812 37430 30864
rect 29178 30744 29184 30796
rect 29236 30784 29242 30796
rect 37752 30793 37780 30892
rect 37737 30787 37795 30793
rect 29236 30756 35112 30784
rect 29236 30744 29242 30756
rect 35084 30725 35112 30756
rect 37737 30753 37749 30787
rect 37783 30753 37795 30787
rect 37737 30747 37795 30753
rect 27249 30719 27307 30725
rect 27249 30716 27261 30719
rect 26712 30688 27261 30716
rect 26605 30679 26663 30685
rect 27249 30685 27261 30688
rect 27295 30685 27307 30719
rect 27249 30679 27307 30685
rect 27893 30719 27951 30725
rect 27893 30685 27905 30719
rect 27939 30685 27951 30719
rect 27893 30679 27951 30685
rect 28537 30719 28595 30725
rect 28537 30685 28549 30719
rect 28583 30685 28595 30719
rect 28537 30679 28595 30685
rect 35069 30719 35127 30725
rect 35069 30685 35081 30719
rect 35115 30685 35127 30719
rect 37458 30716 37464 30728
rect 37419 30688 37464 30716
rect 35069 30679 35127 30685
rect 21928 30620 22968 30648
rect 23017 30651 23075 30657
rect 23017 30617 23029 30651
rect 23063 30648 23075 30651
rect 23106 30648 23112 30660
rect 23063 30620 23112 30648
rect 23063 30617 23075 30620
rect 23017 30611 23075 30617
rect 23106 30608 23112 30620
rect 23164 30608 23170 30660
rect 25498 30648 25504 30660
rect 25459 30620 25504 30648
rect 25498 30608 25504 30620
rect 25556 30608 25562 30660
rect 25590 30608 25596 30660
rect 25648 30648 25654 30660
rect 27908 30648 27936 30679
rect 37458 30676 37464 30688
rect 37516 30676 37522 30728
rect 29822 30648 29828 30660
rect 25648 30620 25693 30648
rect 27908 30620 29684 30648
rect 29783 30620 29828 30648
rect 25648 30608 25654 30620
rect 9858 30540 9864 30592
rect 9916 30580 9922 30592
rect 17770 30580 17776 30592
rect 9916 30552 17776 30580
rect 9916 30540 9922 30552
rect 17770 30540 17776 30552
rect 17828 30540 17834 30592
rect 18230 30540 18236 30592
rect 18288 30580 18294 30592
rect 19797 30583 19855 30589
rect 19797 30580 19809 30583
rect 18288 30552 19809 30580
rect 18288 30540 18294 30552
rect 19797 30549 19809 30552
rect 19843 30549 19855 30583
rect 19797 30543 19855 30549
rect 20162 30540 20168 30592
rect 20220 30580 20226 30592
rect 23753 30583 23811 30589
rect 23753 30580 23765 30583
rect 20220 30552 23765 30580
rect 20220 30540 20226 30552
rect 23753 30549 23765 30552
rect 23799 30549 23811 30583
rect 23753 30543 23811 30549
rect 24673 30583 24731 30589
rect 24673 30549 24685 30583
rect 24719 30580 24731 30583
rect 25682 30580 25688 30592
rect 24719 30552 25688 30580
rect 24719 30549 24731 30552
rect 24673 30543 24731 30549
rect 25682 30540 25688 30552
rect 25740 30540 25746 30592
rect 26694 30580 26700 30592
rect 26655 30552 26700 30580
rect 26694 30540 26700 30552
rect 26752 30540 26758 30592
rect 27341 30583 27399 30589
rect 27341 30549 27353 30583
rect 27387 30580 27399 30583
rect 27706 30580 27712 30592
rect 27387 30552 27712 30580
rect 27387 30549 27399 30552
rect 27341 30543 27399 30549
rect 27706 30540 27712 30552
rect 27764 30540 27770 30592
rect 27890 30540 27896 30592
rect 27948 30580 27954 30592
rect 27985 30583 28043 30589
rect 27985 30580 27997 30583
rect 27948 30552 27997 30580
rect 27948 30540 27954 30552
rect 27985 30549 27997 30552
rect 28031 30549 28043 30583
rect 28626 30580 28632 30592
rect 28587 30552 28632 30580
rect 27985 30543 28043 30549
rect 28626 30540 28632 30552
rect 28684 30540 28690 30592
rect 29656 30580 29684 30620
rect 29822 30608 29828 30620
rect 29880 30608 29886 30660
rect 29914 30608 29920 30660
rect 29972 30648 29978 30660
rect 29972 30620 30017 30648
rect 29972 30608 29978 30620
rect 32030 30580 32036 30592
rect 29656 30552 32036 30580
rect 32030 30540 32036 30552
rect 32088 30540 32094 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 7098 30336 7104 30388
rect 7156 30376 7162 30388
rect 16206 30376 16212 30388
rect 7156 30348 16212 30376
rect 7156 30336 7162 30348
rect 16206 30336 16212 30348
rect 16264 30336 16270 30388
rect 16390 30336 16396 30388
rect 16448 30376 16454 30388
rect 18874 30376 18880 30388
rect 16448 30348 18880 30376
rect 16448 30336 16454 30348
rect 18874 30336 18880 30348
rect 18932 30336 18938 30388
rect 19797 30379 19855 30385
rect 19797 30345 19809 30379
rect 19843 30376 19855 30379
rect 20530 30376 20536 30388
rect 19843 30348 20536 30376
rect 19843 30345 19855 30348
rect 19797 30339 19855 30345
rect 20530 30336 20536 30348
rect 20588 30336 20594 30388
rect 22646 30336 22652 30388
rect 22704 30376 22710 30388
rect 27522 30376 27528 30388
rect 22704 30348 27528 30376
rect 22704 30336 22710 30348
rect 27522 30336 27528 30348
rect 27580 30336 27586 30388
rect 16666 30308 16672 30320
rect 13202 30280 16672 30308
rect 16666 30268 16672 30280
rect 16724 30268 16730 30320
rect 17221 30311 17279 30317
rect 17221 30277 17233 30311
rect 17267 30308 17279 30311
rect 17310 30308 17316 30320
rect 17267 30280 17316 30308
rect 17267 30277 17279 30280
rect 17221 30271 17279 30277
rect 17310 30268 17316 30280
rect 17368 30268 17374 30320
rect 20162 30308 20168 30320
rect 18446 30280 20168 30308
rect 20162 30268 20168 30280
rect 20220 30268 20226 30320
rect 22189 30311 22247 30317
rect 22189 30308 22201 30311
rect 20272 30280 22201 30308
rect 1854 30200 1860 30252
rect 1912 30240 1918 30252
rect 2038 30240 2044 30252
rect 1912 30212 2044 30240
rect 1912 30200 1918 30212
rect 2038 30200 2044 30212
rect 2096 30200 2102 30252
rect 13446 30200 13452 30252
rect 13504 30240 13510 30252
rect 16758 30240 16764 30252
rect 13504 30212 16764 30240
rect 13504 30200 13510 30212
rect 16758 30200 16764 30212
rect 16816 30200 16822 30252
rect 16850 30200 16856 30252
rect 16908 30240 16914 30252
rect 16945 30243 17003 30249
rect 16945 30240 16957 30243
rect 16908 30212 16957 30240
rect 16908 30200 16914 30212
rect 16945 30209 16957 30212
rect 16991 30209 17003 30243
rect 16945 30203 17003 30209
rect 19334 30200 19340 30252
rect 19392 30240 19398 30252
rect 19702 30240 19708 30252
rect 19392 30212 19708 30240
rect 19392 30200 19398 30212
rect 19702 30200 19708 30212
rect 19760 30200 19766 30252
rect 11606 30132 11612 30184
rect 11664 30172 11670 30184
rect 11701 30175 11759 30181
rect 11701 30172 11713 30175
rect 11664 30144 11713 30172
rect 11664 30132 11670 30144
rect 11701 30141 11713 30144
rect 11747 30141 11759 30175
rect 11701 30135 11759 30141
rect 11977 30175 12035 30181
rect 11977 30141 11989 30175
rect 12023 30172 12035 30175
rect 17954 30172 17960 30184
rect 12023 30144 17960 30172
rect 12023 30141 12035 30144
rect 11977 30135 12035 30141
rect 17954 30132 17960 30144
rect 18012 30132 18018 30184
rect 20272 30172 20300 30280
rect 22189 30277 22201 30280
rect 22235 30277 22247 30311
rect 22189 30271 22247 30277
rect 23658 30268 23664 30320
rect 23716 30308 23722 30320
rect 23753 30311 23811 30317
rect 23753 30308 23765 30311
rect 23716 30280 23765 30308
rect 23716 30268 23722 30280
rect 23753 30277 23765 30280
rect 23799 30277 23811 30311
rect 23753 30271 23811 30277
rect 24118 30268 24124 30320
rect 24176 30308 24182 30320
rect 24673 30311 24731 30317
rect 24673 30308 24685 30311
rect 24176 30280 24685 30308
rect 24176 30268 24182 30280
rect 24673 30277 24685 30280
rect 24719 30277 24731 30311
rect 26050 30308 26056 30320
rect 26011 30280 26056 30308
rect 24673 30271 24731 30277
rect 26050 30268 26056 30280
rect 26108 30268 26114 30320
rect 28813 30311 28871 30317
rect 28813 30277 28825 30311
rect 28859 30308 28871 30311
rect 29914 30308 29920 30320
rect 28859 30280 29920 30308
rect 28859 30277 28871 30280
rect 28813 30271 28871 30277
rect 29914 30268 29920 30280
rect 29972 30268 29978 30320
rect 20806 30240 20812 30252
rect 20767 30212 20812 30240
rect 20806 30200 20812 30212
rect 20864 30200 20870 30252
rect 25133 30243 25191 30249
rect 25133 30209 25145 30243
rect 25179 30209 25191 30243
rect 25133 30203 25191 30209
rect 25225 30243 25283 30249
rect 25225 30209 25237 30243
rect 25271 30240 25283 30243
rect 25590 30240 25596 30252
rect 25271 30212 25596 30240
rect 25271 30209 25283 30212
rect 25225 30203 25283 30209
rect 22097 30175 22155 30181
rect 22097 30172 22109 30175
rect 18248 30144 20300 30172
rect 20364 30144 22109 30172
rect 12986 30064 12992 30116
rect 13044 30104 13050 30116
rect 13446 30104 13452 30116
rect 13044 30076 13452 30104
rect 13044 30064 13050 30076
rect 13446 30064 13452 30076
rect 13504 30064 13510 30116
rect 15010 30064 15016 30116
rect 15068 30104 15074 30116
rect 16942 30104 16948 30116
rect 15068 30076 16948 30104
rect 15068 30064 15074 30076
rect 16942 30064 16948 30076
rect 17000 30064 17006 30116
rect 2133 30039 2191 30045
rect 2133 30005 2145 30039
rect 2179 30036 2191 30039
rect 4706 30036 4712 30048
rect 2179 30008 4712 30036
rect 2179 30005 2191 30008
rect 2133 29999 2191 30005
rect 4706 29996 4712 30008
rect 4764 29996 4770 30048
rect 13906 29996 13912 30048
rect 13964 30036 13970 30048
rect 18248 30036 18276 30144
rect 18322 30064 18328 30116
rect 18380 30104 18386 30116
rect 20364 30104 20392 30144
rect 22097 30141 22109 30144
rect 22143 30141 22155 30175
rect 22370 30172 22376 30184
rect 22331 30144 22376 30172
rect 22097 30135 22155 30141
rect 22370 30132 22376 30144
rect 22428 30132 22434 30184
rect 23661 30175 23719 30181
rect 23661 30141 23673 30175
rect 23707 30172 23719 30175
rect 25038 30172 25044 30184
rect 23707 30144 25044 30172
rect 23707 30141 23719 30144
rect 23661 30135 23719 30141
rect 25038 30132 25044 30144
rect 25096 30132 25102 30184
rect 18380 30076 20392 30104
rect 18380 30064 18386 30076
rect 20530 30064 20536 30116
rect 20588 30104 20594 30116
rect 25148 30104 25176 30203
rect 25590 30200 25596 30212
rect 25648 30200 25654 30252
rect 27617 30243 27675 30249
rect 27617 30209 27629 30243
rect 27663 30240 27675 30243
rect 28442 30240 28448 30252
rect 27663 30212 28448 30240
rect 27663 30209 27675 30212
rect 27617 30203 27675 30209
rect 28442 30200 28448 30212
rect 28500 30200 28506 30252
rect 28718 30240 28724 30252
rect 28679 30212 28724 30240
rect 28718 30200 28724 30212
rect 28776 30200 28782 30252
rect 29365 30243 29423 30249
rect 29365 30209 29377 30243
rect 29411 30240 29423 30243
rect 34514 30240 34520 30252
rect 29411 30212 34520 30240
rect 29411 30209 29423 30212
rect 29365 30203 29423 30209
rect 34514 30200 34520 30212
rect 34572 30200 34578 30252
rect 25498 30132 25504 30184
rect 25556 30172 25562 30184
rect 25961 30175 26019 30181
rect 25961 30172 25973 30175
rect 25556 30144 25973 30172
rect 25556 30132 25562 30144
rect 25961 30141 25973 30144
rect 26007 30172 26019 30175
rect 27798 30172 27804 30184
rect 26007 30144 27016 30172
rect 27759 30144 27804 30172
rect 26007 30141 26019 30144
rect 25961 30135 26019 30141
rect 20588 30076 25176 30104
rect 26513 30107 26571 30113
rect 20588 30064 20594 30076
rect 26513 30073 26525 30107
rect 26559 30073 26571 30107
rect 26988 30104 27016 30144
rect 27798 30132 27804 30144
rect 27856 30132 27862 30184
rect 29457 30107 29515 30113
rect 29457 30104 29469 30107
rect 26988 30076 29469 30104
rect 26513 30067 26571 30073
rect 29457 30073 29469 30076
rect 29503 30073 29515 30107
rect 29457 30067 29515 30073
rect 18690 30036 18696 30048
rect 13964 30008 18276 30036
rect 18651 30008 18696 30036
rect 13964 29996 13970 30008
rect 18690 29996 18696 30008
rect 18748 29996 18754 30048
rect 19058 29996 19064 30048
rect 19116 30036 19122 30048
rect 20901 30039 20959 30045
rect 20901 30036 20913 30039
rect 19116 30008 20913 30036
rect 19116 29996 19122 30008
rect 20901 30005 20913 30008
rect 20947 30005 20959 30039
rect 20901 29999 20959 30005
rect 22094 29996 22100 30048
rect 22152 30036 22158 30048
rect 22370 30036 22376 30048
rect 22152 30008 22376 30036
rect 22152 29996 22158 30008
rect 22370 29996 22376 30008
rect 22428 29996 22434 30048
rect 24026 29996 24032 30048
rect 24084 30036 24090 30048
rect 26528 30036 26556 30067
rect 27982 30036 27988 30048
rect 24084 30008 26556 30036
rect 27943 30008 27988 30036
rect 24084 29996 24090 30008
rect 27982 29996 27988 30008
rect 28040 30036 28046 30048
rect 29086 30036 29092 30048
rect 28040 30008 29092 30036
rect 28040 29996 28046 30008
rect 29086 29996 29092 30008
rect 29144 29996 29150 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 2746 29804 17724 29832
rect 2314 29724 2320 29776
rect 2372 29764 2378 29776
rect 2746 29764 2774 29804
rect 2372 29736 2774 29764
rect 13357 29767 13415 29773
rect 2372 29724 2378 29736
rect 13357 29733 13369 29767
rect 13403 29764 13415 29767
rect 13998 29764 14004 29776
rect 13403 29736 14004 29764
rect 13403 29733 13415 29736
rect 13357 29727 13415 29733
rect 13998 29724 14004 29736
rect 14056 29724 14062 29776
rect 17696 29764 17724 29804
rect 17770 29792 17776 29844
rect 17828 29832 17834 29844
rect 18141 29835 18199 29841
rect 18141 29832 18153 29835
rect 17828 29804 18153 29832
rect 17828 29792 17834 29804
rect 18141 29801 18153 29804
rect 18187 29832 18199 29835
rect 18414 29832 18420 29844
rect 18187 29804 18420 29832
rect 18187 29801 18199 29804
rect 18141 29795 18199 29801
rect 18414 29792 18420 29804
rect 18472 29792 18478 29844
rect 18874 29792 18880 29844
rect 18932 29832 18938 29844
rect 21542 29832 21548 29844
rect 18932 29804 21548 29832
rect 18932 29792 18938 29804
rect 21542 29792 21548 29804
rect 21600 29792 21606 29844
rect 26605 29767 26663 29773
rect 26605 29764 26617 29767
rect 17696 29736 18460 29764
rect 16393 29699 16451 29705
rect 16393 29665 16405 29699
rect 16439 29696 16451 29699
rect 16758 29696 16764 29708
rect 16439 29668 16764 29696
rect 16439 29665 16451 29668
rect 16393 29659 16451 29665
rect 16758 29656 16764 29668
rect 16816 29656 16822 29708
rect 17034 29656 17040 29708
rect 17092 29696 17098 29708
rect 18432 29696 18460 29736
rect 18892 29736 26617 29764
rect 18892 29696 18920 29736
rect 26605 29733 26617 29736
rect 26651 29733 26663 29767
rect 26605 29727 26663 29733
rect 21634 29696 21640 29708
rect 17092 29668 18368 29696
rect 18432 29668 18920 29696
rect 21595 29668 21640 29696
rect 17092 29656 17098 29668
rect 1762 29628 1768 29640
rect 1723 29600 1768 29628
rect 1762 29588 1768 29600
rect 1820 29588 1826 29640
rect 11606 29628 11612 29640
rect 11567 29600 11612 29628
rect 11606 29588 11612 29600
rect 11664 29588 11670 29640
rect 18230 29628 18236 29640
rect 17802 29600 18236 29628
rect 18230 29588 18236 29600
rect 18288 29588 18294 29640
rect 18340 29628 18368 29668
rect 21634 29656 21640 29668
rect 21692 29656 21698 29708
rect 27617 29699 27675 29705
rect 27617 29665 27629 29699
rect 27663 29696 27675 29699
rect 28626 29696 28632 29708
rect 27663 29668 28632 29696
rect 27663 29665 27675 29668
rect 27617 29659 27675 29665
rect 28626 29656 28632 29668
rect 28684 29656 28690 29708
rect 18693 29631 18751 29637
rect 18693 29628 18705 29631
rect 18340 29600 18705 29628
rect 18693 29597 18705 29600
rect 18739 29597 18751 29631
rect 18693 29591 18751 29597
rect 18782 29588 18788 29640
rect 18840 29628 18846 29640
rect 19521 29631 19579 29637
rect 18840 29600 18885 29628
rect 18840 29588 18846 29600
rect 19521 29597 19533 29631
rect 19567 29628 19579 29631
rect 20162 29628 20168 29640
rect 19567 29600 20168 29628
rect 19567 29597 19579 29600
rect 19521 29591 19579 29597
rect 20162 29588 20168 29600
rect 20220 29588 20226 29640
rect 20257 29631 20315 29637
rect 20257 29597 20269 29631
rect 20303 29628 20315 29631
rect 20346 29628 20352 29640
rect 20303 29600 20352 29628
rect 20303 29597 20315 29600
rect 20257 29591 20315 29597
rect 20346 29588 20352 29600
rect 20404 29628 20410 29640
rect 20898 29628 20904 29640
rect 20404 29600 20904 29628
rect 20404 29588 20410 29600
rect 20898 29588 20904 29600
rect 20956 29588 20962 29640
rect 23106 29628 23112 29640
rect 21284 29600 21496 29628
rect 23067 29600 23112 29628
rect 11790 29520 11796 29572
rect 11848 29560 11854 29572
rect 11885 29563 11943 29569
rect 11885 29560 11897 29563
rect 11848 29532 11897 29560
rect 11848 29520 11854 29532
rect 11885 29529 11897 29532
rect 11931 29529 11943 29563
rect 13722 29560 13728 29572
rect 13110 29532 13728 29560
rect 11885 29523 11943 29529
rect 13722 29520 13728 29532
rect 13780 29520 13786 29572
rect 16666 29560 16672 29572
rect 16627 29532 16672 29560
rect 16666 29520 16672 29532
rect 16724 29520 16730 29572
rect 17972 29532 18276 29560
rect 1581 29495 1639 29501
rect 1581 29461 1593 29495
rect 1627 29492 1639 29495
rect 1946 29492 1952 29504
rect 1627 29464 1952 29492
rect 1627 29461 1639 29464
rect 1581 29455 1639 29461
rect 1946 29452 1952 29464
rect 2004 29452 2010 29504
rect 14182 29452 14188 29504
rect 14240 29492 14246 29504
rect 17972 29492 18000 29532
rect 14240 29464 18000 29492
rect 18248 29492 18276 29532
rect 18414 29520 18420 29572
rect 18472 29560 18478 29572
rect 19426 29560 19432 29572
rect 18472 29532 19432 29560
rect 18472 29520 18478 29532
rect 19426 29520 19432 29532
rect 19484 29520 19490 29572
rect 19613 29563 19671 29569
rect 19613 29529 19625 29563
rect 19659 29560 19671 29563
rect 21284 29560 21312 29600
rect 19659 29532 21312 29560
rect 21468 29560 21496 29600
rect 23106 29588 23112 29600
rect 23164 29588 23170 29640
rect 23750 29628 23756 29640
rect 23711 29600 23756 29628
rect 23750 29588 23756 29600
rect 23808 29588 23814 29640
rect 26421 29631 26479 29637
rect 26421 29597 26433 29631
rect 26467 29628 26479 29631
rect 27154 29628 27160 29640
rect 26467 29600 27160 29628
rect 26467 29597 26479 29600
rect 26421 29591 26479 29597
rect 27154 29588 27160 29600
rect 27212 29588 27218 29640
rect 36630 29588 36636 29640
rect 36688 29628 36694 29640
rect 38013 29631 38071 29637
rect 38013 29628 38025 29631
rect 36688 29600 38025 29628
rect 36688 29588 36694 29600
rect 38013 29597 38025 29600
rect 38059 29597 38071 29631
rect 38013 29591 38071 29597
rect 21729 29563 21787 29569
rect 21729 29560 21741 29563
rect 21468 29532 21741 29560
rect 19659 29529 19671 29532
rect 19613 29523 19671 29529
rect 21729 29529 21741 29532
rect 21775 29529 21787 29563
rect 22649 29563 22707 29569
rect 22649 29560 22661 29563
rect 21729 29523 21787 29529
rect 22388 29532 22661 29560
rect 22388 29504 22416 29532
rect 22649 29529 22661 29532
rect 22695 29560 22707 29563
rect 23382 29560 23388 29572
rect 22695 29532 23388 29560
rect 22695 29529 22707 29532
rect 22649 29523 22707 29529
rect 23382 29520 23388 29532
rect 23440 29520 23446 29572
rect 24673 29563 24731 29569
rect 24673 29529 24685 29563
rect 24719 29529 24731 29563
rect 24673 29523 24731 29529
rect 20349 29495 20407 29501
rect 20349 29492 20361 29495
rect 18248 29464 20361 29492
rect 14240 29452 14246 29464
rect 20349 29461 20361 29464
rect 20395 29461 20407 29495
rect 20349 29455 20407 29461
rect 20622 29452 20628 29504
rect 20680 29492 20686 29504
rect 20993 29495 21051 29501
rect 20993 29492 21005 29495
rect 20680 29464 21005 29492
rect 20680 29452 20686 29464
rect 20993 29461 21005 29464
rect 21039 29461 21051 29495
rect 20993 29455 21051 29461
rect 22370 29452 22376 29504
rect 22428 29452 22434 29504
rect 22554 29452 22560 29504
rect 22612 29492 22618 29504
rect 23201 29495 23259 29501
rect 23201 29492 23213 29495
rect 22612 29464 23213 29492
rect 22612 29452 22618 29464
rect 23201 29461 23213 29464
rect 23247 29461 23259 29495
rect 23201 29455 23259 29461
rect 23750 29452 23756 29504
rect 23808 29492 23814 29504
rect 23845 29495 23903 29501
rect 23845 29492 23857 29495
rect 23808 29464 23857 29492
rect 23808 29452 23814 29464
rect 23845 29461 23857 29464
rect 23891 29461 23903 29495
rect 23845 29455 23903 29461
rect 23934 29452 23940 29504
rect 23992 29492 23998 29504
rect 24688 29492 24716 29523
rect 24762 29520 24768 29572
rect 24820 29560 24826 29572
rect 24820 29532 24865 29560
rect 24820 29520 24826 29532
rect 24946 29520 24952 29572
rect 25004 29560 25010 29572
rect 25222 29560 25228 29572
rect 25004 29532 25228 29560
rect 25004 29520 25010 29532
rect 25222 29520 25228 29532
rect 25280 29560 25286 29572
rect 25685 29563 25743 29569
rect 25685 29560 25697 29563
rect 25280 29532 25697 29560
rect 25280 29520 25286 29532
rect 25685 29529 25697 29532
rect 25731 29529 25743 29563
rect 25685 29523 25743 29529
rect 27706 29520 27712 29572
rect 27764 29560 27770 29572
rect 28629 29563 28687 29569
rect 27764 29532 27809 29560
rect 27764 29520 27770 29532
rect 28629 29529 28641 29563
rect 28675 29529 28687 29563
rect 28629 29523 28687 29529
rect 27338 29492 27344 29504
rect 23992 29464 27344 29492
rect 23992 29452 23998 29464
rect 27338 29452 27344 29464
rect 27396 29452 27402 29504
rect 27798 29452 27804 29504
rect 27856 29492 27862 29504
rect 28644 29492 28672 29523
rect 38194 29492 38200 29504
rect 27856 29464 28672 29492
rect 38155 29464 38200 29492
rect 27856 29452 27862 29464
rect 38194 29452 38200 29464
rect 38252 29452 38258 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 4062 29248 4068 29300
rect 4120 29288 4126 29300
rect 8297 29291 8355 29297
rect 8297 29288 8309 29291
rect 4120 29260 8309 29288
rect 4120 29248 4126 29260
rect 8297 29257 8309 29260
rect 8343 29257 8355 29291
rect 8297 29251 8355 29257
rect 8941 29291 8999 29297
rect 8941 29257 8953 29291
rect 8987 29288 8999 29291
rect 13906 29288 13912 29300
rect 8987 29260 13912 29288
rect 8987 29257 8999 29260
rect 8941 29251 8999 29257
rect 5626 29180 5632 29232
rect 5684 29220 5690 29232
rect 5684 29192 7314 29220
rect 5684 29180 5690 29192
rect 1762 29152 1768 29164
rect 1723 29124 1768 29152
rect 1762 29112 1768 29124
rect 1820 29112 1826 29164
rect 3237 29155 3295 29161
rect 3237 29121 3249 29155
rect 3283 29152 3295 29155
rect 3786 29152 3792 29164
rect 3283 29124 3792 29152
rect 3283 29121 3295 29124
rect 3237 29115 3295 29121
rect 3786 29112 3792 29124
rect 3844 29112 3850 29164
rect 8312 29152 8340 29251
rect 13906 29248 13912 29260
rect 13964 29248 13970 29300
rect 16758 29288 16764 29300
rect 14292 29260 16764 29288
rect 10229 29223 10287 29229
rect 10229 29189 10241 29223
rect 10275 29220 10287 29223
rect 11054 29220 11060 29232
rect 10275 29192 11060 29220
rect 10275 29189 10287 29192
rect 10229 29183 10287 29189
rect 11054 29180 11060 29192
rect 11112 29180 11118 29232
rect 14182 29220 14188 29232
rect 13202 29192 14188 29220
rect 14182 29180 14188 29192
rect 14240 29180 14246 29232
rect 14292 29161 14320 29260
rect 16758 29248 16764 29260
rect 16816 29248 16822 29300
rect 19058 29288 19064 29300
rect 17052 29260 19064 29288
rect 17052 29220 17080 29260
rect 19058 29248 19064 29260
rect 19116 29248 19122 29300
rect 19150 29248 19156 29300
rect 19208 29288 19214 29300
rect 19208 29260 20760 29288
rect 19208 29248 19214 29260
rect 15778 29192 17080 29220
rect 17129 29223 17187 29229
rect 17129 29189 17141 29223
rect 17175 29220 17187 29223
rect 17218 29220 17224 29232
rect 17175 29192 17224 29220
rect 17175 29189 17187 29192
rect 17129 29183 17187 29189
rect 17218 29180 17224 29192
rect 17276 29180 17282 29232
rect 20622 29220 20628 29232
rect 18354 29192 20628 29220
rect 20622 29180 20628 29192
rect 20680 29180 20686 29232
rect 20732 29229 20760 29260
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 22278 29288 22284 29300
rect 20956 29260 22284 29288
rect 20956 29248 20962 29260
rect 22278 29248 22284 29260
rect 22336 29288 22342 29300
rect 23106 29288 23112 29300
rect 22336 29260 23112 29288
rect 22336 29248 22342 29260
rect 23106 29248 23112 29260
rect 23164 29248 23170 29300
rect 23934 29288 23940 29300
rect 23584 29260 23940 29288
rect 23584 29229 23612 29260
rect 23934 29248 23940 29260
rect 23992 29248 23998 29300
rect 27801 29291 27859 29297
rect 27801 29257 27813 29291
rect 27847 29288 27859 29291
rect 27982 29288 27988 29300
rect 27847 29260 27988 29288
rect 27847 29257 27859 29260
rect 27801 29251 27859 29257
rect 27982 29248 27988 29260
rect 28040 29248 28046 29300
rect 20717 29223 20775 29229
rect 20717 29189 20729 29223
rect 20763 29189 20775 29223
rect 20717 29183 20775 29189
rect 23569 29223 23627 29229
rect 23569 29189 23581 29223
rect 23615 29189 23627 29223
rect 23569 29183 23627 29189
rect 23661 29223 23719 29229
rect 23661 29189 23673 29223
rect 23707 29220 23719 29223
rect 24670 29220 24676 29232
rect 23707 29192 24676 29220
rect 23707 29189 23719 29192
rect 23661 29183 23719 29189
rect 24670 29180 24676 29192
rect 24728 29180 24734 29232
rect 25314 29180 25320 29232
rect 25372 29220 25378 29232
rect 25777 29223 25835 29229
rect 25777 29220 25789 29223
rect 25372 29192 25789 29220
rect 25372 29180 25378 29192
rect 25777 29189 25789 29192
rect 25823 29189 25835 29223
rect 25777 29183 25835 29189
rect 26329 29223 26387 29229
rect 26329 29189 26341 29223
rect 26375 29220 26387 29223
rect 26418 29220 26424 29232
rect 26375 29192 26424 29220
rect 26375 29189 26387 29192
rect 26329 29183 26387 29189
rect 26418 29180 26424 29192
rect 26476 29220 26482 29232
rect 26476 29192 30604 29220
rect 26476 29180 26482 29192
rect 8849 29155 8907 29161
rect 8849 29152 8861 29155
rect 8312 29124 8861 29152
rect 8849 29121 8861 29124
rect 8895 29121 8907 29155
rect 8849 29115 8907 29121
rect 9493 29155 9551 29161
rect 9493 29121 9505 29155
rect 9539 29121 9551 29155
rect 9493 29115 9551 29121
rect 14277 29155 14335 29161
rect 14277 29121 14289 29155
rect 14323 29121 14335 29155
rect 14277 29115 14335 29121
rect 1854 29044 1860 29096
rect 1912 29084 1918 29096
rect 4798 29084 4804 29096
rect 1912 29056 4804 29084
rect 1912 29044 1918 29056
rect 4798 29044 4804 29056
rect 4856 29044 4862 29096
rect 6546 29084 6552 29096
rect 6507 29056 6552 29084
rect 6546 29044 6552 29056
rect 6604 29044 6610 29096
rect 9508 29084 9536 29115
rect 21634 29112 21640 29164
rect 21692 29152 21698 29164
rect 22005 29155 22063 29161
rect 22005 29152 22017 29155
rect 21692 29124 22017 29152
rect 21692 29112 21698 29124
rect 22005 29121 22017 29124
rect 22051 29121 22063 29155
rect 22005 29115 22063 29121
rect 22281 29155 22339 29161
rect 22281 29121 22293 29155
rect 22327 29152 22339 29155
rect 22462 29152 22468 29164
rect 22327 29124 22468 29152
rect 22327 29121 22339 29124
rect 22281 29115 22339 29121
rect 22462 29112 22468 29124
rect 22520 29112 22526 29164
rect 26694 29112 26700 29164
rect 26752 29152 26758 29164
rect 27341 29155 27399 29161
rect 27341 29152 27353 29155
rect 26752 29124 27353 29152
rect 26752 29112 26758 29124
rect 27341 29121 27353 29124
rect 27387 29121 27399 29155
rect 27341 29115 27399 29121
rect 27982 29112 27988 29164
rect 28040 29152 28046 29164
rect 30576 29161 30604 29192
rect 28261 29155 28319 29161
rect 28261 29152 28273 29155
rect 28040 29124 28273 29152
rect 28040 29112 28046 29124
rect 28261 29121 28273 29124
rect 28307 29121 28319 29155
rect 28261 29115 28319 29121
rect 30561 29155 30619 29161
rect 30561 29121 30573 29155
rect 30607 29121 30619 29155
rect 30561 29115 30619 29121
rect 6656 29056 9536 29084
rect 11057 29087 11115 29093
rect 3142 28976 3148 29028
rect 3200 29016 3206 29028
rect 3329 29019 3387 29025
rect 3329 29016 3341 29019
rect 3200 28988 3341 29016
rect 3200 28976 3206 28988
rect 3329 28985 3341 28988
rect 3375 28985 3387 29019
rect 4816 29016 4844 29044
rect 6656 29016 6684 29056
rect 11057 29053 11069 29087
rect 11103 29084 11115 29087
rect 11238 29084 11244 29096
rect 11103 29056 11244 29084
rect 11103 29053 11115 29056
rect 11057 29047 11115 29053
rect 11238 29044 11244 29056
rect 11296 29084 11302 29096
rect 11606 29084 11612 29096
rect 11296 29056 11612 29084
rect 11296 29044 11302 29056
rect 11606 29044 11612 29056
rect 11664 29084 11670 29096
rect 11701 29087 11759 29093
rect 11701 29084 11713 29087
rect 11664 29056 11713 29084
rect 11664 29044 11670 29056
rect 11701 29053 11713 29056
rect 11747 29053 11759 29087
rect 11701 29047 11759 29053
rect 13725 29087 13783 29093
rect 13725 29053 13737 29087
rect 13771 29084 13783 29087
rect 16114 29084 16120 29096
rect 13771 29056 16120 29084
rect 13771 29053 13783 29056
rect 13725 29047 13783 29053
rect 16114 29044 16120 29056
rect 16172 29044 16178 29096
rect 16850 29084 16856 29096
rect 16811 29056 16856 29084
rect 16850 29044 16856 29056
rect 16908 29044 16914 29096
rect 17862 29084 17868 29096
rect 16960 29056 17868 29084
rect 4816 28988 6684 29016
rect 9585 29019 9643 29025
rect 3329 28979 3387 28985
rect 9585 28985 9597 29019
rect 9631 29016 9643 29019
rect 11146 29016 11152 29028
rect 9631 28988 11152 29016
rect 9631 28985 9643 28988
rect 9585 28979 9643 28985
rect 11146 28976 11152 28988
rect 11204 28976 11210 29028
rect 16025 29019 16083 29025
rect 16025 28985 16037 29019
rect 16071 29016 16083 29019
rect 16666 29016 16672 29028
rect 16071 28988 16672 29016
rect 16071 28985 16083 28988
rect 16025 28979 16083 28985
rect 16666 28976 16672 28988
rect 16724 29016 16730 29028
rect 16960 29016 16988 29056
rect 17862 29044 17868 29056
rect 17920 29044 17926 29096
rect 18138 29044 18144 29096
rect 18196 29084 18202 29096
rect 18601 29087 18659 29093
rect 18601 29084 18613 29087
rect 18196 29056 18613 29084
rect 18196 29044 18202 29056
rect 18601 29053 18613 29056
rect 18647 29053 18659 29087
rect 18601 29047 18659 29053
rect 20438 29044 20444 29096
rect 20496 29084 20502 29096
rect 20625 29087 20683 29093
rect 20625 29084 20637 29087
rect 20496 29056 20637 29084
rect 20496 29044 20502 29056
rect 20625 29053 20637 29056
rect 20671 29053 20683 29087
rect 20625 29047 20683 29053
rect 23382 29044 23388 29096
rect 23440 29084 23446 29096
rect 23845 29087 23903 29093
rect 23845 29084 23857 29087
rect 23440 29056 23857 29084
rect 23440 29044 23446 29056
rect 23845 29053 23857 29056
rect 23891 29053 23903 29087
rect 23845 29047 23903 29053
rect 25685 29087 25743 29093
rect 25685 29053 25697 29087
rect 25731 29084 25743 29087
rect 26050 29084 26056 29096
rect 25731 29056 26056 29084
rect 25731 29053 25743 29056
rect 25685 29047 25743 29053
rect 26050 29044 26056 29056
rect 26108 29044 26114 29096
rect 27157 29087 27215 29093
rect 27157 29053 27169 29087
rect 27203 29084 27215 29087
rect 28445 29087 28503 29093
rect 27203 29056 28212 29084
rect 27203 29053 27215 29056
rect 27157 29047 27215 29053
rect 16724 28988 16988 29016
rect 21177 29019 21235 29025
rect 16724 28976 16730 28988
rect 21177 28985 21189 29019
rect 21223 29016 21235 29019
rect 24026 29016 24032 29028
rect 21223 28988 24032 29016
rect 21223 28985 21235 28988
rect 21177 28979 21235 28985
rect 24026 28976 24032 28988
rect 24084 28976 24090 29028
rect 28184 28960 28212 29056
rect 28445 29053 28457 29087
rect 28491 29084 28503 29087
rect 28994 29084 29000 29096
rect 28491 29056 29000 29084
rect 28491 29053 28503 29056
rect 28445 29047 28503 29053
rect 28994 29044 29000 29056
rect 29052 29044 29058 29096
rect 1578 28948 1584 28960
rect 1539 28920 1584 28948
rect 1578 28908 1584 28920
rect 1636 28908 1642 28960
rect 6812 28951 6870 28957
rect 6812 28917 6824 28951
rect 6858 28948 6870 28951
rect 9674 28948 9680 28960
rect 6858 28920 9680 28948
rect 6858 28917 6870 28920
rect 6812 28911 6870 28917
rect 9674 28908 9680 28920
rect 9732 28908 9738 28960
rect 11964 28951 12022 28957
rect 11964 28917 11976 28951
rect 12010 28948 12022 28951
rect 14366 28948 14372 28960
rect 12010 28920 14372 28948
rect 12010 28917 12022 28920
rect 11964 28911 12022 28917
rect 14366 28908 14372 28920
rect 14424 28908 14430 28960
rect 14540 28951 14598 28957
rect 14540 28917 14552 28951
rect 14586 28948 14598 28951
rect 15930 28948 15936 28960
rect 14586 28920 15936 28948
rect 14586 28917 14598 28920
rect 14540 28911 14598 28917
rect 15930 28908 15936 28920
rect 15988 28908 15994 28960
rect 16114 28908 16120 28960
rect 16172 28948 16178 28960
rect 27798 28948 27804 28960
rect 16172 28920 27804 28948
rect 16172 28908 16178 28920
rect 27798 28908 27804 28920
rect 27856 28908 27862 28960
rect 28166 28908 28172 28960
rect 28224 28948 28230 28960
rect 28629 28951 28687 28957
rect 28629 28948 28641 28951
rect 28224 28920 28641 28948
rect 28224 28908 28230 28920
rect 28629 28917 28641 28920
rect 28675 28917 28687 28951
rect 28629 28911 28687 28917
rect 30653 28951 30711 28957
rect 30653 28917 30665 28951
rect 30699 28948 30711 28951
rect 31478 28948 31484 28960
rect 30699 28920 31484 28948
rect 30699 28917 30711 28920
rect 30653 28911 30711 28917
rect 31478 28908 31484 28920
rect 31536 28908 31542 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 9674 28704 9680 28756
rect 9732 28744 9738 28756
rect 13998 28744 14004 28756
rect 9732 28716 14004 28744
rect 9732 28704 9738 28716
rect 13998 28704 14004 28716
rect 14056 28704 14062 28756
rect 14090 28704 14096 28756
rect 14148 28744 14154 28756
rect 14277 28747 14335 28753
rect 14277 28744 14289 28747
rect 14148 28716 14289 28744
rect 14148 28704 14154 28716
rect 14277 28713 14289 28716
rect 14323 28713 14335 28747
rect 14277 28707 14335 28713
rect 15930 28704 15936 28756
rect 15988 28744 15994 28756
rect 18598 28744 18604 28756
rect 15988 28716 18604 28744
rect 15988 28704 15994 28716
rect 18598 28704 18604 28716
rect 18656 28704 18662 28756
rect 22094 28704 22100 28756
rect 22152 28744 22158 28756
rect 23198 28744 23204 28756
rect 22152 28716 23204 28744
rect 22152 28704 22158 28716
rect 23198 28704 23204 28716
rect 23256 28704 23262 28756
rect 28166 28744 28172 28756
rect 28127 28716 28172 28744
rect 28166 28704 28172 28716
rect 28224 28704 28230 28756
rect 12526 28636 12532 28688
rect 12584 28676 12590 28688
rect 14550 28676 14556 28688
rect 12584 28648 14556 28676
rect 12584 28636 12590 28648
rect 14550 28636 14556 28648
rect 14608 28636 14614 28688
rect 17218 28636 17224 28688
rect 17276 28676 17282 28688
rect 19334 28676 19340 28688
rect 17276 28648 19340 28676
rect 17276 28636 17282 28648
rect 19334 28636 19340 28648
rect 19392 28636 19398 28688
rect 19426 28636 19432 28688
rect 19484 28676 19490 28688
rect 26418 28676 26424 28688
rect 19484 28648 24624 28676
rect 26379 28648 26424 28676
rect 19484 28636 19490 28648
rect 5994 28608 6000 28620
rect 2792 28580 6000 28608
rect 1854 28540 1860 28552
rect 1815 28512 1860 28540
rect 1854 28500 1860 28512
rect 1912 28500 1918 28552
rect 2792 28549 2820 28580
rect 5994 28568 6000 28580
rect 6052 28568 6058 28620
rect 21637 28611 21695 28617
rect 21637 28608 21649 28611
rect 12636 28580 21649 28608
rect 2777 28543 2835 28549
rect 2777 28509 2789 28543
rect 2823 28509 2835 28543
rect 2777 28503 2835 28509
rect 3970 28500 3976 28552
rect 4028 28540 4034 28552
rect 6546 28540 6552 28552
rect 4028 28512 6552 28540
rect 4028 28500 4034 28512
rect 6546 28500 6552 28512
rect 6604 28540 6610 28552
rect 6917 28543 6975 28549
rect 6917 28540 6929 28543
rect 6604 28512 6929 28540
rect 6604 28500 6610 28512
rect 6917 28509 6929 28512
rect 6963 28509 6975 28543
rect 11238 28540 11244 28552
rect 11199 28512 11244 28540
rect 6917 28503 6975 28509
rect 11238 28500 11244 28512
rect 11296 28500 11302 28552
rect 12636 28526 12664 28580
rect 21637 28577 21649 28580
rect 21683 28577 21695 28611
rect 21637 28571 21695 28577
rect 23017 28611 23075 28617
rect 23017 28577 23029 28611
rect 23063 28608 23075 28611
rect 23063 28580 24532 28608
rect 23063 28577 23075 28580
rect 23017 28571 23075 28577
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28540 13599 28543
rect 13814 28540 13820 28552
rect 13587 28512 13820 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 13814 28500 13820 28512
rect 13872 28500 13878 28552
rect 14458 28540 14464 28552
rect 14419 28512 14464 28540
rect 14458 28500 14464 28512
rect 14516 28500 14522 28552
rect 15194 28549 15200 28552
rect 15186 28543 15200 28549
rect 15186 28540 15198 28543
rect 15155 28512 15198 28540
rect 15186 28509 15198 28512
rect 15186 28503 15200 28509
rect 15194 28500 15200 28503
rect 15252 28500 15258 28552
rect 16574 28500 16580 28552
rect 16632 28500 16638 28552
rect 16850 28500 16856 28552
rect 16908 28540 16914 28552
rect 18233 28543 18291 28549
rect 18233 28540 18245 28543
rect 16908 28512 18245 28540
rect 16908 28500 16914 28512
rect 18233 28509 18245 28512
rect 18279 28509 18291 28543
rect 18233 28503 18291 28509
rect 19981 28543 20039 28549
rect 19981 28509 19993 28543
rect 20027 28540 20039 28543
rect 20070 28540 20076 28552
rect 20027 28512 20076 28540
rect 20027 28509 20039 28512
rect 19981 28503 20039 28509
rect 20070 28500 20076 28512
rect 20128 28540 20134 28552
rect 20346 28540 20352 28552
rect 20128 28512 20352 28540
rect 20128 28500 20134 28512
rect 20346 28500 20352 28512
rect 20404 28500 20410 28552
rect 20622 28540 20628 28552
rect 20583 28512 20628 28540
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 21545 28543 21603 28549
rect 20732 28512 21036 28540
rect 1949 28475 2007 28481
rect 1949 28441 1961 28475
rect 1995 28472 2007 28475
rect 3326 28472 3332 28484
rect 1995 28444 3332 28472
rect 1995 28441 2007 28444
rect 1949 28435 2007 28441
rect 3326 28432 3332 28444
rect 3384 28432 3390 28484
rect 5626 28432 5632 28484
rect 5684 28472 5690 28484
rect 6181 28475 6239 28481
rect 6181 28472 6193 28475
rect 5684 28444 6193 28472
rect 5684 28432 5690 28444
rect 6181 28441 6193 28444
rect 6227 28441 6239 28475
rect 6181 28435 6239 28441
rect 11517 28475 11575 28481
rect 11517 28441 11529 28475
rect 11563 28472 11575 28475
rect 11606 28472 11612 28484
rect 11563 28444 11612 28472
rect 11563 28441 11575 28444
rect 11517 28435 11575 28441
rect 11606 28432 11612 28444
rect 11664 28432 11670 28484
rect 15473 28475 15531 28481
rect 15473 28441 15485 28475
rect 15519 28472 15531 28475
rect 15746 28472 15752 28484
rect 15519 28444 15752 28472
rect 15519 28441 15531 28444
rect 15473 28435 15531 28441
rect 15746 28432 15752 28444
rect 15804 28432 15810 28484
rect 16758 28432 16764 28484
rect 16816 28472 16822 28484
rect 17494 28472 17500 28484
rect 16816 28444 17080 28472
rect 17455 28444 17500 28472
rect 16816 28432 16822 28444
rect 2866 28404 2872 28416
rect 2827 28376 2872 28404
rect 2866 28364 2872 28376
rect 2924 28364 2930 28416
rect 5994 28364 6000 28416
rect 6052 28404 6058 28416
rect 12526 28404 12532 28416
rect 6052 28376 12532 28404
rect 6052 28364 6058 28376
rect 12526 28364 12532 28376
rect 12584 28364 12590 28416
rect 12986 28404 12992 28416
rect 12947 28376 12992 28404
rect 12986 28364 12992 28376
rect 13044 28364 13050 28416
rect 13630 28404 13636 28416
rect 13591 28376 13636 28404
rect 13630 28364 13636 28376
rect 13688 28364 13694 28416
rect 13998 28364 14004 28416
rect 14056 28404 14062 28416
rect 16942 28404 16948 28416
rect 14056 28376 16948 28404
rect 14056 28364 14062 28376
rect 16942 28364 16948 28376
rect 17000 28364 17006 28416
rect 17052 28404 17080 28444
rect 17494 28432 17500 28444
rect 17552 28432 17558 28484
rect 20732 28472 20760 28512
rect 20898 28472 20904 28484
rect 17604 28444 20760 28472
rect 20859 28444 20904 28472
rect 17604 28404 17632 28444
rect 20898 28432 20904 28444
rect 20956 28432 20962 28484
rect 21008 28472 21036 28512
rect 21545 28509 21557 28543
rect 21591 28540 21603 28543
rect 21818 28540 21824 28552
rect 21591 28512 21824 28540
rect 21591 28509 21603 28512
rect 21545 28503 21603 28509
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 22189 28543 22247 28549
rect 22189 28509 22201 28543
rect 22235 28540 22247 28543
rect 22278 28540 22284 28552
rect 22235 28512 22284 28540
rect 22235 28509 22247 28512
rect 22189 28503 22247 28509
rect 22278 28500 22284 28512
rect 22336 28500 22342 28552
rect 22002 28472 22008 28484
rect 21008 28444 22008 28472
rect 22002 28432 22008 28444
rect 22060 28432 22066 28484
rect 23109 28475 23167 28481
rect 23109 28441 23121 28475
rect 23155 28472 23167 28475
rect 23934 28472 23940 28484
rect 23155 28444 23940 28472
rect 23155 28441 23167 28444
rect 23109 28435 23167 28441
rect 23934 28432 23940 28444
rect 23992 28432 23998 28484
rect 24029 28475 24087 28481
rect 24029 28441 24041 28475
rect 24075 28472 24087 28475
rect 24118 28472 24124 28484
rect 24075 28444 24124 28472
rect 24075 28441 24087 28444
rect 24029 28435 24087 28441
rect 24118 28432 24124 28444
rect 24176 28432 24182 28484
rect 24504 28472 24532 28580
rect 24596 28549 24624 28648
rect 26418 28636 26424 28648
rect 26476 28636 26482 28688
rect 27798 28636 27804 28688
rect 27856 28676 27862 28688
rect 28350 28676 28356 28688
rect 27856 28648 28356 28676
rect 27856 28636 27862 28648
rect 28350 28636 28356 28648
rect 28408 28636 28414 28688
rect 25869 28611 25927 28617
rect 25869 28577 25881 28611
rect 25915 28608 25927 28611
rect 27614 28608 27620 28620
rect 25915 28580 27620 28608
rect 25915 28577 25927 28580
rect 25869 28571 25927 28577
rect 27614 28568 27620 28580
rect 27672 28568 27678 28620
rect 27709 28611 27767 28617
rect 27709 28577 27721 28611
rect 27755 28608 27767 28611
rect 28721 28611 28779 28617
rect 28721 28608 28733 28611
rect 27755 28580 28733 28608
rect 27755 28577 27767 28580
rect 27709 28571 27767 28577
rect 28721 28577 28733 28580
rect 28767 28577 28779 28611
rect 37274 28608 37280 28620
rect 28721 28571 28779 28577
rect 29748 28580 37280 28608
rect 24581 28543 24639 28549
rect 24581 28509 24593 28543
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 27525 28543 27583 28549
rect 27525 28509 27537 28543
rect 27571 28509 27583 28543
rect 27525 28503 27583 28509
rect 24504 28444 25544 28472
rect 17052 28376 17632 28404
rect 17862 28364 17868 28416
rect 17920 28404 17926 28416
rect 19426 28404 19432 28416
rect 17920 28376 19432 28404
rect 17920 28364 17926 28376
rect 19426 28364 19432 28376
rect 19484 28364 19490 28416
rect 20070 28404 20076 28416
rect 20031 28376 20076 28404
rect 20070 28364 20076 28376
rect 20128 28364 20134 28416
rect 20162 28364 20168 28416
rect 20220 28404 20226 28416
rect 22281 28407 22339 28413
rect 22281 28404 22293 28407
rect 20220 28376 22293 28404
rect 20220 28364 20226 28376
rect 22281 28373 22293 28376
rect 22327 28373 22339 28407
rect 22281 28367 22339 28373
rect 24486 28364 24492 28416
rect 24544 28404 24550 28416
rect 24673 28407 24731 28413
rect 24673 28404 24685 28407
rect 24544 28376 24685 28404
rect 24544 28364 24550 28376
rect 24673 28373 24685 28376
rect 24719 28373 24731 28407
rect 25516 28404 25544 28444
rect 25590 28432 25596 28484
rect 25648 28472 25654 28484
rect 25961 28475 26019 28481
rect 25961 28472 25973 28475
rect 25648 28444 25973 28472
rect 25648 28432 25654 28444
rect 25961 28441 25973 28444
rect 26007 28441 26019 28475
rect 25961 28435 26019 28441
rect 27246 28432 27252 28484
rect 27304 28472 27310 28484
rect 27540 28472 27568 28503
rect 28534 28500 28540 28552
rect 28592 28540 28598 28552
rect 28629 28543 28687 28549
rect 28629 28540 28641 28543
rect 28592 28512 28641 28540
rect 28592 28500 28598 28512
rect 28629 28509 28641 28512
rect 28675 28509 28687 28543
rect 28629 28503 28687 28509
rect 29638 28500 29644 28552
rect 29696 28540 29702 28552
rect 29748 28549 29776 28580
rect 37274 28568 37280 28580
rect 37332 28568 37338 28620
rect 29733 28543 29791 28549
rect 29733 28540 29745 28543
rect 29696 28512 29745 28540
rect 29696 28500 29702 28512
rect 29733 28509 29745 28512
rect 29779 28509 29791 28543
rect 31478 28540 31484 28552
rect 31439 28512 31484 28540
rect 29733 28503 29791 28509
rect 31478 28500 31484 28512
rect 31536 28500 31542 28552
rect 29825 28475 29883 28481
rect 29825 28472 29837 28475
rect 27304 28444 29837 28472
rect 27304 28432 27310 28444
rect 29825 28441 29837 28444
rect 29871 28441 29883 28475
rect 29825 28435 29883 28441
rect 27890 28404 27896 28416
rect 25516 28376 27896 28404
rect 24673 28367 24731 28373
rect 27890 28364 27896 28376
rect 27948 28364 27954 28416
rect 31297 28407 31355 28413
rect 31297 28373 31309 28407
rect 31343 28404 31355 28407
rect 33042 28404 33048 28416
rect 31343 28376 33048 28404
rect 31343 28373 31355 28376
rect 31297 28367 31355 28373
rect 33042 28364 33048 28376
rect 33100 28364 33106 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 22554 28200 22560 28212
rect 12406 28172 22560 28200
rect 5994 28132 6000 28144
rect 5955 28104 6000 28132
rect 5994 28092 6000 28104
rect 6052 28092 6058 28144
rect 12406 28132 12434 28172
rect 22554 28160 22560 28172
rect 22612 28160 22618 28212
rect 26418 28200 26424 28212
rect 24320 28172 26424 28200
rect 9706 28104 12434 28132
rect 13630 28092 13636 28144
rect 13688 28092 13694 28144
rect 15010 28092 15016 28144
rect 15068 28132 15074 28144
rect 17218 28132 17224 28144
rect 15068 28104 17224 28132
rect 15068 28092 15074 28104
rect 17218 28092 17224 28104
rect 17276 28092 17282 28144
rect 20070 28132 20076 28144
rect 18354 28104 20076 28132
rect 20070 28092 20076 28104
rect 20128 28092 20134 28144
rect 20993 28135 21051 28141
rect 20993 28101 21005 28135
rect 21039 28132 21051 28135
rect 22189 28135 22247 28141
rect 22189 28132 22201 28135
rect 21039 28104 22201 28132
rect 21039 28101 21051 28104
rect 20993 28095 21051 28101
rect 22189 28101 22201 28104
rect 22235 28101 22247 28135
rect 22189 28095 22247 28101
rect 22278 28092 22284 28144
rect 22336 28132 22342 28144
rect 23750 28132 23756 28144
rect 22336 28104 23336 28132
rect 23711 28104 23756 28132
rect 22336 28092 22342 28104
rect 1762 28064 1768 28076
rect 1723 28036 1768 28064
rect 1762 28024 1768 28036
rect 1820 28024 1826 28076
rect 5382 28036 5488 28064
rect 5460 28008 5488 28036
rect 6546 28024 6552 28076
rect 6604 28064 6610 28076
rect 8205 28067 8263 28073
rect 8205 28064 8217 28067
rect 6604 28036 8217 28064
rect 6604 28024 6610 28036
rect 8205 28033 8217 28036
rect 8251 28033 8263 28067
rect 12802 28064 12808 28076
rect 12763 28036 12808 28064
rect 8205 28027 8263 28033
rect 12802 28024 12808 28036
rect 12860 28024 12866 28076
rect 14550 28024 14556 28076
rect 14608 28064 14614 28076
rect 16758 28064 16764 28076
rect 14608 28036 16764 28064
rect 14608 28024 14614 28036
rect 16758 28024 16764 28036
rect 16816 28024 16822 28076
rect 19058 28064 19064 28076
rect 19019 28036 19064 28064
rect 19058 28024 19064 28036
rect 19116 28024 19122 28076
rect 19150 28024 19156 28076
rect 19208 28064 19214 28076
rect 19208 28036 19253 28064
rect 19208 28024 19214 28036
rect 20806 28024 20812 28076
rect 20864 28064 20870 28076
rect 20901 28067 20959 28073
rect 20901 28064 20913 28067
rect 20864 28036 20913 28064
rect 20864 28024 20870 28036
rect 20901 28033 20913 28036
rect 20947 28033 20959 28067
rect 20901 28027 20959 28033
rect 3970 27996 3976 28008
rect 3931 27968 3976 27996
rect 3970 27956 3976 27968
rect 4028 27956 4034 28008
rect 4249 27999 4307 28005
rect 4249 27965 4261 27999
rect 4295 27996 4307 27999
rect 4982 27996 4988 28008
rect 4295 27968 4988 27996
rect 4295 27965 4307 27968
rect 4249 27959 4307 27965
rect 4982 27956 4988 27968
rect 5040 27956 5046 28008
rect 5442 27956 5448 28008
rect 5500 27956 5506 28008
rect 8481 27999 8539 28005
rect 8481 27965 8493 27999
rect 8527 27996 8539 27999
rect 13081 27999 13139 28005
rect 8527 27968 12434 27996
rect 8527 27965 8539 27968
rect 8481 27959 8539 27965
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 2222 27860 2228 27872
rect 1627 27832 2228 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 2222 27820 2228 27832
rect 2280 27820 2286 27872
rect 9950 27860 9956 27872
rect 9911 27832 9956 27860
rect 9950 27820 9956 27832
rect 10008 27820 10014 27872
rect 12406 27860 12434 27968
rect 13081 27965 13093 27999
rect 13127 27996 13139 27999
rect 13127 27968 15148 27996
rect 13127 27965 13139 27968
rect 13081 27959 13139 27965
rect 15120 27928 15148 27968
rect 15194 27956 15200 28008
rect 15252 27996 15258 28008
rect 16850 27996 16856 28008
rect 15252 27968 16856 27996
rect 15252 27956 15258 27968
rect 16850 27956 16856 27968
rect 16908 27956 16914 28008
rect 17129 27999 17187 28005
rect 17129 27965 17141 27999
rect 17175 27996 17187 27999
rect 17678 27996 17684 28008
rect 17175 27968 17684 27996
rect 17175 27965 17187 27968
rect 17129 27959 17187 27965
rect 17678 27956 17684 27968
rect 17736 27956 17742 28008
rect 17862 27956 17868 28008
rect 17920 27996 17926 28008
rect 20824 27996 20852 28024
rect 17920 27968 20852 27996
rect 22097 27999 22155 28005
rect 17920 27956 17926 27968
rect 22097 27965 22109 27999
rect 22143 27965 22155 27999
rect 22097 27959 22155 27965
rect 23109 27999 23167 28005
rect 23109 27965 23121 27999
rect 23155 27996 23167 27999
rect 23198 27996 23204 28008
rect 23155 27968 23204 27996
rect 23155 27965 23167 27968
rect 23109 27959 23167 27965
rect 16298 27928 16304 27940
rect 14108 27900 14688 27928
rect 15120 27900 16304 27928
rect 14108 27860 14136 27900
rect 14550 27860 14556 27872
rect 12406 27832 14136 27860
rect 14511 27832 14556 27860
rect 14550 27820 14556 27832
rect 14608 27820 14614 27872
rect 14660 27860 14688 27900
rect 16298 27888 16304 27900
rect 16356 27888 16362 27940
rect 18230 27888 18236 27940
rect 18288 27928 18294 27940
rect 21910 27928 21916 27940
rect 18288 27900 21916 27928
rect 18288 27888 18294 27900
rect 21910 27888 21916 27900
rect 21968 27888 21974 27940
rect 22112 27928 22140 27959
rect 23198 27956 23204 27968
rect 23256 27956 23262 28008
rect 23308 27996 23336 28104
rect 23750 28092 23756 28104
rect 23808 28092 23814 28144
rect 24320 28141 24348 28172
rect 26418 28160 26424 28172
rect 26476 28160 26482 28212
rect 28994 28200 29000 28212
rect 28955 28172 29000 28200
rect 28994 28160 29000 28172
rect 29052 28160 29058 28212
rect 24305 28135 24363 28141
rect 24305 28101 24317 28135
rect 24351 28101 24363 28135
rect 25682 28132 25688 28144
rect 25643 28104 25688 28132
rect 24305 28095 24363 28101
rect 25682 28092 25688 28104
rect 25740 28092 25746 28144
rect 26510 28092 26516 28144
rect 26568 28132 26574 28144
rect 26605 28135 26663 28141
rect 26605 28132 26617 28135
rect 26568 28104 26617 28132
rect 26568 28092 26574 28104
rect 26605 28101 26617 28104
rect 26651 28101 26663 28135
rect 27338 28132 27344 28144
rect 27299 28104 27344 28132
rect 26605 28095 26663 28101
rect 27338 28092 27344 28104
rect 27396 28092 27402 28144
rect 27893 28135 27951 28141
rect 27893 28101 27905 28135
rect 27939 28132 27951 28135
rect 28258 28132 28264 28144
rect 27939 28104 28264 28132
rect 27939 28101 27951 28104
rect 27893 28095 27951 28101
rect 28258 28092 28264 28104
rect 28316 28092 28322 28144
rect 29270 28132 29276 28144
rect 28368 28104 29276 28132
rect 24765 28067 24823 28073
rect 24765 28033 24777 28067
rect 24811 28064 24823 28067
rect 25038 28064 25044 28076
rect 24811 28036 25044 28064
rect 24811 28033 24823 28036
rect 24765 28027 24823 28033
rect 23661 27999 23719 28005
rect 23308 27968 23612 27996
rect 23290 27928 23296 27940
rect 22112 27900 23296 27928
rect 23290 27888 23296 27900
rect 23348 27888 23354 27940
rect 23584 27928 23612 27968
rect 23661 27965 23673 27999
rect 23707 27996 23719 27999
rect 24026 27996 24032 28008
rect 23707 27968 24032 27996
rect 23707 27965 23719 27968
rect 23661 27959 23719 27965
rect 24026 27956 24032 27968
rect 24084 27956 24090 28008
rect 24780 27928 24808 28027
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 28368 28073 28396 28104
rect 29270 28092 29276 28104
rect 29328 28092 29334 28144
rect 28353 28067 28411 28073
rect 28353 28033 28365 28067
rect 28399 28033 28411 28067
rect 29178 28064 29184 28076
rect 29139 28036 29184 28064
rect 28353 28027 28411 28033
rect 29178 28024 29184 28036
rect 29236 28024 29242 28076
rect 38010 28064 38016 28076
rect 37971 28036 38016 28064
rect 38010 28024 38016 28036
rect 38068 28024 38074 28076
rect 25590 27996 25596 28008
rect 25551 27968 25596 27996
rect 25590 27956 25596 27968
rect 25648 27956 25654 28008
rect 27246 27996 27252 28008
rect 27207 27968 27252 27996
rect 27246 27956 27252 27968
rect 27304 27956 27310 28008
rect 23584 27900 24808 27928
rect 24854 27888 24860 27940
rect 24912 27928 24918 27940
rect 38194 27928 38200 27940
rect 24912 27900 24957 27928
rect 38155 27900 38200 27928
rect 24912 27888 24918 27900
rect 38194 27888 38200 27900
rect 38252 27888 38258 27940
rect 17862 27860 17868 27872
rect 14660 27832 17868 27860
rect 17862 27820 17868 27832
rect 17920 27820 17926 27872
rect 18138 27820 18144 27872
rect 18196 27860 18202 27872
rect 18601 27863 18659 27869
rect 18601 27860 18613 27863
rect 18196 27832 18613 27860
rect 18196 27820 18202 27832
rect 18601 27829 18613 27832
rect 18647 27829 18659 27863
rect 18601 27823 18659 27829
rect 19426 27820 19432 27872
rect 19484 27860 19490 27872
rect 25222 27860 25228 27872
rect 19484 27832 25228 27860
rect 19484 27820 19490 27832
rect 25222 27820 25228 27832
rect 25280 27820 25286 27872
rect 28074 27820 28080 27872
rect 28132 27860 28138 27872
rect 28442 27860 28448 27872
rect 28132 27832 28448 27860
rect 28132 27820 28138 27832
rect 28442 27820 28448 27832
rect 28500 27820 28506 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1578 27616 1584 27668
rect 1636 27656 1642 27668
rect 1838 27659 1896 27665
rect 1838 27656 1850 27659
rect 1636 27628 1850 27656
rect 1636 27616 1642 27628
rect 1838 27625 1850 27628
rect 1884 27625 1896 27659
rect 1838 27619 1896 27625
rect 12986 27616 12992 27668
rect 13044 27656 13050 27668
rect 17954 27656 17960 27668
rect 13044 27628 17960 27656
rect 13044 27616 13050 27628
rect 17954 27616 17960 27628
rect 18012 27616 18018 27668
rect 18046 27616 18052 27668
rect 18104 27656 18110 27668
rect 18690 27656 18696 27668
rect 18104 27628 18696 27656
rect 18104 27616 18110 27628
rect 18690 27616 18696 27628
rect 18748 27616 18754 27668
rect 18782 27616 18788 27668
rect 18840 27656 18846 27668
rect 20254 27656 20260 27668
rect 18840 27628 20260 27656
rect 18840 27616 18846 27628
rect 20254 27616 20260 27628
rect 20312 27616 20318 27668
rect 21542 27616 21548 27668
rect 21600 27656 21606 27668
rect 27157 27659 27215 27665
rect 27157 27656 27169 27659
rect 21600 27628 27169 27656
rect 21600 27616 21606 27628
rect 27157 27625 27169 27628
rect 27203 27625 27215 27659
rect 27157 27619 27215 27625
rect 3329 27591 3387 27597
rect 3329 27557 3341 27591
rect 3375 27588 3387 27591
rect 4890 27588 4896 27600
rect 3375 27560 4896 27588
rect 3375 27557 3387 27560
rect 3329 27551 3387 27557
rect 4890 27548 4896 27560
rect 4948 27548 4954 27600
rect 17126 27548 17132 27600
rect 17184 27588 17190 27600
rect 19242 27588 19248 27600
rect 17184 27560 19248 27588
rect 17184 27548 17190 27560
rect 19242 27548 19248 27560
rect 19300 27548 19306 27600
rect 21818 27548 21824 27600
rect 21876 27548 21882 27600
rect 24670 27588 24676 27600
rect 24631 27560 24676 27588
rect 24670 27548 24676 27560
rect 24728 27548 24734 27600
rect 24762 27548 24768 27600
rect 24820 27588 24826 27600
rect 25961 27591 26019 27597
rect 24820 27560 25912 27588
rect 24820 27548 24826 27560
rect 1581 27523 1639 27529
rect 1581 27489 1593 27523
rect 1627 27520 1639 27523
rect 3970 27520 3976 27532
rect 1627 27492 3976 27520
rect 1627 27489 1639 27492
rect 1581 27483 1639 27489
rect 3970 27480 3976 27492
rect 4028 27480 4034 27532
rect 12802 27480 12808 27532
rect 12860 27520 12866 27532
rect 15194 27520 15200 27532
rect 12860 27492 15200 27520
rect 12860 27480 12866 27492
rect 15194 27480 15200 27492
rect 15252 27520 15258 27532
rect 15841 27523 15899 27529
rect 15841 27520 15853 27523
rect 15252 27492 15853 27520
rect 15252 27480 15258 27492
rect 15841 27489 15853 27492
rect 15887 27489 15899 27523
rect 15841 27483 15899 27489
rect 16104 27523 16162 27529
rect 16104 27489 16116 27523
rect 16150 27520 16162 27523
rect 16206 27520 16212 27532
rect 16150 27492 16212 27520
rect 16150 27489 16162 27492
rect 16104 27483 16162 27489
rect 16206 27480 16212 27492
rect 16264 27480 16270 27532
rect 16482 27480 16488 27532
rect 16540 27520 16546 27532
rect 21358 27520 21364 27532
rect 16540 27492 21364 27520
rect 16540 27480 16546 27492
rect 21358 27480 21364 27492
rect 21416 27480 21422 27532
rect 21836 27520 21864 27548
rect 21913 27523 21971 27529
rect 21913 27520 21925 27523
rect 21836 27492 21925 27520
rect 21913 27489 21925 27492
rect 21959 27489 21971 27523
rect 21913 27483 21971 27489
rect 4433 27455 4491 27461
rect 4433 27421 4445 27455
rect 4479 27452 4491 27455
rect 4798 27452 4804 27464
rect 4479 27424 4804 27452
rect 4479 27421 4491 27424
rect 4433 27415 4491 27421
rect 4798 27412 4804 27424
rect 4856 27452 4862 27464
rect 5258 27452 5264 27464
rect 4856 27424 5264 27452
rect 4856 27412 4862 27424
rect 5258 27412 5264 27424
rect 5316 27412 5322 27464
rect 18230 27452 18236 27464
rect 17250 27424 18236 27452
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27452 18383 27455
rect 18598 27452 18604 27464
rect 18371 27424 18604 27452
rect 18371 27421 18383 27424
rect 18325 27415 18383 27421
rect 18598 27412 18604 27424
rect 18656 27412 18662 27464
rect 19426 27412 19432 27464
rect 19484 27452 19490 27464
rect 19521 27455 19579 27461
rect 19521 27452 19533 27455
rect 19484 27424 19533 27452
rect 19484 27412 19490 27424
rect 19521 27421 19533 27424
rect 19567 27421 19579 27455
rect 23382 27452 23388 27464
rect 23343 27424 23388 27452
rect 19521 27415 19579 27421
rect 23382 27412 23388 27424
rect 23440 27412 23446 27464
rect 24578 27452 24584 27464
rect 24539 27424 24584 27452
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 24854 27412 24860 27464
rect 24912 27452 24918 27464
rect 25225 27455 25283 27461
rect 25225 27452 25237 27455
rect 24912 27424 25237 27452
rect 24912 27412 24918 27424
rect 25225 27421 25237 27424
rect 25271 27421 25283 27455
rect 25225 27415 25283 27421
rect 25314 27412 25320 27464
rect 25372 27452 25378 27464
rect 25884 27461 25912 27560
rect 25961 27557 25973 27591
rect 26007 27588 26019 27591
rect 27338 27588 27344 27600
rect 26007 27560 27344 27588
rect 26007 27557 26019 27560
rect 25961 27551 26019 27557
rect 27338 27548 27344 27560
rect 27396 27548 27402 27600
rect 28445 27591 28503 27597
rect 28445 27557 28457 27591
rect 28491 27588 28503 27591
rect 29178 27588 29184 27600
rect 28491 27560 29184 27588
rect 28491 27557 28503 27560
rect 28445 27551 28503 27557
rect 29178 27548 29184 27560
rect 29236 27548 29242 27600
rect 32401 27591 32459 27597
rect 32401 27557 32413 27591
rect 32447 27588 32459 27591
rect 36630 27588 36636 27600
rect 32447 27560 36636 27588
rect 32447 27557 32459 27560
rect 32401 27551 32459 27557
rect 36630 27548 36636 27560
rect 36688 27548 36694 27600
rect 28350 27520 28356 27532
rect 27816 27492 28356 27520
rect 25869 27455 25927 27461
rect 25372 27424 25417 27452
rect 25372 27412 25378 27424
rect 25869 27421 25881 27455
rect 25915 27421 25927 27455
rect 25869 27415 25927 27421
rect 26513 27455 26571 27461
rect 26513 27421 26525 27455
rect 26559 27452 26571 27455
rect 27341 27455 27399 27461
rect 26559 27424 27292 27452
rect 26559 27421 26571 27424
rect 26513 27415 26571 27421
rect 3142 27384 3148 27396
rect 3082 27356 3148 27384
rect 3142 27344 3148 27356
rect 3200 27344 3206 27396
rect 3510 27344 3516 27396
rect 3568 27384 3574 27396
rect 10229 27387 10287 27393
rect 10229 27384 10241 27387
rect 3568 27356 10241 27384
rect 3568 27344 3574 27356
rect 10229 27353 10241 27356
rect 10275 27353 10287 27387
rect 10229 27347 10287 27353
rect 10502 27344 10508 27396
rect 10560 27384 10566 27396
rect 16390 27384 16396 27396
rect 10560 27356 16396 27384
rect 10560 27344 10566 27356
rect 16390 27344 16396 27356
rect 16448 27344 16454 27396
rect 17402 27344 17408 27396
rect 17460 27384 17466 27396
rect 17865 27387 17923 27393
rect 17865 27384 17877 27387
rect 17460 27356 17877 27384
rect 17460 27344 17466 27356
rect 17865 27353 17877 27356
rect 17911 27353 17923 27387
rect 17865 27347 17923 27353
rect 18417 27387 18475 27393
rect 18417 27353 18429 27387
rect 18463 27384 18475 27387
rect 19705 27387 19763 27393
rect 19705 27384 19717 27387
rect 18463 27356 19717 27384
rect 18463 27353 18475 27356
rect 18417 27347 18475 27353
rect 19705 27353 19717 27356
rect 19751 27353 19763 27387
rect 21358 27384 21364 27396
rect 21319 27356 21364 27384
rect 19705 27347 19763 27353
rect 21358 27344 21364 27356
rect 21416 27344 21422 27396
rect 22002 27344 22008 27396
rect 22060 27384 22066 27396
rect 22922 27384 22928 27396
rect 22060 27356 22105 27384
rect 22883 27356 22928 27384
rect 22060 27344 22066 27356
rect 22922 27344 22928 27356
rect 22980 27344 22986 27396
rect 27264 27384 27292 27424
rect 27341 27421 27353 27455
rect 27387 27452 27399 27455
rect 27430 27452 27436 27464
rect 27387 27424 27436 27452
rect 27387 27421 27399 27424
rect 27341 27415 27399 27421
rect 27430 27412 27436 27424
rect 27488 27412 27494 27464
rect 27816 27461 27844 27492
rect 28350 27480 28356 27492
rect 28408 27480 28414 27532
rect 27801 27455 27859 27461
rect 27801 27421 27813 27455
rect 27847 27421 27859 27455
rect 27801 27415 27859 27421
rect 28534 27412 28540 27464
rect 28592 27452 28598 27464
rect 28629 27455 28687 27461
rect 28629 27452 28641 27455
rect 28592 27424 28641 27452
rect 28592 27412 28598 27424
rect 28629 27421 28641 27424
rect 28675 27421 28687 27455
rect 28629 27415 28687 27421
rect 29733 27455 29791 27461
rect 29733 27421 29745 27455
rect 29779 27421 29791 27455
rect 30374 27452 30380 27464
rect 30335 27424 30380 27452
rect 29733 27415 29791 27421
rect 28350 27384 28356 27396
rect 27264 27356 28356 27384
rect 28350 27344 28356 27356
rect 28408 27344 28414 27396
rect 29748 27384 29776 27415
rect 30374 27412 30380 27424
rect 30432 27412 30438 27464
rect 31570 27412 31576 27464
rect 31628 27452 31634 27464
rect 32585 27455 32643 27461
rect 32585 27452 32597 27455
rect 31628 27424 32597 27452
rect 31628 27412 31634 27424
rect 32585 27421 32597 27424
rect 32631 27421 32643 27455
rect 32585 27415 32643 27421
rect 33042 27412 33048 27464
rect 33100 27452 33106 27464
rect 38013 27455 38071 27461
rect 38013 27452 38025 27455
rect 33100 27424 38025 27452
rect 33100 27412 33106 27424
rect 38013 27421 38025 27424
rect 38059 27421 38071 27455
rect 38013 27415 38071 27421
rect 37458 27384 37464 27396
rect 29748 27356 37464 27384
rect 37458 27344 37464 27356
rect 37516 27384 37522 27396
rect 37918 27384 37924 27396
rect 37516 27356 37924 27384
rect 37516 27344 37522 27356
rect 37918 27344 37924 27356
rect 37976 27344 37982 27396
rect 4525 27319 4583 27325
rect 4525 27285 4537 27319
rect 4571 27316 4583 27319
rect 7006 27316 7012 27328
rect 4571 27288 7012 27316
rect 4571 27285 4583 27288
rect 4525 27279 4583 27285
rect 7006 27276 7012 27288
rect 7064 27276 7070 27328
rect 11514 27316 11520 27328
rect 11475 27288 11520 27316
rect 11514 27276 11520 27288
rect 11572 27276 11578 27328
rect 12986 27276 12992 27328
rect 13044 27316 13050 27328
rect 21818 27316 21824 27328
rect 13044 27288 21824 27316
rect 13044 27276 13050 27288
rect 21818 27276 21824 27288
rect 21876 27276 21882 27328
rect 23474 27276 23480 27328
rect 23532 27316 23538 27328
rect 23532 27288 23577 27316
rect 23532 27276 23538 27288
rect 24210 27276 24216 27328
rect 24268 27316 24274 27328
rect 24762 27316 24768 27328
rect 24268 27288 24768 27316
rect 24268 27276 24274 27288
rect 24762 27276 24768 27288
rect 24820 27276 24826 27328
rect 26418 27276 26424 27328
rect 26476 27316 26482 27328
rect 26605 27319 26663 27325
rect 26605 27316 26617 27319
rect 26476 27288 26617 27316
rect 26476 27276 26482 27288
rect 26605 27285 26617 27288
rect 26651 27285 26663 27319
rect 26605 27279 26663 27285
rect 27338 27276 27344 27328
rect 27396 27316 27402 27328
rect 27893 27319 27951 27325
rect 27893 27316 27905 27319
rect 27396 27288 27905 27316
rect 27396 27276 27402 27288
rect 27893 27285 27905 27288
rect 27939 27285 27951 27319
rect 27893 27279 27951 27285
rect 27982 27276 27988 27328
rect 28040 27316 28046 27328
rect 29825 27319 29883 27325
rect 29825 27316 29837 27319
rect 28040 27288 29837 27316
rect 28040 27276 28046 27288
rect 29825 27285 29837 27288
rect 29871 27285 29883 27319
rect 30466 27316 30472 27328
rect 30427 27288 30472 27316
rect 29825 27279 29883 27285
rect 30466 27276 30472 27288
rect 30524 27276 30530 27328
rect 38194 27316 38200 27328
rect 38155 27288 38200 27316
rect 38194 27276 38200 27288
rect 38252 27276 38258 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 20073 27115 20131 27121
rect 20073 27081 20085 27115
rect 20119 27112 20131 27115
rect 22002 27112 22008 27124
rect 20119 27084 22008 27112
rect 20119 27081 20131 27084
rect 20073 27075 20131 27081
rect 22002 27072 22008 27084
rect 22060 27072 22066 27124
rect 22094 27072 22100 27124
rect 22152 27112 22158 27124
rect 31570 27112 31576 27124
rect 22152 27084 25912 27112
rect 31531 27084 31576 27112
rect 22152 27072 22158 27084
rect 3697 27047 3755 27053
rect 3697 27013 3709 27047
rect 3743 27044 3755 27047
rect 3970 27044 3976 27056
rect 3743 27016 3976 27044
rect 3743 27013 3755 27016
rect 3697 27007 3755 27013
rect 3970 27004 3976 27016
rect 4028 27004 4034 27056
rect 4706 27004 4712 27056
rect 4764 27004 4770 27056
rect 13722 27044 13728 27056
rect 13683 27016 13728 27044
rect 13722 27004 13728 27016
rect 13780 27004 13786 27056
rect 17126 27044 17132 27056
rect 17087 27016 17132 27044
rect 17126 27004 17132 27016
rect 17184 27004 17190 27056
rect 19150 27044 19156 27056
rect 18354 27016 19156 27044
rect 19150 27004 19156 27016
rect 19208 27004 19214 27056
rect 19334 27004 19340 27056
rect 19392 27044 19398 27056
rect 22189 27047 22247 27053
rect 22189 27044 22201 27047
rect 19392 27016 22201 27044
rect 19392 27004 19398 27016
rect 22189 27013 22201 27016
rect 22235 27013 22247 27047
rect 22189 27007 22247 27013
rect 22462 27004 22468 27056
rect 22520 27044 22526 27056
rect 24210 27044 24216 27056
rect 22520 27016 24216 27044
rect 22520 27004 22526 27016
rect 24210 27004 24216 27016
rect 24268 27004 24274 27056
rect 24486 27044 24492 27056
rect 24447 27016 24492 27044
rect 24486 27004 24492 27016
rect 24544 27004 24550 27056
rect 1670 26976 1676 26988
rect 1631 26948 1676 26976
rect 1670 26936 1676 26948
rect 1728 26936 1734 26988
rect 11238 26936 11244 26988
rect 11296 26976 11302 26988
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11296 26948 11713 26976
rect 11296 26936 11302 26948
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 13078 26936 13084 26988
rect 13136 26936 13142 26988
rect 14185 26979 14243 26985
rect 14185 26945 14197 26979
rect 14231 26945 14243 26979
rect 16850 26976 16856 26988
rect 16811 26948 16856 26976
rect 14185 26939 14243 26945
rect 3421 26911 3479 26917
rect 3421 26877 3433 26911
rect 3467 26908 3479 26911
rect 3467 26880 3556 26908
rect 3467 26877 3479 26880
rect 3421 26871 3479 26877
rect 1854 26840 1860 26852
rect 1815 26812 1860 26840
rect 1854 26800 1860 26812
rect 1912 26800 1918 26852
rect 3528 26772 3556 26880
rect 9214 26868 9220 26920
rect 9272 26908 9278 26920
rect 11977 26911 12035 26917
rect 11977 26908 11989 26911
rect 9272 26880 11989 26908
rect 9272 26868 9278 26880
rect 11977 26877 11989 26880
rect 12023 26877 12035 26911
rect 11977 26871 12035 26877
rect 14200 26840 14228 26939
rect 16850 26936 16856 26948
rect 16908 26936 16914 26988
rect 18506 26936 18512 26988
rect 18564 26976 18570 26988
rect 18966 26976 18972 26988
rect 18564 26948 18972 26976
rect 18564 26936 18570 26948
rect 18966 26936 18972 26948
rect 19024 26976 19030 26988
rect 19061 26979 19119 26985
rect 19061 26976 19073 26979
rect 19024 26948 19073 26976
rect 19024 26936 19030 26948
rect 19061 26945 19073 26948
rect 19107 26945 19119 26979
rect 19061 26939 19119 26945
rect 19242 26936 19248 26988
rect 19300 26976 19306 26988
rect 25884 26985 25912 27084
rect 31570 27072 31576 27084
rect 31628 27072 31634 27124
rect 37829 27115 37887 27121
rect 37829 27081 37841 27115
rect 37875 27112 37887 27115
rect 38378 27112 38384 27124
rect 37875 27084 38384 27112
rect 37875 27081 37887 27084
rect 37829 27075 37887 27081
rect 38378 27072 38384 27084
rect 38436 27072 38442 27124
rect 27338 27044 27344 27056
rect 27299 27016 27344 27044
rect 27338 27004 27344 27016
rect 27396 27004 27402 27056
rect 19981 26979 20039 26985
rect 19981 26976 19993 26979
rect 19300 26948 19993 26976
rect 19300 26936 19306 26948
rect 19981 26945 19993 26948
rect 20027 26945 20039 26979
rect 19981 26939 20039 26945
rect 25869 26979 25927 26985
rect 25869 26945 25881 26979
rect 25915 26945 25927 26979
rect 25869 26939 25927 26945
rect 29178 26936 29184 26988
rect 29236 26976 29242 26988
rect 31481 26979 31539 26985
rect 31481 26976 31493 26979
rect 29236 26948 31493 26976
rect 29236 26936 29242 26948
rect 31481 26945 31493 26948
rect 31527 26945 31539 26979
rect 31481 26939 31539 26945
rect 37918 26936 37924 26988
rect 37976 26976 37982 26988
rect 38013 26979 38071 26985
rect 38013 26976 38025 26979
rect 37976 26948 38025 26976
rect 37976 26936 37982 26948
rect 38013 26945 38025 26948
rect 38059 26945 38071 26979
rect 38013 26939 38071 26945
rect 19337 26911 19395 26917
rect 19337 26908 19349 26911
rect 18524 26880 19349 26908
rect 14200 26812 16988 26840
rect 4062 26772 4068 26784
rect 3528 26744 4068 26772
rect 4062 26732 4068 26744
rect 4120 26732 4126 26784
rect 5169 26775 5227 26781
rect 5169 26741 5181 26775
rect 5215 26772 5227 26775
rect 5350 26772 5356 26784
rect 5215 26744 5356 26772
rect 5215 26741 5227 26744
rect 5169 26735 5227 26741
rect 5350 26732 5356 26744
rect 5408 26732 5414 26784
rect 11054 26732 11060 26784
rect 11112 26772 11118 26784
rect 14277 26775 14335 26781
rect 14277 26772 14289 26775
rect 11112 26744 14289 26772
rect 11112 26732 11118 26744
rect 14277 26741 14289 26744
rect 14323 26741 14335 26775
rect 16960 26772 16988 26812
rect 18524 26772 18552 26880
rect 19337 26877 19349 26880
rect 19383 26908 19395 26911
rect 19886 26908 19892 26920
rect 19383 26880 19892 26908
rect 19383 26877 19395 26880
rect 19337 26871 19395 26877
rect 19886 26868 19892 26880
rect 19944 26868 19950 26920
rect 21634 26908 21640 26920
rect 21284 26880 21640 26908
rect 18966 26800 18972 26852
rect 19024 26840 19030 26852
rect 21284 26840 21312 26880
rect 21634 26868 21640 26880
rect 21692 26868 21698 26920
rect 22005 26911 22063 26917
rect 22005 26877 22017 26911
rect 22051 26908 22063 26911
rect 23198 26908 23204 26920
rect 22051 26880 23204 26908
rect 22051 26877 22063 26880
rect 22005 26871 22063 26877
rect 23198 26868 23204 26880
rect 23256 26868 23262 26920
rect 23842 26908 23848 26920
rect 23803 26880 23848 26908
rect 23842 26868 23848 26880
rect 23900 26868 23906 26920
rect 24397 26911 24455 26917
rect 24397 26877 24409 26911
rect 24443 26877 24455 26911
rect 24397 26871 24455 26877
rect 19024 26812 21312 26840
rect 19024 26800 19030 26812
rect 21358 26800 21364 26852
rect 21416 26840 21422 26852
rect 24210 26840 24216 26852
rect 21416 26812 24216 26840
rect 21416 26800 21422 26812
rect 24210 26800 24216 26812
rect 24268 26800 24274 26852
rect 24412 26840 24440 26871
rect 24946 26868 24952 26920
rect 25004 26908 25010 26920
rect 25409 26911 25467 26917
rect 25409 26908 25421 26911
rect 25004 26880 25421 26908
rect 25004 26868 25010 26880
rect 25409 26877 25421 26880
rect 25455 26908 25467 26911
rect 26510 26908 26516 26920
rect 25455 26880 26516 26908
rect 25455 26877 25467 26880
rect 25409 26871 25467 26877
rect 26510 26868 26516 26880
rect 26568 26868 26574 26920
rect 27249 26911 27307 26917
rect 27249 26877 27261 26911
rect 27295 26908 27307 26911
rect 27890 26908 27896 26920
rect 27295 26880 27896 26908
rect 27295 26877 27307 26880
rect 27249 26871 27307 26877
rect 27890 26868 27896 26880
rect 27948 26868 27954 26920
rect 28166 26908 28172 26920
rect 28127 26880 28172 26908
rect 28166 26868 28172 26880
rect 28224 26868 28230 26920
rect 30466 26840 30472 26852
rect 24412 26812 30472 26840
rect 30466 26800 30472 26812
rect 30524 26800 30530 26852
rect 16960 26744 18552 26772
rect 18601 26775 18659 26781
rect 14277 26735 14335 26741
rect 18601 26741 18613 26775
rect 18647 26772 18659 26775
rect 18782 26772 18788 26784
rect 18647 26744 18788 26772
rect 18647 26741 18659 26744
rect 18601 26735 18659 26741
rect 18782 26732 18788 26744
rect 18840 26772 18846 26784
rect 21634 26772 21640 26784
rect 18840 26744 21640 26772
rect 18840 26732 18846 26744
rect 21634 26732 21640 26744
rect 21692 26772 21698 26784
rect 24578 26772 24584 26784
rect 21692 26744 24584 26772
rect 21692 26732 21698 26744
rect 24578 26732 24584 26744
rect 24636 26732 24642 26784
rect 25961 26775 26019 26781
rect 25961 26741 25973 26775
rect 26007 26772 26019 26775
rect 27522 26772 27528 26784
rect 26007 26744 27528 26772
rect 26007 26741 26019 26744
rect 25961 26735 26019 26741
rect 27522 26732 27528 26744
rect 27580 26732 27586 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 5442 26528 5448 26580
rect 5500 26568 5506 26580
rect 12986 26568 12992 26580
rect 5500 26540 12992 26568
rect 5500 26528 5506 26540
rect 12986 26528 12992 26540
rect 13044 26528 13050 26580
rect 13078 26528 13084 26580
rect 13136 26568 13142 26580
rect 21085 26571 21143 26577
rect 21085 26568 21097 26571
rect 13136 26540 21097 26568
rect 13136 26528 13142 26540
rect 21085 26537 21097 26540
rect 21131 26537 21143 26571
rect 21085 26531 21143 26537
rect 23934 26528 23940 26580
rect 23992 26568 23998 26580
rect 24673 26571 24731 26577
rect 24673 26568 24685 26571
rect 23992 26540 24685 26568
rect 23992 26528 23998 26540
rect 24673 26537 24685 26540
rect 24719 26537 24731 26571
rect 24673 26531 24731 26537
rect 26881 26571 26939 26577
rect 26881 26537 26893 26571
rect 26927 26568 26939 26571
rect 29178 26568 29184 26580
rect 26927 26540 29184 26568
rect 26927 26537 26939 26540
rect 26881 26531 26939 26537
rect 29178 26528 29184 26540
rect 29236 26528 29242 26580
rect 30374 26528 30380 26580
rect 30432 26568 30438 26580
rect 38105 26571 38163 26577
rect 38105 26568 38117 26571
rect 30432 26540 38117 26568
rect 30432 26528 30438 26540
rect 38105 26537 38117 26540
rect 38151 26537 38163 26571
rect 38105 26531 38163 26537
rect 11977 26503 12035 26509
rect 11977 26469 11989 26503
rect 12023 26500 12035 26503
rect 15746 26500 15752 26512
rect 12023 26472 15752 26500
rect 12023 26469 12035 26472
rect 11977 26463 12035 26469
rect 15746 26460 15752 26472
rect 15804 26460 15810 26512
rect 19242 26500 19248 26512
rect 18432 26472 19248 26500
rect 2406 26432 2412 26444
rect 2367 26404 2412 26432
rect 2406 26392 2412 26404
rect 2464 26392 2470 26444
rect 7926 26392 7932 26444
rect 7984 26432 7990 26444
rect 8021 26435 8079 26441
rect 8021 26432 8033 26435
rect 7984 26404 8033 26432
rect 7984 26392 7990 26404
rect 8021 26401 8033 26404
rect 8067 26401 8079 26435
rect 8021 26395 8079 26401
rect 10229 26435 10287 26441
rect 10229 26401 10241 26435
rect 10275 26432 10287 26435
rect 12250 26432 12256 26444
rect 10275 26404 12256 26432
rect 10275 26401 10287 26404
rect 10229 26395 10287 26401
rect 6086 26324 6092 26376
rect 6144 26364 6150 26376
rect 6273 26367 6331 26373
rect 6273 26364 6285 26367
rect 6144 26336 6285 26364
rect 6144 26324 6150 26336
rect 6273 26333 6285 26336
rect 6319 26333 6331 26367
rect 6273 26327 6331 26333
rect 2501 26299 2559 26305
rect 2501 26265 2513 26299
rect 2547 26296 2559 26299
rect 2866 26296 2872 26308
rect 2547 26268 2872 26296
rect 2547 26265 2559 26268
rect 2501 26259 2559 26265
rect 2866 26256 2872 26268
rect 2924 26256 2930 26308
rect 3418 26296 3424 26308
rect 3379 26268 3424 26296
rect 3418 26256 3424 26268
rect 3476 26256 3482 26308
rect 6549 26299 6607 26305
rect 6549 26265 6561 26299
rect 6595 26296 6607 26299
rect 6638 26296 6644 26308
rect 6595 26268 6644 26296
rect 6595 26265 6607 26268
rect 6549 26259 6607 26265
rect 6638 26256 6644 26268
rect 6696 26256 6702 26308
rect 7006 26256 7012 26308
rect 7064 26256 7070 26308
rect 8036 26296 8064 26395
rect 12250 26392 12256 26404
rect 12308 26392 12314 26444
rect 16577 26435 16635 26441
rect 16577 26401 16589 26435
rect 16623 26432 16635 26435
rect 16850 26432 16856 26444
rect 16623 26404 16856 26432
rect 16623 26401 16635 26404
rect 16577 26395 16635 26401
rect 16850 26392 16856 26404
rect 16908 26392 16914 26444
rect 17310 26392 17316 26444
rect 17368 26432 17374 26444
rect 18432 26432 18460 26472
rect 19242 26460 19248 26472
rect 19300 26460 19306 26512
rect 19521 26503 19579 26509
rect 19521 26469 19533 26503
rect 19567 26500 19579 26503
rect 19978 26500 19984 26512
rect 19567 26472 19984 26500
rect 19567 26469 19579 26472
rect 19521 26463 19579 26469
rect 19978 26460 19984 26472
rect 20036 26460 20042 26512
rect 29733 26503 29791 26509
rect 25332 26472 26556 26500
rect 20162 26432 20168 26444
rect 17368 26404 18460 26432
rect 18708 26404 20168 26432
rect 17368 26392 17374 26404
rect 18708 26364 18736 26404
rect 20162 26392 20168 26404
rect 20220 26392 20226 26444
rect 22738 26392 22744 26444
rect 22796 26432 22802 26444
rect 25332 26432 25360 26472
rect 26418 26432 26424 26444
rect 22796 26404 25360 26432
rect 26379 26404 26424 26432
rect 22796 26392 22802 26404
rect 17986 26336 18736 26364
rect 18782 26324 18788 26376
rect 18840 26364 18846 26376
rect 19421 26367 19479 26373
rect 19421 26364 19433 26367
rect 18840 26336 19433 26364
rect 18840 26324 18846 26336
rect 19421 26333 19433 26336
rect 19467 26333 19479 26367
rect 20070 26364 20076 26376
rect 19421 26327 19479 26333
rect 19536 26336 20076 26364
rect 10502 26296 10508 26308
rect 8036 26268 10508 26296
rect 10502 26256 10508 26268
rect 10560 26256 10566 26308
rect 11146 26256 11152 26308
rect 11204 26256 11210 26308
rect 16574 26256 16580 26308
rect 16632 26296 16638 26308
rect 16853 26299 16911 26305
rect 16853 26296 16865 26299
rect 16632 26268 16865 26296
rect 16632 26256 16638 26268
rect 16853 26265 16865 26268
rect 16899 26296 16911 26299
rect 16942 26296 16948 26308
rect 16899 26268 16948 26296
rect 16899 26265 16911 26268
rect 16853 26259 16911 26265
rect 16942 26256 16948 26268
rect 17000 26256 17006 26308
rect 18601 26299 18659 26305
rect 18601 26265 18613 26299
rect 18647 26296 18659 26299
rect 19242 26296 19248 26308
rect 18647 26268 19248 26296
rect 18647 26265 18659 26268
rect 18601 26259 18659 26265
rect 19242 26256 19248 26268
rect 19300 26296 19306 26308
rect 19536 26296 19564 26336
rect 20070 26324 20076 26336
rect 20128 26324 20134 26376
rect 20346 26324 20352 26376
rect 20404 26364 20410 26376
rect 20993 26367 21051 26373
rect 20404 26336 20449 26364
rect 20404 26324 20410 26336
rect 20993 26333 21005 26367
rect 21039 26364 21051 26367
rect 21637 26367 21695 26373
rect 21637 26364 21649 26367
rect 21039 26336 21649 26364
rect 21039 26333 21051 26336
rect 20993 26327 21051 26333
rect 21637 26333 21649 26336
rect 21683 26364 21695 26367
rect 22462 26364 22468 26376
rect 21683 26336 22468 26364
rect 21683 26333 21695 26336
rect 21637 26327 21695 26333
rect 22462 26324 22468 26336
rect 22520 26324 22526 26376
rect 22646 26324 22652 26376
rect 22704 26364 22710 26376
rect 22830 26364 22836 26376
rect 22704 26336 22836 26364
rect 22704 26324 22710 26336
rect 22830 26324 22836 26336
rect 22888 26324 22894 26376
rect 23308 26373 23336 26404
rect 26418 26392 26424 26404
rect 26476 26392 26482 26444
rect 26528 26432 26556 26472
rect 29733 26469 29745 26503
rect 29779 26500 29791 26503
rect 38010 26500 38016 26512
rect 29779 26472 38016 26500
rect 29779 26469 29791 26472
rect 29733 26463 29791 26469
rect 38010 26460 38016 26472
rect 38068 26460 38074 26512
rect 36354 26432 36360 26444
rect 26528 26404 36360 26432
rect 36354 26392 36360 26404
rect 36412 26392 36418 26444
rect 23293 26367 23351 26373
rect 23293 26333 23305 26367
rect 23339 26333 23351 26367
rect 23293 26327 23351 26333
rect 23382 26324 23388 26376
rect 23440 26364 23446 26376
rect 23440 26336 23485 26364
rect 23440 26324 23446 26336
rect 24486 26324 24492 26376
rect 24544 26366 24550 26376
rect 24581 26367 24639 26373
rect 24581 26366 24593 26367
rect 24544 26338 24593 26366
rect 24544 26324 24550 26338
rect 24581 26333 24593 26338
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 25038 26324 25044 26376
rect 25096 26364 25102 26376
rect 25225 26367 25283 26373
rect 25225 26364 25237 26367
rect 25096 26336 25237 26364
rect 25096 26324 25102 26336
rect 25225 26333 25237 26336
rect 25271 26333 25283 26367
rect 25225 26327 25283 26333
rect 26237 26367 26295 26373
rect 26237 26333 26249 26367
rect 26283 26364 26295 26367
rect 26510 26364 26516 26376
rect 26283 26336 26516 26364
rect 26283 26333 26295 26336
rect 26237 26327 26295 26333
rect 26510 26324 26516 26336
rect 26568 26324 26574 26376
rect 28534 26364 28540 26376
rect 28495 26336 28540 26364
rect 28534 26324 28540 26336
rect 28592 26324 28598 26376
rect 28718 26364 28724 26376
rect 28679 26336 28724 26364
rect 28718 26324 28724 26336
rect 28776 26324 28782 26376
rect 29086 26324 29092 26376
rect 29144 26364 29150 26376
rect 29917 26367 29975 26373
rect 29917 26364 29929 26367
rect 29144 26336 29929 26364
rect 29144 26324 29150 26336
rect 29917 26333 29929 26336
rect 29963 26333 29975 26367
rect 38286 26364 38292 26376
rect 38247 26336 38292 26364
rect 29917 26327 29975 26333
rect 38286 26324 38292 26336
rect 38344 26324 38350 26376
rect 20438 26296 20444 26308
rect 19300 26268 19564 26296
rect 20399 26268 20444 26296
rect 19300 26256 19306 26268
rect 20438 26256 20444 26268
rect 20496 26256 20502 26308
rect 21729 26299 21787 26305
rect 21729 26296 21741 26299
rect 20732 26268 21741 26296
rect 17218 26188 17224 26240
rect 17276 26228 17282 26240
rect 20732 26228 20760 26268
rect 21729 26265 21741 26268
rect 21775 26265 21787 26299
rect 21729 26259 21787 26265
rect 22741 26299 22799 26305
rect 22741 26265 22753 26299
rect 22787 26296 22799 26299
rect 24762 26296 24768 26308
rect 22787 26268 24768 26296
rect 22787 26265 22799 26268
rect 22741 26259 22799 26265
rect 24762 26256 24768 26268
rect 24820 26256 24826 26308
rect 17276 26200 20760 26228
rect 17276 26188 17282 26200
rect 22278 26188 22284 26240
rect 22336 26228 22342 26240
rect 24946 26228 24952 26240
rect 22336 26200 24952 26228
rect 22336 26188 22342 26200
rect 24946 26188 24952 26200
rect 25004 26188 25010 26240
rect 25314 26228 25320 26240
rect 25275 26200 25320 26228
rect 25314 26188 25320 26200
rect 25372 26188 25378 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 10778 26024 10784 26036
rect 10739 25996 10784 26024
rect 10778 25984 10784 25996
rect 10836 25984 10842 26036
rect 18414 26024 18420 26036
rect 12912 25996 18420 26024
rect 3878 25916 3884 25968
rect 3936 25956 3942 25968
rect 12912 25956 12940 25996
rect 18414 25984 18420 25996
rect 18472 25984 18478 26036
rect 19150 26024 19156 26036
rect 19111 25996 19156 26024
rect 19150 25984 19156 25996
rect 19208 25984 19214 26036
rect 24486 26024 24492 26036
rect 22066 25996 24492 26024
rect 17218 25956 17224 25968
rect 3936 25928 4922 25956
rect 10534 25928 12940 25956
rect 13754 25928 17224 25956
rect 3936 25916 3942 25928
rect 17218 25916 17224 25928
rect 17276 25916 17282 25968
rect 20438 25956 20444 25968
rect 18354 25928 20444 25956
rect 20438 25916 20444 25928
rect 20496 25916 20502 25968
rect 20530 25916 20536 25968
rect 20588 25956 20594 25968
rect 22066 25956 22094 25996
rect 24486 25984 24492 25996
rect 24544 25984 24550 26036
rect 28534 25984 28540 26036
rect 28592 26024 28598 26036
rect 28721 26027 28779 26033
rect 28721 26024 28733 26027
rect 28592 25996 28733 26024
rect 28592 25984 28598 25996
rect 28721 25993 28733 25996
rect 28767 25993 28779 26027
rect 28721 25987 28779 25993
rect 20588 25928 22094 25956
rect 20588 25916 20594 25928
rect 23474 25916 23480 25968
rect 23532 25956 23538 25968
rect 24765 25959 24823 25965
rect 24765 25956 24777 25959
rect 23532 25928 24777 25956
rect 23532 25916 23538 25928
rect 24765 25925 24777 25928
rect 24811 25925 24823 25959
rect 24765 25919 24823 25925
rect 25685 25959 25743 25965
rect 25685 25925 25697 25959
rect 25731 25956 25743 25959
rect 26602 25956 26608 25968
rect 25731 25928 26608 25956
rect 25731 25925 25743 25928
rect 25685 25919 25743 25925
rect 26602 25916 26608 25928
rect 26660 25916 26666 25968
rect 27522 25916 27528 25968
rect 27580 25956 27586 25968
rect 29917 25959 29975 25965
rect 29917 25956 29929 25959
rect 27580 25928 29929 25956
rect 27580 25916 27586 25928
rect 29917 25925 29929 25928
rect 29963 25925 29975 25959
rect 29917 25919 29975 25925
rect 3513 25891 3571 25897
rect 3513 25857 3525 25891
rect 3559 25888 3571 25891
rect 3786 25888 3792 25900
rect 3559 25860 3792 25888
rect 3559 25857 3571 25860
rect 3513 25851 3571 25857
rect 3786 25848 3792 25860
rect 3844 25848 3850 25900
rect 12250 25888 12256 25900
rect 12211 25860 12256 25888
rect 12250 25848 12256 25860
rect 12308 25848 12314 25900
rect 18782 25848 18788 25900
rect 18840 25888 18846 25900
rect 19061 25891 19119 25897
rect 19061 25888 19073 25891
rect 18840 25860 19073 25888
rect 18840 25848 18846 25860
rect 19061 25857 19073 25860
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 19150 25848 19156 25900
rect 19208 25888 19214 25900
rect 19705 25891 19763 25897
rect 19705 25888 19717 25891
rect 19208 25860 19717 25888
rect 19208 25848 19214 25860
rect 19705 25857 19717 25860
rect 19751 25857 19763 25891
rect 22278 25888 22284 25900
rect 22239 25860 22284 25888
rect 19705 25851 19763 25857
rect 22278 25848 22284 25860
rect 22336 25848 22342 25900
rect 26145 25891 26203 25897
rect 26145 25857 26157 25891
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 4062 25780 4068 25832
rect 4120 25820 4126 25832
rect 4157 25823 4215 25829
rect 4157 25820 4169 25823
rect 4120 25792 4169 25820
rect 4120 25780 4126 25792
rect 4157 25789 4169 25792
rect 4203 25789 4215 25823
rect 4157 25783 4215 25789
rect 4433 25823 4491 25829
rect 4433 25789 4445 25823
rect 4479 25820 4491 25823
rect 4522 25820 4528 25832
rect 4479 25792 4528 25820
rect 4479 25789 4491 25792
rect 4433 25783 4491 25789
rect 4522 25780 4528 25792
rect 4580 25780 4586 25832
rect 6086 25780 6092 25832
rect 6144 25820 6150 25832
rect 7466 25820 7472 25832
rect 6144 25792 7472 25820
rect 6144 25780 6150 25792
rect 7466 25780 7472 25792
rect 7524 25820 7530 25832
rect 9033 25823 9091 25829
rect 9033 25820 9045 25823
rect 7524 25792 9045 25820
rect 7524 25780 7530 25792
rect 9033 25789 9045 25792
rect 9079 25789 9091 25823
rect 9033 25783 9091 25789
rect 9309 25823 9367 25829
rect 9309 25789 9321 25823
rect 9355 25820 9367 25823
rect 9950 25820 9956 25832
rect 9355 25792 9956 25820
rect 9355 25789 9367 25792
rect 9309 25783 9367 25789
rect 9950 25780 9956 25792
rect 10008 25820 10014 25832
rect 12529 25823 12587 25829
rect 10008 25792 10548 25820
rect 10008 25780 10014 25792
rect 3605 25687 3663 25693
rect 3605 25653 3617 25687
rect 3651 25684 3663 25687
rect 3694 25684 3700 25696
rect 3651 25656 3700 25684
rect 3651 25653 3663 25656
rect 3605 25647 3663 25653
rect 3694 25644 3700 25656
rect 3752 25644 3758 25696
rect 5905 25687 5963 25693
rect 5905 25653 5917 25687
rect 5951 25684 5963 25687
rect 6638 25684 6644 25696
rect 5951 25656 6644 25684
rect 5951 25653 5963 25656
rect 5905 25647 5963 25653
rect 6638 25644 6644 25656
rect 6696 25644 6702 25696
rect 10520 25684 10548 25792
rect 12529 25789 12541 25823
rect 12575 25820 12587 25823
rect 12618 25820 12624 25832
rect 12575 25792 12624 25820
rect 12575 25789 12587 25792
rect 12529 25783 12587 25789
rect 12618 25780 12624 25792
rect 12676 25780 12682 25832
rect 12894 25780 12900 25832
rect 12952 25820 12958 25832
rect 14277 25823 14335 25829
rect 14277 25820 14289 25823
rect 12952 25792 14289 25820
rect 12952 25780 12958 25792
rect 14277 25789 14289 25792
rect 14323 25820 14335 25823
rect 16022 25820 16028 25832
rect 14323 25792 16028 25820
rect 14323 25789 14335 25792
rect 14277 25783 14335 25789
rect 16022 25780 16028 25792
rect 16080 25780 16086 25832
rect 16850 25820 16856 25832
rect 16811 25792 16856 25820
rect 16850 25780 16856 25792
rect 16908 25780 16914 25832
rect 17129 25823 17187 25829
rect 17129 25789 17141 25823
rect 17175 25820 17187 25823
rect 18138 25820 18144 25832
rect 17175 25792 18144 25820
rect 17175 25789 17187 25792
rect 17129 25783 17187 25789
rect 18138 25780 18144 25792
rect 18196 25780 18202 25832
rect 18414 25780 18420 25832
rect 18472 25820 18478 25832
rect 22462 25820 22468 25832
rect 18472 25792 22094 25820
rect 22423 25792 22468 25820
rect 18472 25780 18478 25792
rect 18322 25712 18328 25764
rect 18380 25752 18386 25764
rect 22066 25752 22094 25792
rect 22462 25780 22468 25792
rect 22520 25780 22526 25832
rect 24121 25823 24179 25829
rect 24121 25789 24133 25823
rect 24167 25820 24179 25823
rect 24210 25820 24216 25832
rect 24167 25792 24216 25820
rect 24167 25789 24179 25792
rect 24121 25783 24179 25789
rect 24210 25780 24216 25792
rect 24268 25780 24274 25832
rect 24302 25780 24308 25832
rect 24360 25820 24366 25832
rect 24673 25823 24731 25829
rect 24673 25820 24685 25823
rect 24360 25792 24685 25820
rect 24360 25780 24366 25792
rect 24673 25789 24685 25792
rect 24719 25789 24731 25823
rect 24673 25783 24731 25789
rect 25314 25752 25320 25764
rect 18380 25724 19932 25752
rect 22066 25724 25320 25752
rect 18380 25712 18386 25724
rect 18230 25684 18236 25696
rect 10520 25656 18236 25684
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 18598 25684 18604 25696
rect 18559 25656 18604 25684
rect 18598 25644 18604 25656
rect 18656 25644 18662 25696
rect 18690 25644 18696 25696
rect 18748 25684 18754 25696
rect 19797 25687 19855 25693
rect 19797 25684 19809 25687
rect 18748 25656 19809 25684
rect 18748 25644 18754 25656
rect 19797 25653 19809 25656
rect 19843 25653 19855 25687
rect 19904 25684 19932 25724
rect 25314 25712 25320 25724
rect 25372 25712 25378 25764
rect 26160 25684 26188 25851
rect 29825 25823 29883 25829
rect 29825 25789 29837 25823
rect 29871 25820 29883 25823
rect 29914 25820 29920 25832
rect 29871 25792 29920 25820
rect 29871 25789 29883 25792
rect 29825 25783 29883 25789
rect 29914 25780 29920 25792
rect 29972 25780 29978 25832
rect 30834 25820 30840 25832
rect 30795 25792 30840 25820
rect 30834 25780 30840 25792
rect 30892 25780 30898 25832
rect 19904 25656 26188 25684
rect 26237 25687 26295 25693
rect 19797 25647 19855 25653
rect 26237 25653 26249 25687
rect 26283 25684 26295 25687
rect 30282 25684 30288 25696
rect 26283 25656 30288 25684
rect 26283 25653 26295 25656
rect 26237 25647 26295 25653
rect 30282 25644 30288 25656
rect 30340 25644 30346 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 15000 25483 15058 25489
rect 15000 25449 15012 25483
rect 15046 25480 15058 25483
rect 18598 25480 18604 25492
rect 15046 25452 18604 25480
rect 15046 25449 15058 25452
rect 15000 25443 15058 25449
rect 18598 25440 18604 25452
rect 18656 25440 18662 25492
rect 22373 25483 22431 25489
rect 19996 25452 22324 25480
rect 16022 25372 16028 25424
rect 16080 25412 16086 25424
rect 19058 25412 19064 25424
rect 16080 25384 19064 25412
rect 16080 25372 16086 25384
rect 19058 25372 19064 25384
rect 19116 25372 19122 25424
rect 19150 25372 19156 25424
rect 19208 25412 19214 25424
rect 19886 25412 19892 25424
rect 19208 25384 19892 25412
rect 19208 25372 19214 25384
rect 19886 25372 19892 25384
rect 19944 25372 19950 25424
rect 6086 25344 6092 25356
rect 6047 25316 6092 25344
rect 6086 25304 6092 25316
rect 6144 25304 6150 25356
rect 8018 25304 8024 25356
rect 8076 25344 8082 25356
rect 19996 25344 20024 25452
rect 8076 25316 20024 25344
rect 8076 25304 8082 25316
rect 20162 25304 20168 25356
rect 20220 25344 20226 25356
rect 22296 25344 22324 25452
rect 22373 25449 22385 25483
rect 22419 25480 22431 25483
rect 23658 25480 23664 25492
rect 22419 25452 23664 25480
rect 22419 25449 22431 25452
rect 22373 25443 22431 25449
rect 23658 25440 23664 25452
rect 23716 25440 23722 25492
rect 25314 25440 25320 25492
rect 25372 25480 25378 25492
rect 27798 25480 27804 25492
rect 25372 25452 27804 25480
rect 25372 25440 25378 25452
rect 27798 25440 27804 25452
rect 27856 25480 27862 25492
rect 28258 25480 28264 25492
rect 27856 25452 28264 25480
rect 27856 25440 27862 25452
rect 28258 25440 28264 25452
rect 28316 25440 28322 25492
rect 28718 25440 28724 25492
rect 28776 25480 28782 25492
rect 28813 25483 28871 25489
rect 28813 25480 28825 25483
rect 28776 25452 28825 25480
rect 28776 25440 28782 25452
rect 28813 25449 28825 25452
rect 28859 25449 28871 25483
rect 28813 25443 28871 25449
rect 23290 25372 23296 25424
rect 23348 25412 23354 25424
rect 26513 25415 26571 25421
rect 26513 25412 26525 25415
rect 23348 25384 26525 25412
rect 23348 25372 23354 25384
rect 26513 25381 26525 25384
rect 26559 25412 26571 25415
rect 26786 25412 26792 25424
rect 26559 25384 26792 25412
rect 26559 25381 26571 25384
rect 26513 25375 26571 25381
rect 26786 25372 26792 25384
rect 26844 25372 26850 25424
rect 29086 25344 29092 25356
rect 20220 25316 20265 25344
rect 22296 25316 29092 25344
rect 20220 25304 20226 25316
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 3602 25236 3608 25288
rect 3660 25276 3666 25288
rect 4062 25276 4068 25288
rect 3660 25248 4068 25276
rect 3660 25236 3666 25248
rect 4062 25236 4068 25248
rect 4120 25276 4126 25288
rect 4893 25279 4951 25285
rect 4893 25276 4905 25279
rect 4120 25248 4905 25276
rect 4120 25236 4126 25248
rect 4893 25245 4905 25248
rect 4939 25245 4951 25279
rect 4893 25239 4951 25245
rect 14274 25236 14280 25288
rect 14332 25276 14338 25288
rect 14737 25279 14795 25285
rect 14737 25276 14749 25279
rect 14332 25248 14749 25276
rect 14332 25236 14338 25248
rect 14737 25245 14749 25248
rect 14783 25245 14795 25279
rect 18046 25276 18052 25288
rect 18007 25248 18052 25276
rect 14737 25239 14795 25245
rect 18046 25236 18052 25248
rect 18104 25236 18110 25288
rect 18230 25236 18236 25288
rect 18288 25276 18294 25288
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 18288 25248 19441 25276
rect 18288 25236 18294 25248
rect 19429 25245 19441 25248
rect 19475 25245 19487 25279
rect 21634 25276 21640 25288
rect 21595 25248 21640 25276
rect 19429 25239 19487 25245
rect 21634 25236 21640 25248
rect 21692 25236 21698 25288
rect 22278 25276 22284 25288
rect 22239 25248 22284 25276
rect 22278 25236 22284 25248
rect 22336 25236 22342 25288
rect 22925 25279 22983 25285
rect 22925 25245 22937 25279
rect 22971 25276 22983 25279
rect 23106 25276 23112 25288
rect 22971 25248 23112 25276
rect 22971 25245 22983 25248
rect 22925 25239 22983 25245
rect 23106 25236 23112 25248
rect 23164 25236 23170 25288
rect 23474 25236 23480 25288
rect 23532 25276 23538 25288
rect 23569 25279 23627 25285
rect 23569 25276 23581 25279
rect 23532 25248 23581 25276
rect 23532 25236 23538 25248
rect 23569 25245 23581 25248
rect 23615 25245 23627 25279
rect 23569 25239 23627 25245
rect 25314 25236 25320 25288
rect 25372 25276 25378 25288
rect 25372 25248 25417 25276
rect 25372 25236 25378 25248
rect 25498 25236 25504 25288
rect 25556 25276 25562 25288
rect 26436 25285 26464 25316
rect 29086 25304 29092 25316
rect 29144 25304 29150 25356
rect 29914 25344 29920 25356
rect 29875 25316 29920 25344
rect 29914 25304 29920 25316
rect 29972 25304 29978 25356
rect 25777 25279 25835 25285
rect 25777 25276 25789 25279
rect 25556 25248 25789 25276
rect 25556 25236 25562 25248
rect 25777 25245 25789 25248
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 26421 25279 26479 25285
rect 26421 25245 26433 25279
rect 26467 25245 26479 25279
rect 27062 25276 27068 25288
rect 27023 25248 27068 25276
rect 26421 25239 26479 25245
rect 27062 25236 27068 25248
rect 27120 25236 27126 25288
rect 28350 25276 28356 25288
rect 28311 25248 28356 25276
rect 28350 25236 28356 25248
rect 28408 25236 28414 25288
rect 28997 25279 29055 25285
rect 28997 25245 29009 25279
rect 29043 25245 29055 25279
rect 28997 25239 29055 25245
rect 31481 25279 31539 25285
rect 31481 25245 31493 25279
rect 31527 25276 31539 25279
rect 31754 25276 31760 25288
rect 31527 25248 31760 25276
rect 31527 25245 31539 25248
rect 31481 25239 31539 25245
rect 4157 25211 4215 25217
rect 4157 25177 4169 25211
rect 4203 25208 4215 25211
rect 5626 25208 5632 25220
rect 4203 25180 5632 25208
rect 4203 25177 4215 25180
rect 4157 25171 4215 25177
rect 5626 25168 5632 25180
rect 5684 25168 5690 25220
rect 6362 25208 6368 25220
rect 6323 25180 6368 25208
rect 6362 25168 6368 25180
rect 6420 25168 6426 25220
rect 11054 25208 11060 25220
rect 7590 25180 11060 25208
rect 11054 25168 11060 25180
rect 11112 25168 11118 25220
rect 18141 25211 18199 25217
rect 16238 25180 18092 25208
rect 1762 25140 1768 25152
rect 1723 25112 1768 25140
rect 1762 25100 1768 25112
rect 1820 25100 1826 25152
rect 7098 25100 7104 25152
rect 7156 25140 7162 25152
rect 7837 25143 7895 25149
rect 7837 25140 7849 25143
rect 7156 25112 7849 25140
rect 7156 25100 7162 25112
rect 7837 25109 7849 25112
rect 7883 25109 7895 25143
rect 16482 25140 16488 25152
rect 16443 25112 16488 25140
rect 7837 25103 7895 25109
rect 16482 25100 16488 25112
rect 16540 25100 16546 25152
rect 18064 25140 18092 25180
rect 18141 25177 18153 25211
rect 18187 25208 18199 25211
rect 19794 25208 19800 25220
rect 18187 25180 19800 25208
rect 18187 25177 18199 25180
rect 18141 25171 18199 25177
rect 19794 25168 19800 25180
rect 19852 25168 19858 25220
rect 20257 25211 20315 25217
rect 20257 25177 20269 25211
rect 20303 25208 20315 25211
rect 20438 25208 20444 25220
rect 20303 25180 20444 25208
rect 20303 25177 20315 25180
rect 20257 25171 20315 25177
rect 20438 25168 20444 25180
rect 20496 25168 20502 25220
rect 21174 25208 21180 25220
rect 21135 25180 21180 25208
rect 21174 25168 21180 25180
rect 21232 25168 21238 25220
rect 21358 25168 21364 25220
rect 21416 25208 21422 25220
rect 23661 25211 23719 25217
rect 23661 25208 23673 25211
rect 21416 25180 23673 25208
rect 21416 25168 21422 25180
rect 23661 25177 23673 25180
rect 23707 25177 23719 25211
rect 23661 25171 23719 25177
rect 23842 25168 23848 25220
rect 23900 25208 23906 25220
rect 24486 25208 24492 25220
rect 23900 25180 24492 25208
rect 23900 25168 23906 25180
rect 24486 25168 24492 25180
rect 24544 25208 24550 25220
rect 24673 25211 24731 25217
rect 24673 25208 24685 25211
rect 24544 25180 24685 25208
rect 24544 25168 24550 25180
rect 24673 25177 24685 25180
rect 24719 25177 24731 25211
rect 24673 25171 24731 25177
rect 24762 25168 24768 25220
rect 24820 25208 24826 25220
rect 29012 25208 29040 25239
rect 31754 25236 31760 25248
rect 31812 25236 31818 25288
rect 24820 25180 24865 25208
rect 28184 25180 29040 25208
rect 24820 25168 24826 25180
rect 19242 25140 19248 25152
rect 18064 25112 19248 25140
rect 19242 25100 19248 25112
rect 19300 25100 19306 25152
rect 19521 25143 19579 25149
rect 19521 25109 19533 25143
rect 19567 25140 19579 25143
rect 19978 25140 19984 25152
rect 19567 25112 19984 25140
rect 19567 25109 19579 25112
rect 19521 25103 19579 25109
rect 19978 25100 19984 25112
rect 20036 25100 20042 25152
rect 21729 25143 21787 25149
rect 21729 25109 21741 25143
rect 21775 25140 21787 25143
rect 21910 25140 21916 25152
rect 21775 25112 21916 25140
rect 21775 25109 21787 25112
rect 21729 25103 21787 25109
rect 21910 25100 21916 25112
rect 21968 25100 21974 25152
rect 23017 25143 23075 25149
rect 23017 25109 23029 25143
rect 23063 25140 23075 25143
rect 23566 25140 23572 25152
rect 23063 25112 23572 25140
rect 23063 25109 23075 25112
rect 23017 25103 23075 25109
rect 23566 25100 23572 25112
rect 23624 25100 23630 25152
rect 24854 25100 24860 25152
rect 24912 25140 24918 25152
rect 25869 25143 25927 25149
rect 25869 25140 25881 25143
rect 24912 25112 25881 25140
rect 24912 25100 24918 25112
rect 25869 25109 25881 25112
rect 25915 25109 25927 25143
rect 27154 25140 27160 25152
rect 27115 25112 27160 25140
rect 25869 25103 25927 25109
rect 27154 25100 27160 25112
rect 27212 25100 27218 25152
rect 28184 25149 28212 25180
rect 28169 25143 28227 25149
rect 28169 25109 28181 25143
rect 28215 25109 28227 25143
rect 31570 25140 31576 25152
rect 31531 25112 31576 25140
rect 28169 25103 28227 25109
rect 31570 25100 31576 25112
rect 31628 25100 31634 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 5353 24939 5411 24945
rect 5353 24905 5365 24939
rect 5399 24905 5411 24939
rect 5353 24899 5411 24905
rect 4614 24828 4620 24880
rect 4672 24828 4678 24880
rect 1394 24760 1400 24812
rect 1452 24800 1458 24812
rect 1765 24803 1823 24809
rect 1765 24800 1777 24803
rect 1452 24772 1777 24800
rect 1452 24760 1458 24772
rect 1765 24769 1777 24772
rect 1811 24769 1823 24803
rect 5368 24800 5396 24899
rect 16298 24896 16304 24948
rect 16356 24936 16362 24948
rect 18046 24936 18052 24948
rect 16356 24908 18052 24936
rect 16356 24896 16362 24908
rect 18046 24896 18052 24908
rect 18104 24896 18110 24948
rect 18138 24896 18144 24948
rect 18196 24936 18202 24948
rect 23106 24936 23112 24948
rect 18196 24908 23112 24936
rect 18196 24896 18202 24908
rect 23106 24896 23112 24908
rect 23164 24896 23170 24948
rect 24210 24896 24216 24948
rect 24268 24936 24274 24948
rect 27890 24936 27896 24948
rect 24268 24908 27896 24936
rect 24268 24896 24274 24908
rect 27890 24896 27896 24908
rect 27948 24896 27954 24948
rect 16482 24828 16488 24880
rect 16540 24868 16546 24880
rect 16540 24840 17632 24868
rect 16540 24828 16546 24840
rect 7742 24800 7748 24812
rect 5368 24772 7748 24800
rect 1765 24763 1823 24769
rect 7742 24760 7748 24772
rect 7800 24760 7806 24812
rect 3602 24732 3608 24744
rect 3563 24704 3608 24732
rect 3602 24692 3608 24704
rect 3660 24692 3666 24744
rect 3881 24735 3939 24741
rect 3881 24701 3893 24735
rect 3927 24732 3939 24735
rect 13262 24732 13268 24744
rect 3927 24704 6868 24732
rect 13223 24704 13268 24732
rect 3927 24701 3939 24704
rect 3881 24695 3939 24701
rect 6840 24608 6868 24704
rect 13262 24692 13268 24704
rect 13320 24692 13326 24744
rect 13541 24735 13599 24741
rect 13541 24701 13553 24735
rect 13587 24732 13599 24735
rect 14182 24732 14188 24744
rect 13587 24704 14188 24732
rect 13587 24701 13599 24704
rect 13541 24695 13599 24701
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 14660 24664 14688 24786
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 16853 24803 16911 24809
rect 16853 24800 16865 24803
rect 15252 24772 16865 24800
rect 15252 24760 15258 24772
rect 16853 24769 16865 24772
rect 16899 24800 16911 24803
rect 17494 24800 17500 24812
rect 16899 24772 17500 24800
rect 16899 24769 16911 24772
rect 16853 24763 16911 24769
rect 17494 24760 17500 24772
rect 17552 24760 17558 24812
rect 17604 24800 17632 24840
rect 18248 24840 19104 24868
rect 18248 24800 18276 24840
rect 17604 24772 18276 24800
rect 18322 24760 18328 24812
rect 18380 24800 18386 24812
rect 18969 24803 19027 24809
rect 18380 24772 18425 24800
rect 18380 24760 18386 24772
rect 18969 24769 18981 24803
rect 19015 24769 19027 24803
rect 19076 24800 19104 24840
rect 20070 24828 20076 24880
rect 20128 24868 20134 24880
rect 20441 24871 20499 24877
rect 20441 24868 20453 24871
rect 20128 24840 20453 24868
rect 20128 24828 20134 24840
rect 20441 24837 20453 24840
rect 20487 24837 20499 24871
rect 20441 24831 20499 24837
rect 23566 24828 23572 24880
rect 23624 24868 23630 24880
rect 24029 24871 24087 24877
rect 24029 24868 24041 24871
rect 23624 24840 24041 24868
rect 23624 24828 23630 24840
rect 24029 24837 24041 24840
rect 24075 24837 24087 24871
rect 24946 24868 24952 24880
rect 24907 24840 24952 24868
rect 24029 24831 24087 24837
rect 24946 24828 24952 24840
rect 25004 24828 25010 24880
rect 27264 24840 27476 24868
rect 19613 24803 19671 24809
rect 19613 24800 19625 24803
rect 19076 24772 19625 24800
rect 18969 24763 19027 24769
rect 19613 24769 19625 24772
rect 19659 24769 19671 24803
rect 21634 24800 21640 24812
rect 19613 24763 19671 24769
rect 21376 24772 21640 24800
rect 15010 24732 15016 24744
rect 14971 24704 15016 24732
rect 15010 24692 15016 24704
rect 15068 24692 15074 24744
rect 16942 24692 16948 24744
rect 17000 24732 17006 24744
rect 17589 24735 17647 24741
rect 17589 24732 17601 24735
rect 17000 24704 17601 24732
rect 17000 24692 17006 24704
rect 17589 24701 17601 24704
rect 17635 24701 17647 24735
rect 17589 24695 17647 24701
rect 17678 24692 17684 24744
rect 17736 24732 17742 24744
rect 18984 24732 19012 24763
rect 17736 24704 19012 24732
rect 19061 24735 19119 24741
rect 17736 24692 17742 24704
rect 19061 24701 19073 24735
rect 19107 24732 19119 24735
rect 19334 24732 19340 24744
rect 19107 24704 19340 24732
rect 19107 24701 19119 24704
rect 19061 24695 19119 24701
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 20349 24735 20407 24741
rect 20349 24701 20361 24735
rect 20395 24732 20407 24735
rect 20438 24732 20444 24744
rect 20395 24704 20444 24732
rect 20395 24701 20407 24704
rect 20349 24695 20407 24701
rect 20438 24692 20444 24704
rect 20496 24692 20502 24744
rect 21174 24732 21180 24744
rect 21135 24704 21180 24732
rect 21174 24692 21180 24704
rect 21232 24732 21238 24744
rect 21376 24732 21404 24772
rect 21634 24760 21640 24772
rect 21692 24760 21698 24812
rect 22186 24800 22192 24812
rect 22147 24772 22192 24800
rect 22186 24760 22192 24772
rect 22244 24760 22250 24812
rect 22554 24760 22560 24812
rect 22612 24800 22618 24812
rect 22649 24803 22707 24809
rect 22649 24800 22661 24803
rect 22612 24772 22661 24800
rect 22612 24760 22618 24772
rect 22649 24769 22661 24772
rect 22695 24800 22707 24803
rect 23474 24800 23480 24812
rect 22695 24772 23480 24800
rect 22695 24769 22707 24772
rect 22649 24763 22707 24769
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 25501 24803 25559 24809
rect 25501 24769 25513 24803
rect 25547 24800 25559 24803
rect 25590 24800 25596 24812
rect 25547 24772 25596 24800
rect 25547 24769 25559 24772
rect 25501 24763 25559 24769
rect 25590 24760 25596 24772
rect 25648 24760 25654 24812
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24800 25743 24803
rect 27154 24800 27160 24812
rect 25731 24772 27160 24800
rect 25731 24769 25743 24772
rect 25685 24763 25743 24769
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 22462 24732 22468 24744
rect 21232 24704 21404 24732
rect 21468 24704 22468 24732
rect 21232 24692 21238 24704
rect 19705 24667 19763 24673
rect 14660 24636 17632 24664
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 2682 24596 2688 24608
rect 1627 24568 2688 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 6822 24556 6828 24608
rect 6880 24596 6886 24608
rect 17494 24596 17500 24608
rect 6880 24568 17500 24596
rect 6880 24556 6886 24568
rect 17494 24556 17500 24568
rect 17552 24556 17558 24608
rect 17604 24596 17632 24636
rect 18248 24636 19656 24664
rect 18248 24596 18276 24636
rect 18414 24596 18420 24608
rect 17604 24568 18276 24596
rect 18375 24568 18420 24596
rect 18414 24556 18420 24568
rect 18472 24556 18478 24608
rect 19628 24596 19656 24636
rect 19705 24633 19717 24667
rect 19751 24664 19763 24667
rect 21468 24664 21496 24704
rect 22462 24692 22468 24704
rect 22520 24692 22526 24744
rect 23382 24692 23388 24744
rect 23440 24732 23446 24744
rect 23937 24735 23995 24741
rect 23937 24732 23949 24735
rect 23440 24704 23949 24732
rect 23440 24692 23446 24704
rect 23937 24701 23949 24704
rect 23983 24701 23995 24735
rect 23937 24695 23995 24701
rect 22741 24667 22799 24673
rect 22741 24664 22753 24667
rect 19751 24636 21496 24664
rect 21560 24636 22753 24664
rect 19751 24633 19763 24636
rect 19705 24627 19763 24633
rect 21560 24596 21588 24636
rect 22741 24633 22753 24636
rect 22787 24633 22799 24667
rect 22741 24627 22799 24633
rect 22830 24624 22836 24676
rect 22888 24664 22894 24676
rect 27264 24664 27292 24840
rect 27341 24803 27399 24809
rect 27341 24769 27353 24803
rect 27387 24769 27399 24803
rect 27448 24800 27476 24840
rect 27985 24803 28043 24809
rect 27985 24800 27997 24803
rect 27448 24772 27997 24800
rect 27341 24763 27399 24769
rect 27985 24769 27997 24772
rect 28031 24769 28043 24803
rect 27985 24763 28043 24769
rect 28997 24803 29055 24809
rect 28997 24769 29009 24803
rect 29043 24800 29055 24803
rect 37826 24800 37832 24812
rect 29043 24772 37832 24800
rect 29043 24769 29055 24772
rect 28997 24763 29055 24769
rect 27356 24732 27384 24763
rect 37826 24760 37832 24772
rect 37884 24760 37890 24812
rect 38010 24800 38016 24812
rect 37971 24772 38016 24800
rect 38010 24760 38016 24772
rect 38068 24760 38074 24812
rect 29270 24732 29276 24744
rect 27356 24704 29276 24732
rect 29270 24692 29276 24704
rect 29328 24692 29334 24744
rect 22888 24636 27292 24664
rect 22888 24624 22894 24636
rect 19628 24568 21588 24596
rect 22005 24599 22063 24605
rect 22005 24565 22017 24599
rect 22051 24596 22063 24599
rect 22094 24596 22100 24608
rect 22051 24568 22100 24596
rect 22051 24565 22063 24568
rect 22005 24559 22063 24565
rect 22094 24556 22100 24568
rect 22152 24556 22158 24608
rect 25498 24556 25504 24608
rect 25556 24596 25562 24608
rect 25869 24599 25927 24605
rect 25869 24596 25881 24599
rect 25556 24568 25881 24596
rect 25556 24556 25562 24568
rect 25869 24565 25881 24568
rect 25915 24565 25927 24599
rect 27154 24596 27160 24608
rect 27115 24568 27160 24596
rect 25869 24559 25927 24565
rect 27154 24556 27160 24568
rect 27212 24556 27218 24608
rect 28077 24599 28135 24605
rect 28077 24565 28089 24599
rect 28123 24596 28135 24599
rect 28350 24596 28356 24608
rect 28123 24568 28356 24596
rect 28123 24565 28135 24568
rect 28077 24559 28135 24565
rect 28350 24556 28356 24568
rect 28408 24556 28414 24608
rect 29086 24596 29092 24608
rect 29047 24568 29092 24596
rect 29086 24556 29092 24568
rect 29144 24556 29150 24608
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 6822 24392 6828 24404
rect 2746 24364 6408 24392
rect 6783 24364 6828 24392
rect 2225 24327 2283 24333
rect 2225 24293 2237 24327
rect 2271 24324 2283 24327
rect 2746 24324 2774 24364
rect 2271 24296 2774 24324
rect 6380 24324 6408 24364
rect 6822 24352 6828 24364
rect 6880 24352 6886 24404
rect 6914 24352 6920 24404
rect 6972 24392 6978 24404
rect 9398 24392 9404 24404
rect 6972 24364 9404 24392
rect 6972 24352 6978 24364
rect 9398 24352 9404 24364
rect 9456 24392 9462 24404
rect 22186 24392 22192 24404
rect 9456 24364 22192 24392
rect 9456 24352 9462 24364
rect 22186 24352 22192 24364
rect 22244 24352 22250 24404
rect 23032 24364 23888 24392
rect 18690 24324 18696 24336
rect 6380 24296 12434 24324
rect 2271 24293 2283 24296
rect 2225 24287 2283 24293
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24188 1639 24191
rect 2240 24188 2268 24287
rect 3602 24216 3608 24268
rect 3660 24256 3666 24268
rect 5077 24259 5135 24265
rect 5077 24256 5089 24259
rect 3660 24228 5089 24256
rect 3660 24216 3666 24228
rect 5077 24225 5089 24228
rect 5123 24225 5135 24259
rect 5350 24256 5356 24268
rect 5311 24228 5356 24256
rect 5077 24219 5135 24225
rect 5350 24216 5356 24228
rect 5408 24216 5414 24268
rect 7466 24216 7472 24268
rect 7524 24256 7530 24268
rect 9861 24259 9919 24265
rect 9861 24256 9873 24259
rect 7524 24228 9873 24256
rect 7524 24216 7530 24228
rect 9861 24225 9873 24228
rect 9907 24225 9919 24259
rect 9861 24219 9919 24225
rect 12161 24259 12219 24265
rect 12161 24225 12173 24259
rect 12207 24256 12219 24259
rect 12250 24256 12256 24268
rect 12207 24228 12256 24256
rect 12207 24225 12219 24228
rect 12161 24219 12219 24225
rect 12250 24216 12256 24228
rect 12308 24216 12314 24268
rect 1627 24160 2268 24188
rect 4433 24191 4491 24197
rect 1627 24157 1639 24160
rect 1581 24151 1639 24157
rect 4433 24157 4445 24191
rect 4479 24188 4491 24191
rect 4706 24188 4712 24200
rect 4479 24160 4712 24188
rect 4479 24157 4491 24160
rect 4433 24151 4491 24157
rect 4706 24148 4712 24160
rect 4764 24148 4770 24200
rect 3326 24080 3332 24132
rect 3384 24120 3390 24132
rect 3384 24092 5842 24120
rect 3384 24080 3390 24092
rect 6730 24080 6736 24132
rect 6788 24120 6794 24132
rect 9125 24123 9183 24129
rect 9125 24120 9137 24123
rect 6788 24092 9137 24120
rect 6788 24080 6794 24092
rect 9125 24089 9137 24092
rect 9171 24120 9183 24123
rect 11333 24123 11391 24129
rect 11333 24120 11345 24123
rect 9171 24092 11345 24120
rect 9171 24089 9183 24092
rect 9125 24083 9183 24089
rect 11333 24089 11345 24092
rect 11379 24120 11391 24123
rect 11514 24120 11520 24132
rect 11379 24092 11520 24120
rect 11379 24089 11391 24092
rect 11333 24083 11391 24089
rect 11514 24080 11520 24092
rect 11572 24120 11578 24132
rect 11882 24120 11888 24132
rect 11572 24092 11888 24120
rect 11572 24080 11578 24092
rect 11882 24080 11888 24092
rect 11940 24080 11946 24132
rect 12268 24120 12296 24216
rect 12406 24188 12434 24296
rect 17972 24296 18696 24324
rect 14274 24216 14280 24268
rect 14332 24256 14338 24268
rect 16485 24259 16543 24265
rect 16485 24256 16497 24259
rect 14332 24228 16497 24256
rect 14332 24216 14338 24228
rect 16485 24225 16497 24228
rect 16531 24256 16543 24259
rect 16850 24256 16856 24268
rect 16531 24228 16856 24256
rect 16531 24225 16543 24228
rect 16485 24219 16543 24225
rect 16850 24216 16856 24228
rect 16908 24216 16914 24268
rect 17972 24188 18000 24296
rect 18690 24284 18696 24296
rect 18748 24284 18754 24336
rect 19242 24284 19248 24336
rect 19300 24324 19306 24336
rect 20073 24327 20131 24333
rect 20073 24324 20085 24327
rect 19300 24296 20085 24324
rect 19300 24284 19306 24296
rect 20073 24293 20085 24296
rect 20119 24293 20131 24327
rect 20073 24287 20131 24293
rect 21913 24327 21971 24333
rect 21913 24293 21925 24327
rect 21959 24324 21971 24327
rect 22830 24324 22836 24336
rect 21959 24296 22836 24324
rect 21959 24293 21971 24296
rect 21913 24287 21971 24293
rect 22830 24284 22836 24296
rect 22888 24284 22894 24336
rect 23032 24256 23060 24364
rect 23106 24284 23112 24336
rect 23164 24324 23170 24336
rect 23860 24324 23888 24364
rect 25590 24352 25596 24404
rect 25648 24392 25654 24404
rect 26237 24395 26295 24401
rect 26237 24392 26249 24395
rect 25648 24364 26249 24392
rect 25648 24352 25654 24364
rect 26237 24361 26249 24364
rect 26283 24361 26295 24395
rect 32490 24392 32496 24404
rect 26237 24355 26295 24361
rect 26344 24364 32496 24392
rect 26344 24324 26372 24364
rect 32490 24352 32496 24364
rect 32548 24352 32554 24404
rect 37826 24352 37832 24404
rect 37884 24392 37890 24404
rect 38105 24395 38163 24401
rect 38105 24392 38117 24395
rect 37884 24364 38117 24392
rect 37884 24352 37890 24364
rect 38105 24361 38117 24364
rect 38151 24361 38163 24395
rect 38105 24355 38163 24361
rect 23164 24296 23796 24324
rect 23860 24296 26372 24324
rect 23164 24284 23170 24296
rect 12406 24160 15332 24188
rect 17894 24160 18000 24188
rect 18064 24228 23060 24256
rect 13262 24120 13268 24132
rect 12268 24092 13268 24120
rect 13262 24080 13268 24092
rect 13320 24080 13326 24132
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 4525 24055 4583 24061
rect 4525 24021 4537 24055
rect 4571 24052 4583 24055
rect 8110 24052 8116 24064
rect 4571 24024 8116 24052
rect 4571 24021 4583 24024
rect 4525 24015 4583 24021
rect 8110 24012 8116 24024
rect 8168 24012 8174 24064
rect 11900 24052 11928 24080
rect 15194 24052 15200 24064
rect 11900 24024 15200 24052
rect 15194 24012 15200 24024
rect 15252 24012 15258 24064
rect 15304 24052 15332 24160
rect 16758 24120 16764 24132
rect 16719 24092 16764 24120
rect 16758 24080 16764 24092
rect 16816 24080 16822 24132
rect 18064 24052 18092 24228
rect 18690 24188 18696 24200
rect 18651 24160 18696 24188
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 19242 24148 19248 24200
rect 19300 24188 19306 24200
rect 19981 24191 20039 24197
rect 19981 24188 19993 24191
rect 19300 24160 19993 24188
rect 19300 24148 19306 24160
rect 19981 24157 19993 24160
rect 20027 24188 20039 24191
rect 20346 24188 20352 24200
rect 20027 24160 20352 24188
rect 20027 24157 20039 24160
rect 19981 24151 20039 24157
rect 20346 24148 20352 24160
rect 20404 24148 20410 24200
rect 21361 24191 21419 24197
rect 21361 24157 21373 24191
rect 21407 24188 21419 24191
rect 21450 24188 21456 24200
rect 21407 24160 21456 24188
rect 21407 24157 21419 24160
rect 21361 24151 21419 24157
rect 21450 24148 21456 24160
rect 21508 24148 21514 24200
rect 21818 24188 21824 24200
rect 21779 24160 21824 24188
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 21910 24148 21916 24200
rect 21968 24188 21974 24200
rect 22554 24188 22560 24200
rect 21968 24160 22560 24188
rect 21968 24148 21974 24160
rect 22554 24148 22560 24160
rect 22612 24148 22618 24200
rect 22649 24191 22707 24197
rect 22649 24157 22661 24191
rect 22695 24157 22707 24191
rect 23106 24188 23112 24200
rect 23067 24160 23112 24188
rect 22649 24151 22707 24157
rect 19150 24120 19156 24132
rect 18248 24092 19156 24120
rect 15304 24024 18092 24052
rect 18138 24012 18144 24064
rect 18196 24052 18202 24064
rect 18248 24061 18276 24092
rect 19150 24080 19156 24092
rect 19208 24080 19214 24132
rect 20714 24120 20720 24132
rect 20675 24092 20720 24120
rect 20714 24080 20720 24092
rect 20772 24080 20778 24132
rect 20809 24123 20867 24129
rect 20809 24089 20821 24123
rect 20855 24089 20867 24123
rect 20809 24083 20867 24089
rect 21468 24092 22094 24120
rect 18233 24055 18291 24061
rect 18233 24052 18245 24055
rect 18196 24024 18245 24052
rect 18196 24012 18202 24024
rect 18233 24021 18245 24024
rect 18279 24021 18291 24055
rect 18782 24052 18788 24064
rect 18743 24024 18788 24052
rect 18233 24015 18291 24021
rect 18782 24012 18788 24024
rect 18840 24012 18846 24064
rect 18874 24012 18880 24064
rect 18932 24052 18938 24064
rect 20622 24052 20628 24064
rect 18932 24024 20628 24052
rect 18932 24012 18938 24024
rect 20622 24012 20628 24024
rect 20680 24012 20686 24064
rect 20824 24052 20852 24083
rect 21468 24052 21496 24092
rect 20824 24024 21496 24052
rect 22066 24052 22094 24092
rect 22186 24080 22192 24132
rect 22244 24120 22250 24132
rect 22664 24120 22692 24151
rect 23106 24148 23112 24160
rect 23164 24148 23170 24200
rect 23768 24197 23796 24296
rect 27154 24284 27160 24336
rect 27212 24324 27218 24336
rect 38010 24324 38016 24336
rect 27212 24296 38016 24324
rect 27212 24284 27218 24296
rect 38010 24284 38016 24296
rect 38068 24284 38074 24336
rect 24946 24216 24952 24268
rect 25004 24256 25010 24268
rect 26878 24256 26884 24268
rect 25004 24228 26884 24256
rect 25004 24216 25010 24228
rect 26878 24216 26884 24228
rect 26936 24216 26942 24268
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24157 23811 24191
rect 26142 24188 26148 24200
rect 26103 24160 26148 24188
rect 23753 24151 23811 24157
rect 26142 24148 26148 24160
rect 26200 24148 26206 24200
rect 26789 24191 26847 24197
rect 26789 24188 26801 24191
rect 26252 24160 26801 24188
rect 22244 24092 22692 24120
rect 24673 24123 24731 24129
rect 22244 24080 22250 24092
rect 24673 24089 24685 24123
rect 24719 24089 24731 24123
rect 24673 24083 24731 24089
rect 24765 24123 24823 24129
rect 24765 24089 24777 24123
rect 24811 24120 24823 24123
rect 24854 24120 24860 24132
rect 24811 24092 24860 24120
rect 24811 24089 24823 24092
rect 24765 24083 24823 24089
rect 22465 24055 22523 24061
rect 22465 24052 22477 24055
rect 22066 24024 22477 24052
rect 22465 24021 22477 24024
rect 22511 24021 22523 24055
rect 22465 24015 22523 24021
rect 22738 24012 22744 24064
rect 22796 24052 22802 24064
rect 23201 24055 23259 24061
rect 23201 24052 23213 24055
rect 22796 24024 23213 24052
rect 22796 24012 22802 24024
rect 23201 24021 23213 24024
rect 23247 24021 23259 24055
rect 23201 24015 23259 24021
rect 23290 24012 23296 24064
rect 23348 24052 23354 24064
rect 23845 24055 23903 24061
rect 23845 24052 23857 24055
rect 23348 24024 23857 24052
rect 23348 24012 23354 24024
rect 23845 24021 23857 24024
rect 23891 24021 23903 24055
rect 24688 24052 24716 24083
rect 24854 24080 24860 24092
rect 24912 24080 24918 24132
rect 25682 24120 25688 24132
rect 25643 24092 25688 24120
rect 25682 24080 25688 24092
rect 25740 24080 25746 24132
rect 25498 24052 25504 24064
rect 24688 24024 25504 24052
rect 23845 24015 23903 24021
rect 25498 24012 25504 24024
rect 25556 24012 25562 24064
rect 25590 24012 25596 24064
rect 25648 24052 25654 24064
rect 26252 24052 26280 24160
rect 26789 24157 26801 24160
rect 26835 24157 26847 24191
rect 38286 24188 38292 24200
rect 38247 24160 38292 24188
rect 26789 24151 26847 24157
rect 38286 24148 38292 24160
rect 38344 24148 38350 24200
rect 26878 24052 26884 24064
rect 25648 24024 26280 24052
rect 26839 24024 26884 24052
rect 25648 24012 25654 24024
rect 26878 24012 26884 24024
rect 26936 24012 26942 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1857 23851 1915 23857
rect 1857 23817 1869 23851
rect 1903 23848 1915 23851
rect 4614 23848 4620 23860
rect 1903 23820 4620 23848
rect 1903 23817 1915 23820
rect 1857 23811 1915 23817
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 5534 23848 5540 23860
rect 4764 23820 5540 23848
rect 4764 23808 4770 23820
rect 5534 23808 5540 23820
rect 5592 23848 5598 23860
rect 5718 23848 5724 23860
rect 5592 23820 5724 23848
rect 5592 23808 5598 23820
rect 5718 23808 5724 23820
rect 5776 23808 5782 23860
rect 9214 23848 9220 23860
rect 9175 23820 9220 23848
rect 9214 23808 9220 23820
rect 9272 23808 9278 23860
rect 13906 23848 13912 23860
rect 12268 23820 13912 23848
rect 2774 23780 2780 23792
rect 1780 23752 2780 23780
rect 1780 23721 1808 23752
rect 2774 23740 2780 23752
rect 2832 23740 2838 23792
rect 3694 23740 3700 23792
rect 3752 23740 3758 23792
rect 5353 23783 5411 23789
rect 5353 23749 5365 23783
rect 5399 23780 5411 23783
rect 5399 23752 8234 23780
rect 5399 23749 5411 23752
rect 5353 23743 5411 23749
rect 1765 23715 1823 23721
rect 1765 23681 1777 23715
rect 1811 23681 1823 23715
rect 5258 23712 5264 23724
rect 5219 23684 5264 23712
rect 1765 23675 1823 23681
rect 5258 23672 5264 23684
rect 5316 23672 5322 23724
rect 5718 23672 5724 23724
rect 5776 23712 5782 23724
rect 6546 23712 6552 23724
rect 5776 23684 6552 23712
rect 5776 23672 5782 23684
rect 6546 23672 6552 23684
rect 6604 23672 6610 23724
rect 7466 23712 7472 23724
rect 7427 23684 7472 23712
rect 7466 23672 7472 23684
rect 7524 23672 7530 23724
rect 12066 23672 12072 23724
rect 12124 23712 12130 23724
rect 12268 23721 12296 23820
rect 13906 23808 13912 23820
rect 13964 23808 13970 23860
rect 14366 23808 14372 23860
rect 14424 23848 14430 23860
rect 15010 23848 15016 23860
rect 14424 23820 15016 23848
rect 14424 23808 14430 23820
rect 15010 23808 15016 23820
rect 15068 23808 15074 23860
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 18601 23851 18659 23857
rect 18601 23848 18613 23851
rect 16816 23820 18613 23848
rect 16816 23808 16822 23820
rect 18601 23817 18613 23820
rect 18647 23848 18659 23851
rect 21818 23848 21824 23860
rect 18647 23820 21824 23848
rect 18647 23817 18659 23820
rect 18601 23811 18659 23817
rect 21818 23808 21824 23820
rect 21876 23808 21882 23860
rect 25498 23848 25504 23860
rect 25459 23820 25504 23848
rect 25498 23808 25504 23820
rect 25556 23808 25562 23860
rect 26142 23808 26148 23860
rect 26200 23848 26206 23860
rect 28994 23848 29000 23860
rect 26200 23820 29000 23848
rect 26200 23808 26206 23820
rect 28994 23808 29000 23820
rect 29052 23808 29058 23860
rect 18414 23780 18420 23792
rect 12406 23752 14030 23780
rect 18354 23752 18420 23780
rect 12253 23715 12311 23721
rect 12253 23712 12265 23715
rect 12124 23684 12265 23712
rect 12124 23672 12130 23684
rect 12253 23681 12265 23684
rect 12299 23681 12311 23715
rect 12253 23675 12311 23681
rect 2406 23644 2412 23656
rect 2367 23616 2412 23644
rect 2406 23604 2412 23616
rect 2464 23604 2470 23656
rect 2685 23647 2743 23653
rect 2685 23613 2697 23647
rect 2731 23644 2743 23647
rect 4890 23644 4896 23656
rect 2731 23616 4896 23644
rect 2731 23613 2743 23616
rect 2685 23607 2743 23613
rect 4890 23604 4896 23616
rect 4948 23644 4954 23656
rect 5074 23644 5080 23656
rect 4948 23616 5080 23644
rect 4948 23604 4954 23616
rect 5074 23604 5080 23616
rect 5132 23604 5138 23656
rect 7282 23604 7288 23656
rect 7340 23644 7346 23656
rect 7742 23644 7748 23656
rect 7340 23616 7748 23644
rect 7340 23604 7346 23616
rect 7742 23604 7748 23616
rect 7800 23604 7806 23656
rect 11238 23604 11244 23656
rect 11296 23644 11302 23656
rect 12406 23644 12434 23752
rect 18414 23740 18420 23752
rect 18472 23740 18478 23792
rect 19978 23740 19984 23792
rect 20036 23780 20042 23792
rect 20533 23783 20591 23789
rect 20533 23780 20545 23783
rect 20036 23752 20545 23780
rect 20036 23740 20042 23752
rect 20533 23749 20545 23752
rect 20579 23749 20591 23783
rect 22554 23780 22560 23792
rect 22515 23752 22560 23780
rect 20533 23743 20591 23749
rect 22554 23740 22560 23752
rect 22612 23740 22618 23792
rect 26878 23780 26884 23792
rect 25056 23752 26884 23780
rect 16850 23712 16856 23724
rect 16811 23684 16856 23712
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 23937 23715 23995 23721
rect 23937 23681 23949 23715
rect 23983 23712 23995 23715
rect 24670 23712 24676 23724
rect 23983 23684 24676 23712
rect 23983 23681 23995 23684
rect 23937 23675 23995 23681
rect 24670 23672 24676 23684
rect 24728 23672 24734 23724
rect 25056 23721 25084 23752
rect 26878 23740 26884 23752
rect 26936 23740 26942 23792
rect 25041 23715 25099 23721
rect 25041 23681 25053 23715
rect 25087 23681 25099 23715
rect 25041 23675 25099 23681
rect 25774 23672 25780 23724
rect 25832 23712 25838 23724
rect 25961 23715 26019 23721
rect 25961 23712 25973 23715
rect 25832 23684 25973 23712
rect 25832 23672 25838 23684
rect 25961 23681 25973 23684
rect 26007 23681 26019 23715
rect 25961 23675 26019 23681
rect 13262 23644 13268 23656
rect 11296 23616 12434 23644
rect 13223 23616 13268 23644
rect 11296 23604 11302 23616
rect 13262 23604 13268 23616
rect 13320 23604 13326 23656
rect 13538 23644 13544 23656
rect 13499 23616 13544 23644
rect 13538 23604 13544 23616
rect 13596 23604 13602 23656
rect 17129 23647 17187 23653
rect 17129 23613 17141 23647
rect 17175 23644 17187 23647
rect 18598 23644 18604 23656
rect 17175 23616 18604 23644
rect 17175 23613 17187 23616
rect 17129 23607 17187 23613
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 19426 23604 19432 23656
rect 19484 23644 19490 23656
rect 19978 23644 19984 23656
rect 19484 23616 19984 23644
rect 19484 23604 19490 23616
rect 19978 23604 19984 23616
rect 20036 23604 20042 23656
rect 20438 23653 20444 23656
rect 20430 23647 20444 23653
rect 20430 23644 20442 23647
rect 20351 23616 20442 23644
rect 20430 23613 20442 23616
rect 20496 23644 20502 23656
rect 21453 23647 21511 23653
rect 20496 23616 21404 23644
rect 20430 23607 20444 23613
rect 20438 23604 20444 23607
rect 20496 23604 20502 23616
rect 4157 23579 4215 23585
rect 4157 23545 4169 23579
rect 4203 23576 4215 23579
rect 4614 23576 4620 23588
rect 4203 23548 4620 23576
rect 4203 23545 4215 23548
rect 4157 23539 4215 23545
rect 4614 23536 4620 23548
rect 4672 23576 4678 23588
rect 21376 23576 21404 23616
rect 21453 23613 21465 23647
rect 21499 23644 21511 23647
rect 21634 23644 21640 23656
rect 21499 23616 21640 23644
rect 21499 23613 21511 23616
rect 21453 23607 21511 23613
rect 21634 23604 21640 23616
rect 21692 23604 21698 23656
rect 22462 23644 22468 23656
rect 22423 23616 22468 23644
rect 22462 23604 22468 23616
rect 22520 23604 22526 23656
rect 22922 23644 22928 23656
rect 22883 23616 22928 23644
rect 22922 23604 22928 23616
rect 22980 23604 22986 23656
rect 24857 23647 24915 23653
rect 24857 23613 24869 23647
rect 24903 23644 24915 23647
rect 29086 23644 29092 23656
rect 24903 23616 29092 23644
rect 24903 23613 24915 23616
rect 24857 23607 24915 23613
rect 29086 23604 29092 23616
rect 29144 23604 29150 23656
rect 31110 23604 31116 23656
rect 31168 23644 31174 23656
rect 31205 23647 31263 23653
rect 31205 23644 31217 23647
rect 31168 23616 31217 23644
rect 31168 23604 31174 23616
rect 31205 23613 31217 23616
rect 31251 23613 31263 23647
rect 31205 23607 31263 23613
rect 26970 23576 26976 23588
rect 4672 23548 6776 23576
rect 21376 23548 26976 23576
rect 4672 23536 4678 23548
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 5258 23508 5264 23520
rect 2832 23480 5264 23508
rect 2832 23468 2838 23480
rect 5258 23468 5264 23480
rect 5316 23468 5322 23520
rect 5350 23468 5356 23520
rect 5408 23508 5414 23520
rect 6641 23511 6699 23517
rect 6641 23508 6653 23511
rect 5408 23480 6653 23508
rect 5408 23468 5414 23480
rect 6641 23477 6653 23480
rect 6687 23477 6699 23511
rect 6748 23508 6776 23548
rect 26970 23536 26976 23548
rect 27028 23536 27034 23588
rect 9122 23508 9128 23520
rect 6748 23480 9128 23508
rect 6641 23471 6699 23477
rect 9122 23468 9128 23480
rect 9180 23468 9186 23520
rect 12345 23511 12403 23517
rect 12345 23477 12357 23511
rect 12391 23508 12403 23511
rect 13722 23508 13728 23520
rect 12391 23480 13728 23508
rect 12391 23477 12403 23480
rect 12345 23471 12403 23477
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 13906 23468 13912 23520
rect 13964 23508 13970 23520
rect 16850 23508 16856 23520
rect 13964 23480 16856 23508
rect 13964 23468 13970 23480
rect 16850 23468 16856 23480
rect 16908 23468 16914 23520
rect 19150 23468 19156 23520
rect 19208 23508 19214 23520
rect 20622 23508 20628 23520
rect 19208 23480 20628 23508
rect 19208 23468 19214 23480
rect 20622 23468 20628 23480
rect 20680 23468 20686 23520
rect 20714 23468 20720 23520
rect 20772 23508 20778 23520
rect 23382 23508 23388 23520
rect 20772 23480 23388 23508
rect 20772 23468 20778 23480
rect 23382 23468 23388 23480
rect 23440 23468 23446 23520
rect 23750 23468 23756 23520
rect 23808 23508 23814 23520
rect 24029 23511 24087 23517
rect 24029 23508 24041 23511
rect 23808 23480 24041 23508
rect 23808 23468 23814 23480
rect 24029 23477 24041 23480
rect 24075 23477 24087 23511
rect 24029 23471 24087 23477
rect 25958 23468 25964 23520
rect 26016 23508 26022 23520
rect 26053 23511 26111 23517
rect 26053 23508 26065 23511
rect 26016 23480 26065 23508
rect 26016 23468 26022 23480
rect 26053 23477 26065 23480
rect 26099 23477 26111 23511
rect 26053 23471 26111 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 5258 23264 5264 23316
rect 5316 23304 5322 23316
rect 20530 23304 20536 23316
rect 5316 23276 12434 23304
rect 5316 23264 5322 23276
rect 3970 23128 3976 23180
rect 4028 23168 4034 23180
rect 6641 23171 6699 23177
rect 6641 23168 6653 23171
rect 4028 23140 6653 23168
rect 4028 23128 4034 23140
rect 6641 23137 6653 23140
rect 6687 23137 6699 23171
rect 6641 23131 6699 23137
rect 10413 23171 10471 23177
rect 10413 23137 10425 23171
rect 10459 23168 10471 23171
rect 12250 23168 12256 23180
rect 10459 23140 12256 23168
rect 10459 23137 10471 23140
rect 10413 23131 10471 23137
rect 12250 23128 12256 23140
rect 12308 23128 12314 23180
rect 1857 23103 1915 23109
rect 1857 23069 1869 23103
rect 1903 23100 1915 23103
rect 1946 23100 1952 23112
rect 1903 23072 1952 23100
rect 1903 23069 1915 23072
rect 1857 23063 1915 23069
rect 1946 23060 1952 23072
rect 2004 23060 2010 23112
rect 5261 23103 5319 23109
rect 5261 23069 5273 23103
rect 5307 23100 5319 23103
rect 5534 23100 5540 23112
rect 5307 23072 5540 23100
rect 5307 23069 5319 23072
rect 5261 23063 5319 23069
rect 5534 23060 5540 23072
rect 5592 23060 5598 23112
rect 5626 23060 5632 23112
rect 5684 23100 5690 23112
rect 5905 23103 5963 23109
rect 5905 23100 5917 23103
rect 5684 23072 5917 23100
rect 5684 23060 5690 23072
rect 5905 23069 5917 23072
rect 5951 23100 5963 23103
rect 6730 23100 6736 23112
rect 5951 23072 6736 23100
rect 5951 23069 5963 23072
rect 5905 23063 5963 23069
rect 6730 23060 6736 23072
rect 6788 23060 6794 23112
rect 7285 23103 7343 23109
rect 7285 23069 7297 23103
rect 7331 23100 7343 23103
rect 9582 23100 9588 23112
rect 7331 23072 9588 23100
rect 7331 23069 7343 23072
rect 7285 23063 7343 23069
rect 9582 23060 9588 23072
rect 9640 23060 9646 23112
rect 12406 23100 12434 23276
rect 13464 23276 20536 23304
rect 13081 23103 13139 23109
rect 13081 23100 13093 23103
rect 12406 23072 13093 23100
rect 13081 23069 13093 23072
rect 13127 23100 13139 23103
rect 13464 23100 13492 23276
rect 20530 23264 20536 23276
rect 20588 23264 20594 23316
rect 21545 23307 21603 23313
rect 21545 23273 21557 23307
rect 21591 23304 21603 23307
rect 24762 23304 24768 23316
rect 21591 23276 24768 23304
rect 21591 23273 21603 23276
rect 21545 23267 21603 23273
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 26970 23264 26976 23316
rect 27028 23304 27034 23316
rect 27246 23304 27252 23316
rect 27028 23276 27252 23304
rect 27028 23264 27034 23276
rect 27246 23264 27252 23276
rect 27304 23264 27310 23316
rect 29822 23304 29828 23316
rect 29783 23276 29828 23304
rect 29822 23264 29828 23276
rect 29880 23264 29886 23316
rect 17218 23196 17224 23248
rect 17276 23236 17282 23248
rect 22094 23236 22100 23248
rect 17276 23208 22100 23236
rect 17276 23196 17282 23208
rect 22094 23196 22100 23208
rect 22152 23236 22158 23248
rect 22278 23236 22284 23248
rect 22152 23208 22284 23236
rect 22152 23196 22158 23208
rect 22278 23196 22284 23208
rect 22336 23196 22342 23248
rect 25130 23196 25136 23248
rect 25188 23236 25194 23248
rect 25225 23239 25283 23245
rect 25225 23236 25237 23239
rect 25188 23208 25237 23236
rect 25188 23196 25194 23208
rect 25225 23205 25237 23208
rect 25271 23205 25283 23239
rect 25225 23199 25283 23205
rect 25682 23196 25688 23248
rect 25740 23236 25746 23248
rect 30834 23236 30840 23248
rect 25740 23208 30840 23236
rect 25740 23196 25746 23208
rect 30834 23196 30840 23208
rect 30892 23196 30898 23248
rect 14553 23171 14611 23177
rect 14553 23137 14565 23171
rect 14599 23168 14611 23171
rect 16482 23168 16488 23180
rect 14599 23140 16488 23168
rect 14599 23137 14611 23140
rect 14553 23131 14611 23137
rect 16482 23128 16488 23140
rect 16540 23128 16546 23180
rect 16850 23128 16856 23180
rect 16908 23168 16914 23180
rect 18693 23171 18751 23177
rect 18693 23168 18705 23171
rect 16908 23140 18705 23168
rect 16908 23128 16914 23140
rect 18693 23137 18705 23140
rect 18739 23168 18751 23171
rect 19242 23168 19248 23180
rect 18739 23140 19248 23168
rect 18739 23137 18751 23140
rect 18693 23131 18751 23137
rect 19242 23128 19248 23140
rect 19300 23128 19306 23180
rect 20530 23168 20536 23180
rect 20491 23140 20536 23168
rect 20530 23128 20536 23140
rect 20588 23128 20594 23180
rect 20990 23128 20996 23180
rect 21048 23168 21054 23180
rect 21910 23168 21916 23180
rect 21048 23140 21916 23168
rect 21048 23128 21054 23140
rect 21910 23128 21916 23140
rect 21968 23128 21974 23180
rect 31110 23168 31116 23180
rect 22066 23140 25820 23168
rect 31071 23140 31116 23168
rect 14274 23100 14280 23112
rect 13127 23072 13492 23100
rect 13556 23072 14280 23100
rect 13127 23069 13139 23072
rect 13081 23063 13139 23069
rect 9490 22992 9496 23044
rect 9548 23032 9554 23044
rect 10689 23035 10747 23041
rect 10689 23032 10701 23035
rect 9548 23004 10701 23032
rect 9548 22992 9554 23004
rect 10689 23001 10701 23004
rect 10735 23032 10747 23035
rect 10778 23032 10784 23044
rect 10735 23004 10784 23032
rect 10735 23001 10747 23004
rect 10689 22995 10747 23001
rect 10778 22992 10784 23004
rect 10836 22992 10842 23044
rect 11698 22992 11704 23044
rect 11756 22992 11762 23044
rect 12250 22992 12256 23044
rect 12308 23032 12314 23044
rect 13556 23032 13584 23072
rect 14274 23060 14280 23072
rect 14332 23060 14338 23112
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23100 18015 23103
rect 18506 23100 18512 23112
rect 18003 23072 18512 23100
rect 18003 23069 18015 23072
rect 17957 23063 18015 23069
rect 18506 23060 18512 23072
rect 18564 23100 18570 23112
rect 18966 23100 18972 23112
rect 18564 23072 18972 23100
rect 18564 23060 18570 23072
rect 18966 23060 18972 23072
rect 19024 23100 19030 23112
rect 20073 23103 20131 23109
rect 20073 23100 20085 23103
rect 19024 23072 20085 23100
rect 19024 23060 19030 23072
rect 20073 23069 20085 23072
rect 20119 23069 20131 23103
rect 20073 23063 20131 23069
rect 20714 23060 20720 23112
rect 20772 23100 20778 23112
rect 21453 23103 21511 23109
rect 21453 23100 21465 23103
rect 20772 23072 21465 23100
rect 20772 23060 20778 23072
rect 21453 23069 21465 23072
rect 21499 23069 21511 23103
rect 21453 23063 21511 23069
rect 12308 23004 13584 23032
rect 13633 23035 13691 23041
rect 12308 22992 12314 23004
rect 13633 23001 13645 23035
rect 13679 23032 13691 23035
rect 13814 23032 13820 23044
rect 13679 23004 13820 23032
rect 13679 23001 13691 23004
rect 13633 22995 13691 23001
rect 13814 22992 13820 23004
rect 13872 23032 13878 23044
rect 14550 23032 14556 23044
rect 13872 23004 14556 23032
rect 13872 22992 13878 23004
rect 14550 22992 14556 23004
rect 14608 22992 14614 23044
rect 14660 23004 15042 23032
rect 1854 22924 1860 22976
rect 1912 22964 1918 22976
rect 1949 22967 2007 22973
rect 1949 22964 1961 22967
rect 1912 22936 1961 22964
rect 1912 22924 1918 22936
rect 1949 22933 1961 22936
rect 1995 22933 2007 22967
rect 1949 22927 2007 22933
rect 5353 22967 5411 22973
rect 5353 22933 5365 22967
rect 5399 22964 5411 22967
rect 5534 22964 5540 22976
rect 5399 22936 5540 22964
rect 5399 22933 5411 22936
rect 5353 22927 5411 22933
rect 5534 22924 5540 22936
rect 5592 22924 5598 22976
rect 7006 22924 7012 22976
rect 7064 22964 7070 22976
rect 7377 22967 7435 22973
rect 7377 22964 7389 22967
rect 7064 22936 7389 22964
rect 7064 22924 7070 22936
rect 7377 22933 7389 22936
rect 7423 22933 7435 22967
rect 7377 22927 7435 22933
rect 7558 22924 7564 22976
rect 7616 22964 7622 22976
rect 12161 22967 12219 22973
rect 12161 22964 12173 22967
rect 7616 22936 12173 22964
rect 7616 22924 7622 22936
rect 12161 22933 12173 22936
rect 12207 22933 12219 22967
rect 12161 22927 12219 22933
rect 13722 22924 13728 22976
rect 13780 22964 13786 22976
rect 14660 22964 14688 23004
rect 20806 22992 20812 23044
rect 20864 23032 20870 23044
rect 20990 23032 20996 23044
rect 20864 23004 20996 23032
rect 20864 22992 20870 23004
rect 20990 22992 20996 23004
rect 21048 22992 21054 23044
rect 13780 22936 14688 22964
rect 13780 22924 13786 22936
rect 14734 22924 14740 22976
rect 14792 22964 14798 22976
rect 16025 22967 16083 22973
rect 16025 22964 16037 22967
rect 14792 22936 16037 22964
rect 14792 22924 14798 22936
rect 16025 22933 16037 22936
rect 16071 22933 16083 22967
rect 16025 22927 16083 22933
rect 16574 22924 16580 22976
rect 16632 22964 16638 22976
rect 17402 22964 17408 22976
rect 16632 22936 17408 22964
rect 16632 22924 16638 22936
rect 17402 22924 17408 22936
rect 17460 22964 17466 22976
rect 22066 22964 22094 23140
rect 24394 23060 24400 23112
rect 24452 23060 24458 23112
rect 25792 23109 25820 23140
rect 31110 23128 31116 23140
rect 31168 23128 31174 23180
rect 25777 23103 25835 23109
rect 25777 23069 25789 23103
rect 25823 23069 25835 23103
rect 25777 23063 25835 23069
rect 29733 23103 29791 23109
rect 29733 23069 29745 23103
rect 29779 23069 29791 23103
rect 29733 23063 29791 23069
rect 22646 23032 22652 23044
rect 22607 23004 22652 23032
rect 22646 22992 22652 23004
rect 22704 22992 22710 23044
rect 22738 22992 22744 23044
rect 22796 23032 22802 23044
rect 22796 23004 22841 23032
rect 22796 22992 22802 23004
rect 23014 22992 23020 23044
rect 23072 23032 23078 23044
rect 23661 23035 23719 23041
rect 23661 23032 23673 23035
rect 23072 23004 23673 23032
rect 23072 22992 23078 23004
rect 23661 23001 23673 23004
rect 23707 23032 23719 23035
rect 23934 23032 23940 23044
rect 23707 23004 23940 23032
rect 23707 23001 23719 23004
rect 23661 22995 23719 23001
rect 23934 22992 23940 23004
rect 23992 22992 23998 23044
rect 24412 23032 24440 23060
rect 24673 23035 24731 23041
rect 24673 23032 24685 23035
rect 24044 23004 24685 23032
rect 17460 22936 22094 22964
rect 17460 22924 17466 22936
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 24044 22964 24072 23004
rect 24673 23001 24685 23004
rect 24719 23001 24731 23035
rect 24673 22995 24731 23001
rect 24762 22992 24768 23044
rect 24820 23032 24826 23044
rect 24820 23004 24865 23032
rect 24820 22992 24826 23004
rect 23532 22936 24072 22964
rect 23532 22924 23538 22936
rect 24394 22924 24400 22976
rect 24452 22964 24458 22976
rect 25869 22967 25927 22973
rect 25869 22964 25881 22967
rect 24452 22936 25881 22964
rect 24452 22924 24458 22936
rect 25869 22933 25881 22936
rect 25915 22933 25927 22967
rect 26418 22964 26424 22976
rect 26379 22936 26424 22964
rect 25869 22927 25927 22933
rect 26418 22924 26424 22936
rect 26476 22924 26482 22976
rect 29748 22964 29776 23063
rect 36078 23060 36084 23112
rect 36136 23100 36142 23112
rect 38013 23103 38071 23109
rect 38013 23100 38025 23103
rect 36136 23072 38025 23100
rect 36136 23060 36142 23072
rect 38013 23069 38025 23072
rect 38059 23069 38071 23103
rect 38013 23063 38071 23069
rect 30282 22992 30288 23044
rect 30340 23032 30346 23044
rect 31205 23035 31263 23041
rect 31205 23032 31217 23035
rect 30340 23004 31217 23032
rect 30340 22992 30346 23004
rect 31205 23001 31217 23004
rect 31251 23001 31263 23035
rect 32122 23032 32128 23044
rect 32083 23004 32128 23032
rect 31205 22995 31263 23001
rect 32122 22992 32128 23004
rect 32180 22992 32186 23044
rect 37642 22964 37648 22976
rect 29748 22936 37648 22964
rect 37642 22924 37648 22936
rect 37700 22924 37706 22976
rect 37829 22967 37887 22973
rect 37829 22933 37841 22967
rect 37875 22964 37887 22967
rect 38010 22964 38016 22976
rect 37875 22936 38016 22964
rect 37875 22933 37887 22936
rect 37829 22927 37887 22933
rect 38010 22924 38016 22936
rect 38068 22924 38074 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 2406 22760 2412 22772
rect 1780 22732 2412 22760
rect 1780 22633 1808 22732
rect 2406 22720 2412 22732
rect 2464 22760 2470 22772
rect 3694 22760 3700 22772
rect 2464 22732 3700 22760
rect 2464 22720 2470 22732
rect 3694 22720 3700 22732
rect 3752 22720 3758 22772
rect 10686 22760 10692 22772
rect 8036 22732 10692 22760
rect 2038 22652 2044 22704
rect 2096 22692 2102 22704
rect 8036 22701 8064 22732
rect 10686 22720 10692 22732
rect 10744 22720 10750 22772
rect 10778 22720 10784 22772
rect 10836 22760 10842 22772
rect 17218 22760 17224 22772
rect 10836 22732 17224 22760
rect 10836 22720 10842 22732
rect 17218 22720 17224 22732
rect 17276 22720 17282 22772
rect 28442 22760 28448 22772
rect 25608 22732 28448 22760
rect 8021 22695 8079 22701
rect 2096 22664 2530 22692
rect 2096 22652 2102 22664
rect 8021 22661 8033 22695
rect 8067 22661 8079 22695
rect 8021 22655 8079 22661
rect 9582 22652 9588 22704
rect 9640 22692 9646 22704
rect 12434 22692 12440 22704
rect 9640 22664 12440 22692
rect 9640 22652 9646 22664
rect 12434 22652 12440 22664
rect 12492 22652 12498 22704
rect 12529 22695 12587 22701
rect 12529 22661 12541 22695
rect 12575 22692 12587 22695
rect 12802 22692 12808 22704
rect 12575 22664 12808 22692
rect 12575 22661 12587 22664
rect 12529 22655 12587 22661
rect 12802 22652 12808 22664
rect 12860 22652 12866 22704
rect 14182 22652 14188 22704
rect 14240 22692 14246 22704
rect 14277 22695 14335 22701
rect 14277 22692 14289 22695
rect 14240 22664 14289 22692
rect 14240 22652 14246 22664
rect 14277 22661 14289 22664
rect 14323 22661 14335 22695
rect 14277 22655 14335 22661
rect 14550 22652 14556 22704
rect 14608 22692 14614 22704
rect 18230 22692 18236 22704
rect 14608 22664 18236 22692
rect 14608 22652 14614 22664
rect 18230 22652 18236 22664
rect 18288 22652 18294 22704
rect 21358 22692 21364 22704
rect 18524 22664 21364 22692
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22593 1823 22627
rect 1765 22587 1823 22593
rect 6914 22584 6920 22636
rect 6972 22624 6978 22636
rect 7466 22624 7472 22636
rect 6972 22596 7472 22624
rect 6972 22584 6978 22596
rect 7466 22584 7472 22596
rect 7524 22624 7530 22636
rect 7745 22627 7803 22633
rect 7745 22624 7757 22627
rect 7524 22596 7757 22624
rect 7524 22584 7530 22596
rect 7745 22593 7757 22596
rect 7791 22593 7803 22627
rect 12250 22624 12256 22636
rect 7745 22587 7803 22593
rect 2041 22559 2099 22565
rect 2041 22525 2053 22559
rect 2087 22556 2099 22559
rect 7098 22556 7104 22568
rect 2087 22528 7104 22556
rect 2087 22525 2099 22528
rect 2041 22519 2099 22525
rect 7098 22516 7104 22528
rect 7156 22516 7162 22568
rect 9140 22488 9168 22610
rect 12211 22596 12256 22624
rect 12250 22584 12256 22596
rect 12308 22584 12314 22636
rect 18524 22624 18552 22664
rect 21358 22652 21364 22664
rect 21416 22652 21422 22704
rect 24394 22692 24400 22704
rect 24355 22664 24400 22692
rect 24394 22652 24400 22664
rect 24452 22652 24458 22704
rect 24946 22692 24952 22704
rect 24907 22664 24952 22692
rect 24946 22652 24952 22664
rect 25004 22652 25010 22704
rect 25608 22701 25636 22732
rect 28442 22720 28448 22732
rect 28500 22720 28506 22772
rect 36078 22760 36084 22772
rect 36039 22732 36084 22760
rect 36078 22720 36084 22732
rect 36136 22720 36142 22772
rect 25593 22695 25651 22701
rect 25593 22661 25605 22695
rect 25639 22661 25651 22695
rect 25593 22655 25651 22661
rect 25685 22695 25743 22701
rect 25685 22661 25697 22695
rect 25731 22692 25743 22695
rect 27249 22695 27307 22701
rect 27249 22692 27261 22695
rect 25731 22664 27261 22692
rect 25731 22661 25743 22664
rect 25685 22655 25743 22661
rect 27249 22661 27261 22664
rect 27295 22661 27307 22695
rect 27249 22655 27307 22661
rect 13662 22596 18552 22624
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22624 18659 22627
rect 18690 22624 18696 22636
rect 18647 22596 18696 22624
rect 18647 22593 18659 22596
rect 18601 22587 18659 22593
rect 9490 22556 9496 22568
rect 9451 22528 9496 22556
rect 9490 22516 9496 22528
rect 9548 22516 9554 22568
rect 12618 22516 12624 22568
rect 12676 22556 12682 22568
rect 18616 22556 18644 22587
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 27157 22627 27215 22633
rect 27157 22593 27169 22627
rect 27203 22624 27215 22627
rect 27338 22624 27344 22636
rect 27203 22596 27344 22624
rect 27203 22593 27215 22596
rect 27157 22587 27215 22593
rect 27338 22584 27344 22596
rect 27396 22584 27402 22636
rect 30834 22584 30840 22636
rect 30892 22624 30898 22636
rect 35989 22627 36047 22633
rect 35989 22624 36001 22627
rect 30892 22596 36001 22624
rect 30892 22584 30898 22596
rect 35989 22593 36001 22596
rect 36035 22593 36047 22627
rect 38010 22624 38016 22636
rect 37971 22596 38016 22624
rect 35989 22587 36047 22593
rect 38010 22584 38016 22596
rect 38068 22584 38074 22636
rect 24302 22556 24308 22568
rect 12676 22528 18644 22556
rect 24263 22528 24308 22556
rect 12676 22516 12682 22528
rect 24302 22516 24308 22528
rect 24360 22516 24366 22568
rect 26602 22556 26608 22568
rect 26563 22528 26608 22556
rect 26602 22516 26608 22528
rect 26660 22516 26666 22568
rect 18782 22488 18788 22500
rect 9140 22460 10824 22488
rect 3418 22380 3424 22432
rect 3476 22420 3482 22432
rect 3513 22423 3571 22429
rect 3513 22420 3525 22423
rect 3476 22392 3525 22420
rect 3476 22380 3482 22392
rect 3513 22389 3525 22392
rect 3559 22389 3571 22423
rect 10796 22420 10824 22460
rect 15580 22460 18788 22488
rect 15580 22420 15608 22460
rect 18782 22448 18788 22460
rect 18840 22448 18846 22500
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 10796 22392 15608 22420
rect 3513 22383 3571 22389
rect 17586 22380 17592 22432
rect 17644 22420 17650 22432
rect 18693 22423 18751 22429
rect 18693 22420 18705 22423
rect 17644 22392 18705 22420
rect 17644 22380 17650 22392
rect 18693 22389 18705 22392
rect 18739 22389 18751 22423
rect 18693 22383 18751 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 3602 22176 3608 22228
rect 3660 22216 3666 22228
rect 4230 22219 4288 22225
rect 4230 22216 4242 22219
rect 3660 22188 4242 22216
rect 3660 22176 3666 22188
rect 4230 22185 4242 22188
rect 4276 22185 4288 22219
rect 4230 22179 4288 22185
rect 7088 22219 7146 22225
rect 7088 22185 7100 22219
rect 7134 22216 7146 22219
rect 7466 22216 7472 22228
rect 7134 22188 7472 22216
rect 7134 22185 7146 22188
rect 7088 22179 7146 22185
rect 7466 22176 7472 22188
rect 7524 22216 7530 22228
rect 8202 22216 8208 22228
rect 7524 22188 8208 22216
rect 7524 22176 7530 22188
rect 8202 22176 8208 22188
rect 8260 22176 8266 22228
rect 12158 22176 12164 22228
rect 12216 22216 12222 22228
rect 14734 22216 14740 22228
rect 12216 22188 14740 22216
rect 12216 22176 12222 22188
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 8110 22108 8116 22160
rect 8168 22148 8174 22160
rect 13814 22148 13820 22160
rect 8168 22120 8248 22148
rect 8168 22108 8174 22120
rect 3694 22040 3700 22092
rect 3752 22080 3758 22092
rect 3973 22083 4031 22089
rect 3973 22080 3985 22083
rect 3752 22052 3985 22080
rect 3752 22040 3758 22052
rect 3973 22049 3985 22052
rect 4019 22049 4031 22083
rect 3973 22043 4031 22049
rect 5258 22040 5264 22092
rect 5316 22080 5322 22092
rect 5721 22083 5779 22089
rect 5721 22080 5733 22083
rect 5316 22052 5733 22080
rect 5316 22040 5322 22052
rect 5721 22049 5733 22052
rect 5767 22049 5779 22083
rect 6822 22080 6828 22092
rect 6783 22052 6828 22080
rect 5721 22043 5779 22049
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 8220 22080 8248 22120
rect 11624 22120 13820 22148
rect 11514 22080 11520 22092
rect 8220 22052 11520 22080
rect 11514 22040 11520 22052
rect 11572 22040 11578 22092
rect 1578 22012 1584 22024
rect 1539 21984 1584 22012
rect 1578 21972 1584 21984
rect 1636 21972 1642 22024
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 10229 22015 10287 22021
rect 10229 22012 10241 22015
rect 8444 21984 10241 22012
rect 8444 21972 8450 21984
rect 10229 21981 10241 21984
rect 10275 22012 10287 22015
rect 11624 22012 11652 22120
rect 13814 22108 13820 22120
rect 13872 22108 13878 22160
rect 26878 22148 26884 22160
rect 25792 22120 26884 22148
rect 23382 22080 23388 22092
rect 13832 22052 23388 22080
rect 10275 21984 11652 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 11790 21972 11796 22024
rect 11848 22012 11854 22024
rect 12342 22012 12348 22024
rect 11848 21984 12348 22012
rect 11848 21972 11854 21984
rect 12342 21972 12348 21984
rect 12400 22012 12406 22024
rect 13832 22012 13860 22052
rect 23382 22040 23388 22052
rect 23440 22040 23446 22092
rect 25792 22080 25820 22120
rect 26878 22108 26884 22120
rect 26936 22108 26942 22160
rect 23952 22052 25820 22080
rect 25869 22083 25927 22089
rect 15102 22012 15108 22024
rect 12400 21984 13860 22012
rect 15063 21984 15108 22012
rect 12400 21972 12406 21984
rect 15102 21972 15108 21984
rect 15160 21972 15166 22024
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 22012 19487 22015
rect 20070 22012 20076 22024
rect 19475 21984 20076 22012
rect 19475 21981 19487 21984
rect 19429 21975 19487 21981
rect 20070 21972 20076 21984
rect 20128 21972 20134 22024
rect 21821 22015 21879 22021
rect 21821 21981 21833 22015
rect 21867 22012 21879 22015
rect 22094 22012 22100 22024
rect 21867 21984 22100 22012
rect 21867 21981 21879 21984
rect 21821 21975 21879 21981
rect 22094 21972 22100 21984
rect 22152 21972 22158 22024
rect 4706 21904 4712 21956
rect 4764 21904 4770 21956
rect 5534 21904 5540 21956
rect 5592 21944 5598 21956
rect 5592 21916 7590 21944
rect 5592 21904 5598 21916
rect 11514 21904 11520 21956
rect 11572 21944 11578 21956
rect 12710 21944 12716 21956
rect 11572 21916 12716 21944
rect 11572 21904 11578 21916
rect 12710 21904 12716 21916
rect 12768 21904 12774 21956
rect 15378 21944 15384 21956
rect 15339 21916 15384 21944
rect 15378 21904 15384 21916
rect 15436 21904 15442 21956
rect 17586 21944 17592 21956
rect 16606 21916 17592 21944
rect 17586 21904 17592 21916
rect 17644 21904 17650 21956
rect 20162 21904 20168 21956
rect 20220 21944 20226 21956
rect 23952 21944 23980 22052
rect 25869 22049 25881 22083
rect 25915 22080 25927 22083
rect 26418 22080 26424 22092
rect 25915 22052 26424 22080
rect 25915 22049 25927 22052
rect 25869 22043 25927 22049
rect 26418 22040 26424 22052
rect 26476 22040 26482 22092
rect 28166 22080 28172 22092
rect 26896 22052 28172 22080
rect 26896 21956 26924 22052
rect 28166 22040 28172 22052
rect 28224 22040 28230 22092
rect 27341 22015 27399 22021
rect 27341 21981 27353 22015
rect 27387 22012 27399 22015
rect 27430 22012 27436 22024
rect 27387 21984 27436 22012
rect 27387 21981 27399 21984
rect 27341 21975 27399 21981
rect 27430 21972 27436 21984
rect 27488 21972 27494 22024
rect 27985 22015 28043 22021
rect 27985 21981 27997 22015
rect 28031 22012 28043 22015
rect 28442 22012 28448 22024
rect 28031 21984 28448 22012
rect 28031 21981 28043 21984
rect 27985 21975 28043 21981
rect 20220 21916 23980 21944
rect 20220 21904 20226 21916
rect 25958 21904 25964 21956
rect 26016 21944 26022 21956
rect 26878 21944 26884 21956
rect 26016 21916 26061 21944
rect 26839 21916 26884 21944
rect 26016 21904 26022 21916
rect 26878 21904 26884 21916
rect 26936 21904 26942 21956
rect 26970 21904 26976 21956
rect 27028 21944 27034 21956
rect 28000 21944 28028 21975
rect 28442 21972 28448 21984
rect 28500 21972 28506 22024
rect 29733 22015 29791 22021
rect 29733 21981 29745 22015
rect 29779 22012 29791 22015
rect 36630 22012 36636 22024
rect 29779 21984 36636 22012
rect 29779 21981 29791 21984
rect 29733 21975 29791 21981
rect 36630 21972 36636 21984
rect 36688 21972 36694 22024
rect 27028 21916 28028 21944
rect 27028 21904 27034 21916
rect 1762 21876 1768 21888
rect 1723 21848 1768 21876
rect 1762 21836 1768 21848
rect 1820 21836 1826 21888
rect 8110 21836 8116 21888
rect 8168 21876 8174 21888
rect 8573 21879 8631 21885
rect 8573 21876 8585 21879
rect 8168 21848 8585 21876
rect 8168 21836 8174 21848
rect 8573 21845 8585 21848
rect 8619 21876 8631 21879
rect 8754 21876 8760 21888
rect 8619 21848 8760 21876
rect 8619 21845 8631 21848
rect 8573 21839 8631 21845
rect 8754 21836 8760 21848
rect 8812 21836 8818 21888
rect 8938 21836 8944 21888
rect 8996 21876 9002 21888
rect 10321 21879 10379 21885
rect 10321 21876 10333 21879
rect 8996 21848 10333 21876
rect 8996 21836 9002 21848
rect 10321 21845 10333 21848
rect 10367 21845 10379 21879
rect 10321 21839 10379 21845
rect 10410 21836 10416 21888
rect 10468 21876 10474 21888
rect 16853 21879 16911 21885
rect 16853 21876 16865 21879
rect 10468 21848 16865 21876
rect 10468 21836 10474 21848
rect 16853 21845 16865 21848
rect 16899 21876 16911 21879
rect 17310 21876 17316 21888
rect 16899 21848 17316 21876
rect 16899 21845 16911 21848
rect 16853 21839 16911 21845
rect 17310 21836 17316 21848
rect 17368 21836 17374 21888
rect 17862 21836 17868 21888
rect 17920 21876 17926 21888
rect 19521 21879 19579 21885
rect 19521 21876 19533 21879
rect 17920 21848 19533 21876
rect 17920 21836 17926 21848
rect 19521 21845 19533 21848
rect 19567 21845 19579 21879
rect 19521 21839 19579 21845
rect 20622 21836 20628 21888
rect 20680 21876 20686 21888
rect 21913 21879 21971 21885
rect 21913 21876 21925 21879
rect 20680 21848 21925 21876
rect 20680 21836 20686 21848
rect 21913 21845 21925 21848
rect 21959 21845 21971 21879
rect 21913 21839 21971 21845
rect 26234 21836 26240 21888
rect 26292 21876 26298 21888
rect 27433 21879 27491 21885
rect 27433 21876 27445 21879
rect 26292 21848 27445 21876
rect 26292 21836 26298 21848
rect 27433 21845 27445 21848
rect 27479 21845 27491 21879
rect 27433 21839 27491 21845
rect 27982 21836 27988 21888
rect 28040 21876 28046 21888
rect 28077 21879 28135 21885
rect 28077 21876 28089 21879
rect 28040 21848 28089 21876
rect 28040 21836 28046 21848
rect 28077 21845 28089 21848
rect 28123 21845 28135 21879
rect 29822 21876 29828 21888
rect 29783 21848 29828 21876
rect 28077 21839 28135 21845
rect 29822 21836 29828 21848
rect 29880 21836 29886 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 4982 21632 4988 21684
rect 5040 21672 5046 21684
rect 5166 21672 5172 21684
rect 5040 21644 5172 21672
rect 5040 21632 5046 21644
rect 5166 21632 5172 21644
rect 5224 21632 5230 21684
rect 5258 21632 5264 21684
rect 5316 21672 5322 21684
rect 7374 21672 7380 21684
rect 5316 21644 7380 21672
rect 5316 21632 5322 21644
rect 7374 21632 7380 21644
rect 7432 21632 7438 21684
rect 7558 21632 7564 21684
rect 7616 21672 7622 21684
rect 8018 21672 8024 21684
rect 7616 21644 8024 21672
rect 7616 21632 7622 21644
rect 8018 21632 8024 21644
rect 8076 21632 8082 21684
rect 8202 21632 8208 21684
rect 8260 21672 8266 21684
rect 17770 21672 17776 21684
rect 8260 21644 11284 21672
rect 8260 21632 8266 21644
rect 7190 21564 7196 21616
rect 7248 21604 7254 21616
rect 7248 21576 7682 21604
rect 7248 21564 7254 21576
rect 9858 21564 9864 21616
rect 9916 21564 9922 21616
rect 1762 21536 1768 21548
rect 1723 21508 1768 21536
rect 1762 21496 1768 21508
rect 1820 21496 1826 21548
rect 3970 21536 3976 21548
rect 3931 21508 3976 21536
rect 3970 21496 3976 21508
rect 4028 21496 4034 21548
rect 5350 21496 5356 21548
rect 5408 21496 5414 21548
rect 4246 21468 4252 21480
rect 4207 21440 4252 21468
rect 4246 21428 4252 21440
rect 4304 21428 4310 21480
rect 4706 21428 4712 21480
rect 4764 21468 4770 21480
rect 4982 21468 4988 21480
rect 4764 21440 4988 21468
rect 4764 21428 4770 21440
rect 4982 21428 4988 21440
rect 5040 21428 5046 21480
rect 5994 21468 6000 21480
rect 5955 21440 6000 21468
rect 5994 21428 6000 21440
rect 6052 21428 6058 21480
rect 6822 21428 6828 21480
rect 6880 21468 6886 21480
rect 6917 21471 6975 21477
rect 6917 21468 6929 21471
rect 6880 21440 6929 21468
rect 6880 21428 6886 21440
rect 6917 21437 6929 21440
rect 6963 21437 6975 21471
rect 6917 21431 6975 21437
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 7558 21468 7564 21480
rect 7239 21440 7564 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 7558 21428 7564 21440
rect 7616 21428 7622 21480
rect 8478 21428 8484 21480
rect 8536 21468 8542 21480
rect 9125 21471 9183 21477
rect 9125 21468 9137 21471
rect 8536 21440 9137 21468
rect 8536 21428 8542 21440
rect 9125 21437 9137 21440
rect 9171 21437 9183 21471
rect 9401 21471 9459 21477
rect 9401 21468 9413 21471
rect 9125 21431 9183 21437
rect 9232 21440 9413 21468
rect 9232 21400 9260 21440
rect 9401 21437 9413 21440
rect 9447 21437 9459 21471
rect 9401 21431 9459 21437
rect 10686 21428 10692 21480
rect 10744 21468 10750 21480
rect 11149 21471 11207 21477
rect 11149 21468 11161 21471
rect 10744 21440 11161 21468
rect 10744 21428 10750 21440
rect 11149 21437 11161 21440
rect 11195 21437 11207 21471
rect 11256 21468 11284 21644
rect 11992 21644 14136 21672
rect 11992 21545 12020 21644
rect 12710 21564 12716 21616
rect 12768 21564 12774 21616
rect 14108 21548 14136 21644
rect 17144 21644 17776 21672
rect 14185 21607 14243 21613
rect 14185 21573 14197 21607
rect 14231 21604 14243 21607
rect 15194 21604 15200 21616
rect 14231 21576 15200 21604
rect 14231 21573 14243 21576
rect 14185 21567 14243 21573
rect 15194 21564 15200 21576
rect 15252 21564 15258 21616
rect 17144 21613 17172 21644
rect 17770 21632 17776 21644
rect 17828 21672 17834 21684
rect 17828 21644 22094 21672
rect 17828 21632 17834 21644
rect 17129 21607 17187 21613
rect 17129 21573 17141 21607
rect 17175 21573 17187 21607
rect 20073 21607 20131 21613
rect 20073 21604 20085 21607
rect 18354 21576 20085 21604
rect 17129 21567 17187 21573
rect 20073 21573 20085 21576
rect 20119 21573 20131 21607
rect 22066 21604 22094 21644
rect 25406 21632 25412 21684
rect 25464 21672 25470 21684
rect 29822 21672 29828 21684
rect 25464 21644 29828 21672
rect 25464 21632 25470 21644
rect 29822 21632 29828 21644
rect 29880 21632 29886 21684
rect 25130 21604 25136 21616
rect 22066 21576 25136 21604
rect 20073 21567 20131 21573
rect 25130 21564 25136 21576
rect 25188 21604 25194 21616
rect 25590 21604 25596 21616
rect 25188 21576 25596 21604
rect 25188 21564 25194 21576
rect 25590 21564 25596 21576
rect 25648 21564 25654 21616
rect 27982 21604 27988 21616
rect 27943 21576 27988 21604
rect 27982 21564 27988 21576
rect 28040 21564 28046 21616
rect 11977 21539 12035 21545
rect 11977 21505 11989 21539
rect 12023 21505 12035 21539
rect 14090 21536 14096 21548
rect 14003 21508 14096 21536
rect 11977 21499 12035 21505
rect 14090 21496 14096 21508
rect 14148 21536 14154 21548
rect 14921 21539 14979 21545
rect 14921 21536 14933 21539
rect 14148 21508 14933 21536
rect 14148 21496 14154 21508
rect 14921 21505 14933 21508
rect 14967 21536 14979 21539
rect 15102 21536 15108 21548
rect 14967 21508 15108 21536
rect 14967 21505 14979 21508
rect 14921 21499 14979 21505
rect 15102 21496 15108 21508
rect 15160 21536 15166 21548
rect 16574 21536 16580 21548
rect 15160 21508 16580 21536
rect 15160 21496 15166 21508
rect 16574 21496 16580 21508
rect 16632 21536 16638 21548
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16632 21508 16865 21536
rect 16632 21496 16638 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 19153 21539 19211 21545
rect 19153 21505 19165 21539
rect 19199 21505 19211 21539
rect 19153 21499 19211 21505
rect 19981 21539 20039 21545
rect 19981 21505 19993 21539
rect 20027 21536 20039 21539
rect 20717 21539 20775 21545
rect 20717 21536 20729 21539
rect 20027 21508 20729 21536
rect 20027 21505 20039 21508
rect 19981 21499 20039 21505
rect 20717 21505 20729 21508
rect 20763 21536 20775 21539
rect 20898 21536 20904 21548
rect 20763 21508 20904 21536
rect 20763 21505 20775 21508
rect 20717 21499 20775 21505
rect 19168 21468 19196 21499
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 23382 21536 23388 21548
rect 23343 21508 23388 21536
rect 23382 21496 23388 21508
rect 23440 21496 23446 21548
rect 26513 21539 26571 21545
rect 26513 21505 26525 21539
rect 26559 21536 26571 21539
rect 26694 21536 26700 21548
rect 26559 21508 26700 21536
rect 26559 21505 26571 21508
rect 26513 21499 26571 21505
rect 26694 21496 26700 21508
rect 26752 21496 26758 21548
rect 38286 21536 38292 21548
rect 38247 21508 38292 21536
rect 38286 21496 38292 21508
rect 38344 21496 38350 21548
rect 11256 21440 15792 21468
rect 11149 21431 11207 21437
rect 8496 21372 9260 21400
rect 11164 21400 11192 21431
rect 11790 21400 11796 21412
rect 11164 21372 11796 21400
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 2222 21332 2228 21344
rect 1627 21304 2228 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 2222 21292 2228 21304
rect 2280 21292 2286 21344
rect 2498 21292 2504 21344
rect 2556 21332 2562 21344
rect 4890 21332 4896 21344
rect 2556 21304 4896 21332
rect 2556 21292 2562 21304
rect 4890 21292 4896 21304
rect 4948 21292 4954 21344
rect 5718 21292 5724 21344
rect 5776 21332 5782 21344
rect 8496 21332 8524 21372
rect 11790 21360 11796 21372
rect 11848 21360 11854 21412
rect 8662 21332 8668 21344
rect 5776 21304 8524 21332
rect 8623 21304 8668 21332
rect 5776 21292 5782 21304
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 8754 21292 8760 21344
rect 8812 21332 8818 21344
rect 12234 21335 12292 21341
rect 12234 21332 12246 21335
rect 8812 21304 12246 21332
rect 8812 21292 8818 21304
rect 12234 21301 12246 21304
rect 12280 21301 12292 21335
rect 12234 21295 12292 21301
rect 12342 21292 12348 21344
rect 12400 21332 12406 21344
rect 13725 21335 13783 21341
rect 13725 21332 13737 21335
rect 12400 21304 13737 21332
rect 12400 21292 12406 21304
rect 13725 21301 13737 21304
rect 13771 21301 13783 21335
rect 15764 21332 15792 21440
rect 18156 21440 19196 21468
rect 18156 21332 18184 21440
rect 19242 21428 19248 21480
rect 19300 21468 19306 21480
rect 20809 21471 20867 21477
rect 20809 21468 20821 21471
rect 19300 21440 20821 21468
rect 19300 21428 19306 21440
rect 20809 21437 20821 21440
rect 20855 21437 20867 21471
rect 20809 21431 20867 21437
rect 27893 21471 27951 21477
rect 27893 21437 27905 21471
rect 27939 21468 27951 21471
rect 28074 21468 28080 21480
rect 27939 21440 28080 21468
rect 27939 21437 27951 21440
rect 27893 21431 27951 21437
rect 28074 21428 28080 21440
rect 28132 21428 28138 21480
rect 28169 21471 28227 21477
rect 28169 21437 28181 21471
rect 28215 21437 28227 21471
rect 28169 21431 28227 21437
rect 22002 21400 22008 21412
rect 18616 21372 22008 21400
rect 15764 21304 18184 21332
rect 13725 21295 13783 21301
rect 18506 21292 18512 21344
rect 18564 21332 18570 21344
rect 18616 21341 18644 21372
rect 22002 21360 22008 21372
rect 22060 21360 22066 21412
rect 23477 21403 23535 21409
rect 23477 21369 23489 21403
rect 23523 21400 23535 21403
rect 26418 21400 26424 21412
rect 23523 21372 26424 21400
rect 23523 21369 23535 21372
rect 23477 21363 23535 21369
rect 26418 21360 26424 21372
rect 26476 21360 26482 21412
rect 27798 21360 27804 21412
rect 27856 21400 27862 21412
rect 28184 21400 28212 21431
rect 27856 21372 28212 21400
rect 27856 21360 27862 21372
rect 18601 21335 18659 21341
rect 18601 21332 18613 21335
rect 18564 21304 18613 21332
rect 18564 21292 18570 21304
rect 18601 21301 18613 21304
rect 18647 21301 18659 21335
rect 18601 21295 18659 21301
rect 19245 21335 19303 21341
rect 19245 21301 19257 21335
rect 19291 21332 19303 21335
rect 19886 21332 19892 21344
rect 19291 21304 19892 21332
rect 19291 21301 19303 21304
rect 19245 21295 19303 21301
rect 19886 21292 19892 21304
rect 19944 21292 19950 21344
rect 26326 21332 26332 21344
rect 26287 21304 26332 21332
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 29730 21292 29736 21344
rect 29788 21332 29794 21344
rect 38105 21335 38163 21341
rect 38105 21332 38117 21335
rect 29788 21304 38117 21332
rect 29788 21292 29794 21304
rect 38105 21301 38117 21304
rect 38151 21301 38163 21335
rect 38105 21295 38163 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1844 21131 1902 21137
rect 1844 21097 1856 21131
rect 1890 21128 1902 21131
rect 6914 21128 6920 21140
rect 1890 21100 4568 21128
rect 1890 21097 1902 21100
rect 1844 21091 1902 21097
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20992 1639 20995
rect 3142 20992 3148 21004
rect 1627 20964 3148 20992
rect 1627 20961 1639 20964
rect 1581 20955 1639 20961
rect 3142 20952 3148 20964
rect 3200 20952 3206 21004
rect 4062 20856 4068 20868
rect 3082 20828 4068 20856
rect 4062 20816 4068 20828
rect 4120 20816 4126 20868
rect 3326 20788 3332 20800
rect 3287 20760 3332 20788
rect 3326 20748 3332 20760
rect 3384 20748 3390 20800
rect 4540 20788 4568 21100
rect 4632 21100 6920 21128
rect 4632 21001 4660 21100
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 9769 21131 9827 21137
rect 9769 21097 9781 21131
rect 9815 21128 9827 21131
rect 9858 21128 9864 21140
rect 9815 21100 9864 21128
rect 9815 21097 9827 21100
rect 9769 21091 9827 21097
rect 9858 21088 9864 21100
rect 9916 21088 9922 21140
rect 14918 21128 14924 21140
rect 10520 21100 14924 21128
rect 8573 21063 8631 21069
rect 8573 21029 8585 21063
rect 8619 21060 8631 21063
rect 10520 21060 10548 21100
rect 14918 21088 14924 21100
rect 14976 21088 14982 21140
rect 16390 21128 16396 21140
rect 16040 21100 16396 21128
rect 16040 21060 16068 21100
rect 16390 21088 16396 21100
rect 16448 21088 16454 21140
rect 17681 21131 17739 21137
rect 17681 21097 17693 21131
rect 17727 21128 17739 21131
rect 17770 21128 17776 21140
rect 17727 21100 17776 21128
rect 17727 21097 17739 21100
rect 17681 21091 17739 21097
rect 17770 21088 17776 21100
rect 17828 21088 17834 21140
rect 8619 21032 10548 21060
rect 12406 21032 16068 21060
rect 8619 21029 8631 21032
rect 8573 21023 8631 21029
rect 4617 20995 4675 21001
rect 4617 20961 4629 20995
rect 4663 20961 4675 20995
rect 4617 20955 4675 20961
rect 4893 20995 4951 21001
rect 4893 20961 4905 20995
rect 4939 20992 4951 20995
rect 10410 20992 10416 21004
rect 4939 20964 10416 20992
rect 4939 20961 4951 20964
rect 4893 20955 4951 20961
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20992 11299 20995
rect 12406 20992 12434 21032
rect 17218 21020 17224 21072
rect 17276 21060 17282 21072
rect 18506 21060 18512 21072
rect 17276 21032 18512 21060
rect 17276 21020 17282 21032
rect 18506 21020 18512 21032
rect 18564 21020 18570 21072
rect 22002 21020 22008 21072
rect 22060 21060 22066 21072
rect 27062 21060 27068 21072
rect 22060 21032 27068 21060
rect 22060 21020 22066 21032
rect 27062 21020 27068 21032
rect 27120 21020 27126 21072
rect 11287 20964 12434 20992
rect 11287 20961 11299 20964
rect 11241 20955 11299 20961
rect 15102 20952 15108 21004
rect 15160 20992 15166 21004
rect 15856 21001 15976 21004
rect 15856 20995 15991 21001
rect 15856 20992 15945 20995
rect 15160 20976 15945 20992
rect 15160 20964 15884 20976
rect 15160 20952 15166 20964
rect 15933 20961 15945 20976
rect 15979 20961 15991 20995
rect 16206 20992 16212 21004
rect 16167 20964 16212 20992
rect 15933 20955 15991 20961
rect 16206 20952 16212 20964
rect 16264 20952 16270 21004
rect 19794 20952 19800 21004
rect 19852 20992 19932 21004
rect 20714 20992 20720 21004
rect 19852 20976 20720 20992
rect 19852 20952 19858 20976
rect 19904 20964 20720 20976
rect 20714 20952 20720 20964
rect 20772 20992 20778 21004
rect 21082 20992 21088 21004
rect 20772 20964 21088 20992
rect 20772 20952 20778 20964
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 26970 20992 26976 21004
rect 22066 20964 26976 20992
rect 6822 20924 6828 20936
rect 6783 20896 6828 20924
rect 6822 20884 6828 20896
rect 6880 20884 6886 20936
rect 8938 20924 8944 20936
rect 8234 20896 8944 20924
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 9582 20884 9588 20936
rect 9640 20924 9646 20936
rect 9677 20927 9735 20933
rect 9677 20924 9689 20927
rect 9640 20896 9689 20924
rect 9640 20884 9646 20896
rect 9677 20893 9689 20896
rect 9723 20893 9735 20927
rect 9677 20887 9735 20893
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20924 10379 20927
rect 10502 20924 10508 20936
rect 10367 20896 10508 20924
rect 10367 20893 10379 20896
rect 10321 20887 10379 20893
rect 10502 20884 10508 20896
rect 10560 20884 10566 20936
rect 10962 20924 10968 20936
rect 10923 20896 10968 20924
rect 10962 20884 10968 20896
rect 11020 20884 11026 20936
rect 19242 20924 19248 20936
rect 17342 20896 19248 20924
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 7006 20856 7012 20868
rect 6118 20828 7012 20856
rect 7006 20816 7012 20828
rect 7064 20816 7070 20868
rect 7101 20859 7159 20865
rect 7101 20825 7113 20859
rect 7147 20856 7159 20859
rect 7374 20856 7380 20868
rect 7147 20828 7380 20856
rect 7147 20825 7159 20828
rect 7101 20819 7159 20825
rect 7374 20816 7380 20828
rect 7432 20816 7438 20868
rect 8570 20816 8576 20868
rect 8628 20856 8634 20868
rect 8628 20828 11468 20856
rect 8628 20816 8634 20828
rect 6270 20788 6276 20800
rect 4540 20760 6276 20788
rect 6270 20748 6276 20760
rect 6328 20788 6334 20800
rect 6365 20791 6423 20797
rect 6365 20788 6377 20791
rect 6328 20760 6377 20788
rect 6328 20748 6334 20760
rect 6365 20757 6377 20760
rect 6411 20757 6423 20791
rect 6365 20751 6423 20757
rect 6822 20748 6828 20800
rect 6880 20788 6886 20800
rect 8478 20788 8484 20800
rect 6880 20760 8484 20788
rect 6880 20748 6886 20760
rect 8478 20748 8484 20760
rect 8536 20748 8542 20800
rect 10413 20791 10471 20797
rect 10413 20757 10425 20791
rect 10459 20788 10471 20791
rect 11330 20788 11336 20800
rect 10459 20760 11336 20788
rect 10459 20757 10471 20760
rect 10413 20751 10471 20757
rect 11330 20748 11336 20760
rect 11388 20748 11394 20800
rect 11440 20788 11468 20828
rect 11698 20816 11704 20868
rect 11756 20816 11762 20868
rect 19794 20856 19800 20868
rect 12636 20828 16620 20856
rect 19755 20828 19800 20856
rect 12636 20788 12664 20828
rect 11440 20760 12664 20788
rect 12713 20791 12771 20797
rect 12713 20757 12725 20791
rect 12759 20788 12771 20791
rect 13814 20788 13820 20800
rect 12759 20760 13820 20788
rect 12759 20757 12771 20760
rect 12713 20751 12771 20757
rect 13814 20748 13820 20760
rect 13872 20748 13878 20800
rect 14918 20748 14924 20800
rect 14976 20788 14982 20800
rect 16206 20788 16212 20800
rect 14976 20760 16212 20788
rect 14976 20748 14982 20760
rect 16206 20748 16212 20760
rect 16264 20748 16270 20800
rect 16592 20788 16620 20828
rect 19794 20816 19800 20828
rect 19852 20816 19858 20868
rect 19886 20816 19892 20868
rect 19944 20856 19950 20868
rect 20809 20859 20867 20865
rect 19944 20828 19989 20856
rect 19944 20816 19950 20828
rect 20809 20825 20821 20859
rect 20855 20856 20867 20859
rect 22066 20856 22094 20964
rect 26970 20952 26976 20964
rect 27028 20952 27034 21004
rect 28261 20995 28319 21001
rect 28261 20961 28273 20995
rect 28307 20992 28319 20995
rect 29546 20992 29552 21004
rect 28307 20964 29552 20992
rect 28307 20961 28319 20964
rect 28261 20955 28319 20961
rect 29546 20952 29552 20964
rect 29604 20992 29610 21004
rect 29825 20995 29883 21001
rect 29825 20992 29837 20995
rect 29604 20964 29837 20992
rect 29604 20952 29610 20964
rect 29825 20961 29837 20964
rect 29871 20961 29883 20995
rect 29825 20955 29883 20961
rect 23658 20924 23664 20936
rect 23619 20896 23664 20924
rect 23658 20884 23664 20896
rect 23716 20884 23722 20936
rect 29730 20924 29736 20936
rect 29691 20896 29736 20924
rect 29730 20884 29736 20896
rect 29788 20884 29794 20936
rect 30377 20927 30435 20933
rect 30377 20893 30389 20927
rect 30423 20924 30435 20927
rect 37550 20924 37556 20936
rect 30423 20896 37556 20924
rect 30423 20893 30435 20896
rect 30377 20887 30435 20893
rect 37550 20884 37556 20896
rect 37608 20884 37614 20936
rect 38286 20924 38292 20936
rect 38247 20896 38292 20924
rect 38286 20884 38292 20896
rect 38344 20884 38350 20936
rect 20855 20828 22094 20856
rect 20855 20825 20867 20828
rect 20809 20819 20867 20825
rect 20824 20788 20852 20819
rect 25222 20816 25228 20868
rect 25280 20856 25286 20868
rect 26329 20859 26387 20865
rect 26329 20856 26341 20859
rect 25280 20828 26341 20856
rect 25280 20816 25286 20828
rect 26329 20825 26341 20828
rect 26375 20825 26387 20859
rect 26329 20819 26387 20825
rect 26418 20816 26424 20868
rect 26476 20856 26482 20868
rect 26476 20828 26521 20856
rect 26476 20816 26482 20828
rect 28350 20816 28356 20868
rect 28408 20856 28414 20868
rect 28902 20856 28908 20868
rect 28408 20828 28453 20856
rect 28863 20828 28908 20856
rect 28408 20816 28414 20828
rect 28902 20816 28908 20828
rect 28960 20816 28966 20868
rect 16592 20760 20852 20788
rect 23477 20791 23535 20797
rect 23477 20757 23489 20791
rect 23523 20788 23535 20791
rect 25774 20788 25780 20800
rect 23523 20760 25780 20788
rect 23523 20757 23535 20760
rect 23477 20751 23535 20757
rect 25774 20748 25780 20760
rect 25832 20748 25838 20800
rect 30466 20788 30472 20800
rect 30427 20760 30472 20788
rect 30466 20748 30472 20760
rect 30524 20748 30530 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1765 20587 1823 20593
rect 1765 20553 1777 20587
rect 1811 20584 1823 20587
rect 1811 20556 10732 20584
rect 1811 20553 1823 20556
rect 1765 20547 1823 20553
rect 1946 20476 1952 20528
rect 2004 20516 2010 20528
rect 2004 20488 3174 20516
rect 2004 20476 2010 20488
rect 6730 20476 6736 20528
rect 6788 20516 6794 20528
rect 7745 20519 7803 20525
rect 7745 20516 7757 20519
rect 6788 20488 7757 20516
rect 6788 20476 6794 20488
rect 7745 20485 7757 20488
rect 7791 20485 7803 20519
rect 8478 20516 8484 20528
rect 8439 20488 8484 20516
rect 7745 20479 7803 20485
rect 8478 20476 8484 20488
rect 8536 20476 8542 20528
rect 9674 20516 9680 20528
rect 9048 20488 9680 20516
rect 1394 20408 1400 20460
rect 1452 20448 1458 20460
rect 1673 20451 1731 20457
rect 1673 20448 1685 20451
rect 1452 20420 1685 20448
rect 1452 20408 1458 20420
rect 1673 20417 1685 20420
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 2409 20383 2467 20389
rect 2409 20349 2421 20383
rect 2455 20380 2467 20383
rect 2685 20383 2743 20389
rect 2455 20352 2544 20380
rect 2455 20349 2467 20352
rect 2409 20343 2467 20349
rect 2516 20244 2544 20352
rect 2685 20349 2697 20383
rect 2731 20380 2743 20383
rect 4614 20380 4620 20392
rect 2731 20352 4620 20380
rect 2731 20349 2743 20352
rect 2685 20343 2743 20349
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 3694 20272 3700 20324
rect 3752 20312 3758 20324
rect 9048 20312 9076 20488
rect 9674 20476 9680 20488
rect 9732 20476 9738 20528
rect 10410 20476 10416 20528
rect 10468 20476 10474 20528
rect 9125 20383 9183 20389
rect 9125 20349 9137 20383
rect 9171 20349 9183 20383
rect 9125 20343 9183 20349
rect 9401 20383 9459 20389
rect 9401 20349 9413 20383
rect 9447 20380 9459 20383
rect 10134 20380 10140 20392
rect 9447 20352 10140 20380
rect 9447 20349 9459 20352
rect 9401 20343 9459 20349
rect 3752 20284 9076 20312
rect 3752 20272 3758 20284
rect 3142 20244 3148 20256
rect 2516 20216 3148 20244
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 4157 20247 4215 20253
rect 4157 20213 4169 20247
rect 4203 20244 4215 20247
rect 4614 20244 4620 20256
rect 4203 20216 4620 20244
rect 4203 20213 4215 20216
rect 4157 20207 4215 20213
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 6638 20204 6644 20256
rect 6696 20244 6702 20256
rect 7742 20244 7748 20256
rect 6696 20216 7748 20244
rect 6696 20204 6702 20216
rect 7742 20204 7748 20216
rect 7800 20204 7806 20256
rect 9140 20244 9168 20343
rect 10134 20340 10140 20352
rect 10192 20340 10198 20392
rect 10704 20312 10732 20556
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 10836 20556 19104 20584
rect 10836 20544 10842 20556
rect 11882 20516 11888 20528
rect 11843 20488 11888 20516
rect 11882 20476 11888 20488
rect 11940 20476 11946 20528
rect 12526 20476 12532 20528
rect 12584 20516 12590 20528
rect 13722 20516 13728 20528
rect 12584 20488 13728 20516
rect 12584 20476 12590 20488
rect 13722 20476 13728 20488
rect 13780 20476 13786 20528
rect 14182 20476 14188 20528
rect 14240 20476 14246 20528
rect 15102 20476 15108 20528
rect 15160 20516 15166 20528
rect 18966 20516 18972 20528
rect 15160 20488 18972 20516
rect 15160 20476 15166 20488
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 12066 20408 12072 20460
rect 12124 20448 12130 20460
rect 12342 20448 12348 20460
rect 12124 20420 12348 20448
rect 12124 20408 12130 20420
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 13262 20408 13268 20460
rect 13320 20448 13326 20460
rect 13357 20451 13415 20457
rect 13357 20448 13369 20451
rect 13320 20420 13369 20448
rect 13320 20408 13326 20420
rect 13357 20417 13369 20420
rect 13403 20417 13415 20451
rect 13357 20411 13415 20417
rect 16482 20408 16488 20460
rect 16540 20448 16546 20460
rect 19076 20457 19104 20556
rect 23658 20544 23664 20596
rect 23716 20584 23722 20596
rect 24765 20587 24823 20593
rect 24765 20584 24777 20587
rect 23716 20556 24777 20584
rect 23716 20544 23722 20556
rect 24765 20553 24777 20556
rect 24811 20553 24823 20587
rect 30466 20584 30472 20596
rect 24765 20547 24823 20553
rect 27448 20556 30472 20584
rect 22554 20476 22560 20528
rect 22612 20516 22618 20528
rect 22925 20519 22983 20525
rect 22925 20516 22937 20519
rect 22612 20488 22937 20516
rect 22612 20476 22618 20488
rect 22925 20485 22937 20488
rect 22971 20485 22983 20519
rect 23750 20516 23756 20528
rect 23711 20488 23756 20516
rect 22925 20479 22983 20485
rect 23750 20476 23756 20488
rect 23808 20476 23814 20528
rect 25774 20516 25780 20528
rect 25735 20488 25780 20516
rect 25774 20476 25780 20488
rect 25832 20476 25838 20528
rect 27448 20516 27476 20556
rect 30466 20544 30472 20556
rect 30524 20544 30530 20596
rect 27264 20488 27476 20516
rect 28261 20519 28319 20525
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 16540 20420 16865 20448
rect 16540 20408 16546 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 19061 20451 19119 20457
rect 19061 20417 19073 20451
rect 19107 20417 19119 20451
rect 21818 20448 21824 20460
rect 19061 20411 19119 20417
rect 19306 20420 21824 20448
rect 10962 20340 10968 20392
rect 11020 20380 11026 20392
rect 12621 20383 12679 20389
rect 12621 20380 12633 20383
rect 11020 20352 12633 20380
rect 11020 20340 11026 20352
rect 12621 20349 12633 20352
rect 12667 20349 12679 20383
rect 13633 20383 13691 20389
rect 13633 20380 13645 20383
rect 12621 20343 12679 20349
rect 13280 20352 13645 20380
rect 13280 20324 13308 20352
rect 13633 20349 13645 20352
rect 13679 20349 13691 20383
rect 13633 20343 13691 20349
rect 13722 20340 13728 20392
rect 13780 20380 13786 20392
rect 19306 20380 19334 20420
rect 21818 20408 21824 20420
rect 21876 20408 21882 20460
rect 22002 20448 22008 20460
rect 21963 20420 22008 20448
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 24854 20408 24860 20460
rect 24912 20448 24918 20460
rect 24949 20451 25007 20457
rect 24949 20448 24961 20451
rect 24912 20420 24961 20448
rect 24912 20408 24918 20420
rect 24949 20417 24961 20420
rect 24995 20417 25007 20451
rect 24949 20411 25007 20417
rect 13780 20352 19334 20380
rect 22112 20352 23244 20380
rect 13780 20340 13786 20352
rect 10704 20284 12434 20312
rect 9766 20244 9772 20256
rect 9140 20216 9772 20244
rect 9766 20204 9772 20216
rect 9824 20244 9830 20256
rect 10594 20244 10600 20256
rect 9824 20216 10600 20244
rect 9824 20204 9830 20216
rect 10594 20204 10600 20216
rect 10652 20204 10658 20256
rect 10870 20244 10876 20256
rect 10831 20216 10876 20244
rect 10870 20204 10876 20216
rect 10928 20204 10934 20256
rect 12406 20244 12434 20284
rect 13262 20272 13268 20324
rect 13320 20272 13326 20324
rect 22112 20312 22140 20352
rect 15028 20284 22140 20312
rect 15028 20244 15056 20284
rect 22186 20272 22192 20324
rect 22244 20312 22250 20324
rect 23109 20315 23167 20321
rect 23109 20312 23121 20315
rect 22244 20284 23121 20312
rect 22244 20272 22250 20284
rect 23109 20281 23121 20284
rect 23155 20281 23167 20315
rect 23109 20275 23167 20281
rect 12406 20216 15056 20244
rect 15105 20247 15163 20253
rect 15105 20213 15117 20247
rect 15151 20244 15163 20247
rect 16666 20244 16672 20256
rect 15151 20216 16672 20244
rect 15151 20213 15163 20216
rect 15105 20207 15163 20213
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 16945 20247 17003 20253
rect 16945 20244 16957 20247
rect 16816 20216 16957 20244
rect 16816 20204 16822 20216
rect 16945 20213 16957 20216
rect 16991 20213 17003 20247
rect 16945 20207 17003 20213
rect 19153 20247 19211 20253
rect 19153 20213 19165 20247
rect 19199 20244 19211 20247
rect 20530 20244 20536 20256
rect 19199 20216 20536 20244
rect 19199 20213 19211 20216
rect 19153 20207 19211 20213
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 23216 20244 23244 20352
rect 23474 20340 23480 20392
rect 23532 20380 23538 20392
rect 23661 20383 23719 20389
rect 23661 20380 23673 20383
rect 23532 20352 23673 20380
rect 23532 20340 23538 20352
rect 23661 20349 23673 20352
rect 23707 20349 23719 20383
rect 24026 20380 24032 20392
rect 23987 20352 24032 20380
rect 23661 20343 23719 20349
rect 24026 20340 24032 20352
rect 24084 20340 24090 20392
rect 25685 20383 25743 20389
rect 25685 20349 25697 20383
rect 25731 20380 25743 20383
rect 26142 20380 26148 20392
rect 25731 20352 26148 20380
rect 25731 20349 25743 20352
rect 25685 20343 25743 20349
rect 26142 20340 26148 20352
rect 26200 20380 26206 20392
rect 27264 20380 27292 20488
rect 28261 20485 28273 20519
rect 28307 20516 28319 20519
rect 29641 20519 29699 20525
rect 29641 20516 29653 20519
rect 28307 20488 29653 20516
rect 28307 20485 28319 20488
rect 28261 20479 28319 20485
rect 29641 20485 29653 20488
rect 29687 20485 29699 20519
rect 29641 20479 29699 20485
rect 27338 20408 27344 20460
rect 27396 20448 27402 20460
rect 28169 20451 28227 20457
rect 28169 20448 28181 20451
rect 27396 20420 28181 20448
rect 27396 20408 27402 20420
rect 28169 20417 28181 20420
rect 28215 20417 28227 20451
rect 28994 20448 29000 20460
rect 28907 20420 29000 20448
rect 28169 20411 28227 20417
rect 28966 20408 29000 20420
rect 29052 20408 29058 20460
rect 26200 20352 27292 20380
rect 26200 20340 26206 20352
rect 26237 20315 26295 20321
rect 26237 20281 26249 20315
rect 26283 20312 26295 20315
rect 26418 20312 26424 20324
rect 26283 20284 26424 20312
rect 26283 20281 26295 20284
rect 26237 20275 26295 20281
rect 26418 20272 26424 20284
rect 26476 20272 26482 20324
rect 28966 20312 28994 20408
rect 29546 20380 29552 20392
rect 29507 20352 29552 20380
rect 29546 20340 29552 20352
rect 29604 20340 29610 20392
rect 30374 20380 30380 20392
rect 30335 20352 30380 20380
rect 30374 20340 30380 20352
rect 30432 20340 30438 20392
rect 26528 20284 28994 20312
rect 26528 20244 26556 20284
rect 22152 20216 22197 20244
rect 23216 20216 26556 20244
rect 28813 20247 28871 20253
rect 22152 20204 22158 20216
rect 28813 20213 28825 20247
rect 28859 20244 28871 20247
rect 29730 20244 29736 20256
rect 28859 20216 29736 20244
rect 28859 20213 28871 20216
rect 28813 20207 28871 20213
rect 29730 20204 29736 20216
rect 29788 20204 29794 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 2130 20000 2136 20052
rect 2188 20040 2194 20052
rect 2188 20012 7696 20040
rect 2188 20000 2194 20012
rect 5718 19972 5724 19984
rect 5679 19944 5724 19972
rect 5718 19932 5724 19944
rect 5776 19932 5782 19984
rect 1673 19907 1731 19913
rect 1673 19873 1685 19907
rect 1719 19904 1731 19907
rect 3142 19904 3148 19916
rect 1719 19876 3148 19904
rect 1719 19873 1731 19876
rect 1673 19867 1731 19873
rect 3142 19864 3148 19876
rect 3200 19904 3206 19916
rect 3970 19904 3976 19916
rect 3200 19876 3976 19904
rect 3200 19864 3206 19876
rect 3970 19864 3976 19876
rect 4028 19864 4034 19916
rect 4249 19907 4307 19913
rect 4249 19873 4261 19907
rect 4295 19904 4307 19907
rect 5534 19904 5540 19916
rect 4295 19876 5540 19904
rect 4295 19873 4307 19876
rect 4249 19867 4307 19873
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 6549 19907 6607 19913
rect 6549 19873 6561 19907
rect 6595 19904 6607 19907
rect 7006 19904 7012 19916
rect 6595 19876 7012 19904
rect 6595 19873 6607 19876
rect 6549 19867 6607 19873
rect 7006 19864 7012 19876
rect 7064 19864 7070 19916
rect 6273 19839 6331 19845
rect 6273 19805 6285 19839
rect 6319 19805 6331 19839
rect 7668 19822 7696 20012
rect 7742 20000 7748 20052
rect 7800 20040 7806 20052
rect 10686 20040 10692 20052
rect 7800 20012 10692 20040
rect 7800 20000 7806 20012
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 10860 20043 10918 20049
rect 10860 20009 10872 20043
rect 10906 20040 10918 20043
rect 15286 20040 15292 20052
rect 10906 20012 15292 20040
rect 10906 20009 10918 20012
rect 10860 20003 10918 20009
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 28258 20040 28264 20052
rect 15383 20012 28264 20040
rect 12250 19932 12256 19984
rect 12308 19972 12314 19984
rect 12345 19975 12403 19981
rect 12345 19972 12357 19975
rect 12308 19944 12357 19972
rect 12308 19932 12314 19944
rect 12345 19941 12357 19944
rect 12391 19941 12403 19975
rect 12345 19935 12403 19941
rect 10594 19904 10600 19916
rect 10507 19876 10600 19904
rect 10594 19864 10600 19876
rect 10652 19904 10658 19916
rect 10962 19904 10968 19916
rect 10652 19876 10968 19904
rect 10652 19864 10658 19876
rect 10962 19864 10968 19876
rect 11020 19864 11026 19916
rect 11882 19864 11888 19916
rect 11940 19904 11946 19916
rect 13004 19904 13216 19920
rect 15102 19904 15108 19916
rect 11940 19892 15108 19904
rect 11940 19876 13032 19892
rect 13188 19876 15108 19892
rect 11940 19864 11946 19876
rect 12912 19845 12940 19876
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 12897 19839 12955 19845
rect 6273 19799 6331 19805
rect 12897 19805 12909 19839
rect 12943 19805 12955 19839
rect 15383 19836 15411 20012
rect 28258 20000 28264 20012
rect 28316 20000 28322 20052
rect 21634 19932 21640 19984
rect 21692 19932 21698 19984
rect 22646 19932 22652 19984
rect 22704 19972 22710 19984
rect 24026 19972 24032 19984
rect 22704 19944 24032 19972
rect 22704 19932 22710 19944
rect 24026 19932 24032 19944
rect 24084 19972 24090 19984
rect 28902 19972 28908 19984
rect 24084 19944 28908 19972
rect 24084 19932 24090 19944
rect 28902 19932 28908 19944
rect 28960 19932 28966 19984
rect 16574 19904 16580 19916
rect 16535 19876 16580 19904
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 16942 19864 16948 19916
rect 17000 19904 17006 19916
rect 20254 19904 20260 19916
rect 17000 19876 20260 19904
rect 17000 19864 17006 19876
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 20530 19904 20536 19916
rect 20491 19876 20536 19904
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 20898 19904 20904 19916
rect 20859 19876 20904 19904
rect 20898 19864 20904 19876
rect 20956 19904 20962 19916
rect 21652 19904 21680 19932
rect 20956 19876 21680 19904
rect 23753 19907 23811 19913
rect 20956 19864 20962 19876
rect 23753 19873 23765 19907
rect 23799 19904 23811 19907
rect 25682 19904 25688 19916
rect 23799 19876 25688 19904
rect 23799 19873 23811 19876
rect 23753 19867 23811 19873
rect 25682 19864 25688 19876
rect 25740 19864 25746 19916
rect 26142 19904 26148 19916
rect 26103 19876 26148 19904
rect 26142 19864 26148 19876
rect 26200 19864 26206 19916
rect 26602 19904 26608 19916
rect 26563 19876 26608 19904
rect 26602 19864 26608 19876
rect 26660 19864 26666 19916
rect 20346 19836 20352 19848
rect 12897 19799 12955 19805
rect 13004 19808 15411 19836
rect 20307 19808 20352 19836
rect 1949 19771 2007 19777
rect 1949 19737 1961 19771
rect 1995 19737 2007 19771
rect 3234 19768 3240 19780
rect 3174 19740 3240 19768
rect 1949 19731 2007 19737
rect 1964 19700 1992 19731
rect 3234 19728 3240 19740
rect 3292 19728 3298 19780
rect 3326 19728 3332 19780
rect 3384 19768 3390 19780
rect 3384 19740 3740 19768
rect 3384 19728 3390 19740
rect 3344 19700 3372 19728
rect 1964 19672 3372 19700
rect 3421 19703 3479 19709
rect 3421 19669 3433 19703
rect 3467 19700 3479 19703
rect 3602 19700 3608 19712
rect 3467 19672 3608 19700
rect 3467 19669 3479 19672
rect 3421 19663 3479 19669
rect 3602 19660 3608 19672
rect 3660 19660 3666 19712
rect 3712 19700 3740 19740
rect 4706 19728 4712 19780
rect 4764 19728 4770 19780
rect 5166 19700 5172 19712
rect 3712 19672 5172 19700
rect 5166 19660 5172 19672
rect 5224 19660 5230 19712
rect 6288 19700 6316 19799
rect 11330 19728 11336 19780
rect 11388 19728 11394 19780
rect 12250 19728 12256 19780
rect 12308 19768 12314 19780
rect 13004 19768 13032 19808
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 24946 19836 24952 19848
rect 24907 19808 24952 19836
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 27430 19796 27436 19848
rect 27488 19836 27494 19848
rect 28353 19839 28411 19845
rect 28353 19836 28365 19839
rect 27488 19808 28365 19836
rect 27488 19796 27494 19808
rect 28353 19805 28365 19808
rect 28399 19805 28411 19839
rect 28353 19799 28411 19805
rect 28442 19796 28448 19848
rect 28500 19836 28506 19848
rect 28997 19839 29055 19845
rect 28997 19836 29009 19839
rect 28500 19808 29009 19836
rect 28500 19796 28506 19808
rect 28997 19805 29009 19808
rect 29043 19805 29055 19839
rect 28997 19799 29055 19805
rect 12308 19740 13032 19768
rect 12308 19728 12314 19740
rect 13170 19728 13176 19780
rect 13228 19768 13234 19780
rect 16482 19768 16488 19780
rect 13228 19740 16488 19768
rect 13228 19728 13234 19740
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 16853 19771 16911 19777
rect 16853 19737 16865 19771
rect 16899 19768 16911 19771
rect 16942 19768 16948 19780
rect 16899 19740 16948 19768
rect 16899 19737 16911 19740
rect 16853 19731 16911 19737
rect 16942 19728 16948 19740
rect 17000 19728 17006 19780
rect 19426 19768 19432 19780
rect 18078 19740 19432 19768
rect 19426 19728 19432 19740
rect 19484 19728 19490 19780
rect 22738 19768 22744 19780
rect 22699 19740 22744 19768
rect 22738 19728 22744 19740
rect 22796 19728 22802 19780
rect 22830 19728 22836 19780
rect 22888 19768 22894 19780
rect 22888 19740 22933 19768
rect 24872 19740 26188 19768
rect 22888 19728 22894 19740
rect 6822 19700 6828 19712
rect 6288 19672 6828 19700
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 7834 19660 7840 19712
rect 7892 19700 7898 19712
rect 8021 19703 8079 19709
rect 8021 19700 8033 19703
rect 7892 19672 8033 19700
rect 7892 19660 7898 19672
rect 8021 19669 8033 19672
rect 8067 19669 8079 19703
rect 8021 19663 8079 19669
rect 13722 19660 13728 19712
rect 13780 19700 13786 19712
rect 17126 19700 17132 19712
rect 13780 19672 17132 19700
rect 13780 19660 13786 19672
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 18322 19700 18328 19712
rect 18283 19672 18328 19700
rect 18322 19660 18328 19672
rect 18380 19700 18386 19712
rect 24872 19700 24900 19740
rect 25038 19700 25044 19712
rect 18380 19672 24900 19700
rect 24999 19672 25044 19700
rect 18380 19660 18386 19672
rect 25038 19660 25044 19672
rect 25096 19660 25102 19712
rect 26160 19700 26188 19740
rect 26234 19728 26240 19780
rect 26292 19768 26298 19780
rect 27709 19771 27767 19777
rect 26292 19740 26337 19768
rect 26292 19728 26298 19740
rect 27709 19737 27721 19771
rect 27755 19768 27767 19771
rect 29638 19768 29644 19780
rect 27755 19740 29644 19768
rect 27755 19737 27767 19740
rect 27709 19731 27767 19737
rect 29638 19728 29644 19740
rect 29696 19728 29702 19780
rect 27338 19700 27344 19712
rect 26160 19672 27344 19700
rect 27338 19660 27344 19672
rect 27396 19660 27402 19712
rect 27798 19700 27804 19712
rect 27759 19672 27804 19700
rect 27798 19660 27804 19672
rect 27856 19660 27862 19712
rect 28445 19703 28503 19709
rect 28445 19669 28457 19703
rect 28491 19700 28503 19703
rect 28994 19700 29000 19712
rect 28491 19672 29000 19700
rect 28491 19669 28503 19672
rect 28445 19663 28503 19669
rect 28994 19660 29000 19672
rect 29052 19660 29058 19712
rect 29089 19703 29147 19709
rect 29089 19669 29101 19703
rect 29135 19700 29147 19703
rect 30558 19700 30564 19712
rect 29135 19672 30564 19700
rect 29135 19669 29147 19672
rect 29089 19663 29147 19669
rect 30558 19660 30564 19672
rect 30616 19660 30622 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 3329 19499 3387 19505
rect 3329 19465 3341 19499
rect 3375 19496 3387 19499
rect 3694 19496 3700 19508
rect 3375 19468 3700 19496
rect 3375 19465 3387 19468
rect 3329 19459 3387 19465
rect 3694 19456 3700 19468
rect 3752 19456 3758 19508
rect 4890 19456 4896 19508
rect 4948 19496 4954 19508
rect 5997 19499 6055 19505
rect 4948 19468 5856 19496
rect 4948 19456 4954 19468
rect 2866 19388 2872 19440
rect 2924 19388 2930 19440
rect 5828 19428 5856 19468
rect 5997 19465 6009 19499
rect 6043 19496 6055 19499
rect 7466 19496 7472 19508
rect 6043 19468 7472 19496
rect 6043 19465 6055 19468
rect 5997 19459 6055 19465
rect 7466 19456 7472 19468
rect 7524 19456 7530 19508
rect 9766 19496 9772 19508
rect 8220 19468 9772 19496
rect 5828 19400 8156 19428
rect 3970 19320 3976 19372
rect 4028 19360 4034 19372
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 4028 19332 4261 19360
rect 4028 19320 4034 19332
rect 4249 19329 4261 19332
rect 4295 19329 4307 19363
rect 5810 19360 5816 19372
rect 5658 19332 5816 19360
rect 4249 19323 4307 19329
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 1581 19295 1639 19301
rect 1581 19261 1593 19295
rect 1627 19292 1639 19295
rect 1857 19295 1915 19301
rect 1627 19264 1716 19292
rect 1627 19261 1639 19264
rect 1581 19255 1639 19261
rect 1688 19168 1716 19264
rect 1857 19261 1869 19295
rect 1903 19292 1915 19295
rect 4525 19295 4583 19301
rect 1903 19264 4384 19292
rect 1903 19261 1915 19264
rect 1857 19255 1915 19261
rect 1670 19116 1676 19168
rect 1728 19116 1734 19168
rect 4356 19156 4384 19264
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 5994 19292 6000 19304
rect 4571 19264 6000 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 5994 19252 6000 19264
rect 6052 19292 6058 19304
rect 6454 19292 6460 19304
rect 6052 19264 6460 19292
rect 6052 19252 6058 19264
rect 6454 19252 6460 19264
rect 6512 19252 6518 19304
rect 8128 19292 8156 19400
rect 8220 19369 8248 19468
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 15841 19499 15899 19505
rect 15841 19465 15853 19499
rect 15887 19496 15899 19499
rect 16666 19496 16672 19508
rect 15887 19468 16672 19496
rect 15887 19465 15899 19468
rect 15841 19459 15899 19465
rect 16666 19456 16672 19468
rect 16724 19496 16730 19508
rect 18601 19499 18659 19505
rect 16724 19468 18460 19496
rect 16724 19456 16730 19468
rect 8938 19388 8944 19440
rect 8996 19388 9002 19440
rect 13630 19428 13636 19440
rect 13386 19400 13636 19428
rect 13630 19388 13636 19400
rect 13688 19388 13694 19440
rect 16758 19428 16764 19440
rect 15594 19400 16764 19428
rect 16758 19388 16764 19400
rect 16816 19388 16822 19440
rect 17770 19388 17776 19440
rect 17828 19388 17834 19440
rect 18432 19428 18460 19468
rect 18601 19465 18613 19499
rect 18647 19496 18659 19499
rect 19242 19496 19248 19508
rect 18647 19468 19248 19496
rect 18647 19465 18659 19468
rect 18601 19459 18659 19465
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 20346 19496 20352 19508
rect 20307 19468 20352 19496
rect 20346 19456 20352 19468
rect 20404 19456 20410 19508
rect 27430 19496 27436 19508
rect 20456 19468 27436 19496
rect 20456 19428 20484 19468
rect 27430 19456 27436 19468
rect 27488 19456 27494 19508
rect 30374 19496 30380 19508
rect 29932 19468 30380 19496
rect 18432 19400 20484 19428
rect 21085 19431 21143 19437
rect 21085 19397 21097 19431
rect 21131 19428 21143 19431
rect 22189 19431 22247 19437
rect 22189 19428 22201 19431
rect 21131 19400 22201 19428
rect 21131 19397 21143 19400
rect 21085 19391 21143 19397
rect 22189 19397 22201 19400
rect 22235 19397 22247 19431
rect 23106 19428 23112 19440
rect 23067 19400 23112 19428
rect 22189 19391 22247 19397
rect 23106 19388 23112 19400
rect 23164 19388 23170 19440
rect 24213 19431 24271 19437
rect 24213 19397 24225 19431
rect 24259 19428 24271 19431
rect 24762 19428 24768 19440
rect 24259 19400 24768 19428
rect 24259 19397 24271 19400
rect 24213 19391 24271 19397
rect 24762 19388 24768 19400
rect 24820 19388 24826 19440
rect 28994 19428 29000 19440
rect 28955 19400 29000 19428
rect 28994 19388 29000 19400
rect 29052 19388 29058 19440
rect 29932 19437 29960 19468
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 37642 19456 37648 19508
rect 37700 19496 37706 19508
rect 38105 19499 38163 19505
rect 38105 19496 38117 19499
rect 37700 19468 38117 19496
rect 37700 19456 37706 19468
rect 38105 19465 38117 19468
rect 38151 19465 38163 19499
rect 38105 19459 38163 19465
rect 29917 19431 29975 19437
rect 29917 19397 29929 19431
rect 29963 19397 29975 19431
rect 30558 19428 30564 19440
rect 30519 19400 30564 19428
rect 29917 19391 29975 19397
rect 30558 19388 30564 19400
rect 30616 19388 30622 19440
rect 8205 19363 8263 19369
rect 8205 19329 8217 19363
rect 8251 19329 8263 19363
rect 13722 19360 13728 19372
rect 8205 19323 8263 19329
rect 13648 19332 13728 19360
rect 8481 19295 8539 19301
rect 8128 19264 8248 19292
rect 5994 19156 6000 19168
rect 4356 19128 6000 19156
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 8220 19156 8248 19264
rect 8481 19261 8493 19295
rect 8527 19292 8539 19295
rect 8527 19264 10456 19292
rect 8527 19261 8539 19264
rect 8481 19255 8539 19261
rect 9953 19159 10011 19165
rect 9953 19156 9965 19159
rect 8220 19128 9965 19156
rect 9953 19125 9965 19128
rect 9999 19125 10011 19159
rect 10428 19156 10456 19264
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11885 19295 11943 19301
rect 11885 19292 11897 19295
rect 11112 19264 11897 19292
rect 11112 19252 11118 19264
rect 11885 19261 11897 19264
rect 11931 19261 11943 19295
rect 12158 19292 12164 19304
rect 12119 19264 12164 19292
rect 11885 19255 11943 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 13648 19301 13676 19332
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 14090 19360 14096 19372
rect 14051 19332 14096 19360
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16632 19332 16865 19360
rect 16632 19320 16638 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 18874 19320 18880 19372
rect 18932 19360 18938 19372
rect 18932 19332 20208 19360
rect 18932 19320 18938 19332
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19292 13691 19295
rect 14369 19295 14427 19301
rect 13679 19264 13713 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 14369 19261 14381 19295
rect 14415 19292 14427 19295
rect 14415 19264 16988 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 13814 19156 13820 19168
rect 10428 19128 13820 19156
rect 9953 19119 10011 19125
rect 13814 19116 13820 19128
rect 13872 19156 13878 19168
rect 14366 19156 14372 19168
rect 13872 19128 14372 19156
rect 13872 19116 13878 19128
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 16960 19156 16988 19264
rect 17126 19252 17132 19304
rect 17184 19292 17190 19304
rect 18690 19292 18696 19304
rect 17184 19264 18696 19292
rect 17184 19252 17190 19264
rect 18690 19252 18696 19264
rect 18748 19252 18754 19304
rect 20180 19292 20208 19332
rect 20254 19320 20260 19372
rect 20312 19360 20318 19372
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 20312 19332 21005 19360
rect 20312 19320 20318 19332
rect 20993 19329 21005 19332
rect 21039 19329 21051 19363
rect 23569 19363 23627 19369
rect 20993 19323 21051 19329
rect 21100 19332 21956 19360
rect 21100 19292 21128 19332
rect 20180 19264 21128 19292
rect 21928 19292 21956 19332
rect 23569 19329 23581 19363
rect 23615 19360 23627 19363
rect 23842 19360 23848 19372
rect 23615 19332 23848 19360
rect 23615 19329 23627 19332
rect 23569 19323 23627 19329
rect 23842 19320 23848 19332
rect 23900 19320 23906 19372
rect 24026 19320 24032 19372
rect 24084 19360 24090 19372
rect 24857 19363 24915 19369
rect 24857 19360 24869 19363
rect 24084 19332 24869 19360
rect 24084 19320 24090 19332
rect 24857 19329 24869 19332
rect 24903 19329 24915 19363
rect 24857 19323 24915 19329
rect 28074 19320 28080 19372
rect 28132 19360 28138 19372
rect 38286 19360 38292 19372
rect 28132 19332 28764 19360
rect 38247 19332 38292 19360
rect 28132 19320 28138 19332
rect 22097 19295 22155 19301
rect 22097 19292 22109 19295
rect 21928 19264 22109 19292
rect 22097 19261 22109 19264
rect 22143 19261 22155 19295
rect 22097 19255 22155 19261
rect 23753 19295 23811 19301
rect 23753 19261 23765 19295
rect 23799 19261 23811 19295
rect 28736 19292 28764 19332
rect 38286 19320 38292 19332
rect 38344 19320 38350 19372
rect 28902 19292 28908 19304
rect 28736 19264 28908 19292
rect 23753 19255 23811 19261
rect 23768 19224 23796 19255
rect 28902 19252 28908 19264
rect 28960 19252 28966 19304
rect 30466 19292 30472 19304
rect 30427 19264 30472 19292
rect 30466 19252 30472 19264
rect 30524 19252 30530 19304
rect 30745 19295 30803 19301
rect 30745 19261 30757 19295
rect 30791 19261 30803 19295
rect 30745 19255 30803 19261
rect 24673 19227 24731 19233
rect 24673 19224 24685 19227
rect 23768 19196 24685 19224
rect 24673 19193 24685 19196
rect 24719 19193 24731 19227
rect 24673 19187 24731 19193
rect 28810 19184 28816 19236
rect 28868 19224 28874 19236
rect 30760 19224 30788 19255
rect 28868 19196 30788 19224
rect 28868 19184 28874 19196
rect 18322 19156 18328 19168
rect 16960 19128 18328 19156
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 22462 19116 22468 19168
rect 22520 19156 22526 19168
rect 30098 19156 30104 19168
rect 22520 19128 30104 19156
rect 22520 19116 22526 19128
rect 30098 19116 30104 19128
rect 30156 19116 30162 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 6546 18912 6552 18964
rect 6604 18952 6610 18964
rect 9950 18952 9956 18964
rect 6604 18924 9956 18952
rect 6604 18912 6610 18924
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 10100 18924 12434 18952
rect 10100 18912 10106 18924
rect 12406 18884 12434 18924
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 12805 18955 12863 18961
rect 12805 18952 12817 18955
rect 12584 18924 12817 18952
rect 12584 18912 12590 18924
rect 12805 18921 12817 18924
rect 12851 18952 12863 18955
rect 13538 18952 13544 18964
rect 12851 18924 13544 18952
rect 12851 18921 12863 18924
rect 12805 18915 12863 18921
rect 13538 18912 13544 18924
rect 13596 18912 13602 18964
rect 15010 18912 15016 18964
rect 15068 18952 15074 18964
rect 15068 18924 16068 18952
rect 15068 18912 15074 18924
rect 16040 18884 16068 18924
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 19484 18924 19533 18952
rect 19484 18912 19490 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 22738 18952 22744 18964
rect 22699 18924 22744 18952
rect 19521 18915 19579 18921
rect 22738 18912 22744 18924
rect 22796 18912 22802 18964
rect 23106 18912 23112 18964
rect 23164 18952 23170 18964
rect 30098 18952 30104 18964
rect 23164 18924 24072 18952
rect 30059 18924 30104 18952
rect 23164 18912 23170 18924
rect 12406 18856 14872 18884
rect 16040 18856 23244 18884
rect 1949 18819 2007 18825
rect 1949 18785 1961 18819
rect 1995 18816 2007 18819
rect 3418 18816 3424 18828
rect 1995 18788 3424 18816
rect 1995 18785 2007 18788
rect 1949 18779 2007 18785
rect 3418 18776 3424 18788
rect 3476 18776 3482 18828
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18816 4675 18819
rect 7101 18819 7159 18825
rect 4663 18788 6868 18816
rect 4663 18785 4675 18788
rect 4617 18779 4675 18785
rect 6840 18760 6868 18788
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 8573 18819 8631 18825
rect 7147 18788 8524 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 1670 18748 1676 18760
rect 1631 18720 1676 18748
rect 1670 18708 1676 18720
rect 1728 18708 1734 18760
rect 3050 18708 3056 18760
rect 3108 18708 3114 18760
rect 6822 18748 6828 18760
rect 6783 18720 6828 18748
rect 6822 18708 6828 18720
rect 6880 18708 6886 18760
rect 8202 18708 8208 18760
rect 8260 18708 8266 18760
rect 8496 18748 8524 18788
rect 8573 18785 8585 18819
rect 8619 18816 8631 18819
rect 11330 18816 11336 18828
rect 8619 18788 11336 18816
rect 8619 18785 8631 18788
rect 8573 18779 8631 18785
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14737 18819 14795 18825
rect 14737 18816 14749 18819
rect 14148 18788 14749 18816
rect 14148 18776 14154 18788
rect 14737 18785 14749 18788
rect 14783 18785 14795 18819
rect 14844 18816 14872 18856
rect 20806 18816 20812 18828
rect 14844 18788 20812 18816
rect 14737 18779 14795 18785
rect 20806 18776 20812 18788
rect 20864 18776 20870 18828
rect 8662 18748 8668 18760
rect 8496 18720 8668 18748
rect 8662 18708 8668 18720
rect 8720 18708 8726 18760
rect 11054 18748 11060 18760
rect 11015 18720 11060 18748
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 16390 18708 16396 18760
rect 16448 18748 16454 18760
rect 16761 18751 16819 18757
rect 16761 18748 16773 18751
rect 16448 18720 16773 18748
rect 16448 18708 16454 18720
rect 16761 18717 16773 18720
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 4893 18683 4951 18689
rect 4893 18649 4905 18683
rect 4939 18649 4951 18683
rect 4893 18643 4951 18649
rect 3421 18615 3479 18621
rect 3421 18581 3433 18615
rect 3467 18612 3479 18615
rect 4614 18612 4620 18624
rect 3467 18584 4620 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 4614 18572 4620 18584
rect 4672 18572 4678 18624
rect 4908 18612 4936 18643
rect 5626 18640 5632 18692
rect 5684 18640 5690 18692
rect 11790 18640 11796 18692
rect 11848 18640 11854 18692
rect 15010 18680 15016 18692
rect 14971 18652 15016 18680
rect 15010 18640 15016 18652
rect 15068 18640 15074 18692
rect 15102 18640 15108 18692
rect 15160 18680 15166 18692
rect 16776 18680 16804 18711
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 19392 18720 19441 18748
rect 19392 18708 19398 18720
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 23216 18757 23244 18856
rect 23937 18819 23995 18825
rect 23937 18816 23949 18819
rect 23308 18788 23949 18816
rect 22097 18751 22155 18757
rect 22097 18748 22109 18751
rect 20036 18720 22109 18748
rect 20036 18708 20042 18720
rect 22097 18717 22109 18720
rect 22143 18717 22155 18751
rect 22097 18711 22155 18717
rect 22281 18751 22339 18757
rect 22281 18717 22293 18751
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 23201 18751 23259 18757
rect 23201 18717 23213 18751
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 21634 18680 21640 18692
rect 15160 18652 15502 18680
rect 16776 18652 21640 18680
rect 15160 18640 15166 18652
rect 21634 18640 21640 18652
rect 21692 18640 21698 18692
rect 22296 18680 22324 18711
rect 23308 18680 23336 18788
rect 23937 18785 23949 18788
rect 23983 18785 23995 18819
rect 23937 18779 23995 18785
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18717 23903 18751
rect 23845 18711 23903 18717
rect 22296 18652 23336 18680
rect 5258 18612 5264 18624
rect 4908 18584 5264 18612
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 6362 18612 6368 18624
rect 5592 18584 6368 18612
rect 5592 18572 5598 18584
rect 6362 18572 6368 18584
rect 6420 18572 6426 18624
rect 6454 18572 6460 18624
rect 6512 18612 6518 18624
rect 9858 18612 9864 18624
rect 6512 18584 9864 18612
rect 6512 18572 6518 18584
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 13538 18572 13544 18624
rect 13596 18612 13602 18624
rect 18506 18612 18512 18624
rect 13596 18584 18512 18612
rect 13596 18572 13602 18584
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 22922 18572 22928 18624
rect 22980 18612 22986 18624
rect 23293 18615 23351 18621
rect 23293 18612 23305 18615
rect 22980 18584 23305 18612
rect 22980 18572 22986 18584
rect 23293 18581 23305 18584
rect 23339 18581 23351 18615
rect 23860 18612 23888 18711
rect 24044 18680 24072 18924
rect 30098 18912 30104 18924
rect 30156 18912 30162 18964
rect 25222 18884 25228 18896
rect 25183 18856 25228 18884
rect 25222 18844 25228 18856
rect 25280 18844 25286 18896
rect 24673 18819 24731 18825
rect 24673 18785 24685 18819
rect 24719 18816 24731 18819
rect 25777 18819 25835 18825
rect 25777 18816 25789 18819
rect 24719 18788 25789 18816
rect 24719 18785 24731 18788
rect 24673 18779 24731 18785
rect 25777 18785 25789 18788
rect 25823 18785 25835 18819
rect 25777 18779 25835 18785
rect 30009 18751 30067 18757
rect 30009 18717 30021 18751
rect 30055 18748 30067 18751
rect 37918 18748 37924 18760
rect 30055 18720 37924 18748
rect 30055 18717 30067 18720
rect 30009 18711 30067 18717
rect 37918 18708 37924 18720
rect 37976 18708 37982 18760
rect 24765 18683 24823 18689
rect 24765 18680 24777 18683
rect 24044 18652 24777 18680
rect 24765 18649 24777 18652
rect 24811 18649 24823 18683
rect 24765 18643 24823 18649
rect 25130 18612 25136 18624
rect 23860 18584 25136 18612
rect 23293 18575 23351 18581
rect 25130 18572 25136 18584
rect 25188 18572 25194 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 3970 18408 3976 18420
rect 1728 18380 3976 18408
rect 1728 18368 1734 18380
rect 2056 18281 2084 18380
rect 3970 18368 3976 18380
rect 4028 18368 4034 18420
rect 5258 18368 5264 18420
rect 5316 18408 5322 18420
rect 5994 18408 6000 18420
rect 5316 18380 5856 18408
rect 5955 18380 6000 18408
rect 5316 18368 5322 18380
rect 3326 18300 3332 18352
rect 3384 18300 3390 18352
rect 3694 18300 3700 18352
rect 3752 18340 3758 18352
rect 3752 18312 5014 18340
rect 3752 18300 3758 18312
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 3970 18232 3976 18284
rect 4028 18272 4034 18284
rect 4249 18275 4307 18281
rect 4249 18272 4261 18275
rect 4028 18244 4261 18272
rect 4028 18232 4034 18244
rect 4249 18241 4261 18244
rect 4295 18241 4307 18275
rect 4249 18235 4307 18241
rect 2317 18207 2375 18213
rect 2317 18173 2329 18207
rect 2363 18204 2375 18207
rect 4154 18204 4160 18216
rect 2363 18176 4160 18204
rect 2363 18173 2375 18176
rect 2317 18167 2375 18173
rect 4154 18164 4160 18176
rect 4212 18164 4218 18216
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 4890 18204 4896 18216
rect 4571 18176 4896 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 4890 18164 4896 18176
rect 4948 18204 4954 18216
rect 5258 18204 5264 18216
rect 4948 18176 5264 18204
rect 4948 18164 4954 18176
rect 5258 18164 5264 18176
rect 5316 18164 5322 18216
rect 5828 18204 5856 18380
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 6641 18411 6699 18417
rect 6641 18377 6653 18411
rect 6687 18408 6699 18411
rect 8938 18408 8944 18420
rect 6687 18380 8944 18408
rect 6687 18377 6699 18380
rect 6641 18371 6699 18377
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 11698 18368 11704 18420
rect 11756 18408 11762 18420
rect 11793 18411 11851 18417
rect 11793 18408 11805 18411
rect 11756 18380 11805 18408
rect 11756 18368 11762 18380
rect 11793 18377 11805 18380
rect 11839 18377 11851 18411
rect 11793 18371 11851 18377
rect 13722 18368 13728 18420
rect 13780 18408 13786 18420
rect 15286 18408 15292 18420
rect 13780 18380 14228 18408
rect 15247 18380 15292 18408
rect 13780 18368 13786 18380
rect 7098 18300 7104 18352
rect 7156 18340 7162 18352
rect 7466 18340 7472 18352
rect 7156 18312 7472 18340
rect 7156 18300 7162 18312
rect 7466 18300 7472 18312
rect 7524 18300 7530 18352
rect 8294 18300 8300 18352
rect 8352 18300 8358 18352
rect 9950 18300 9956 18352
rect 10008 18340 10014 18352
rect 14090 18340 14096 18352
rect 10008 18312 11744 18340
rect 10008 18300 10014 18312
rect 6086 18232 6092 18284
rect 6144 18272 6150 18284
rect 6546 18272 6552 18284
rect 6144 18244 6552 18272
rect 6144 18232 6150 18244
rect 6546 18232 6552 18244
rect 6604 18232 6610 18284
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 11716 18281 11744 18312
rect 13556 18312 14096 18340
rect 11701 18275 11759 18281
rect 9272 18244 10180 18272
rect 9272 18232 9278 18244
rect 5828 18176 6776 18204
rect 6454 18136 6460 18148
rect 5644 18108 6460 18136
rect 3789 18071 3847 18077
rect 3789 18037 3801 18071
rect 3835 18068 3847 18071
rect 5644 18068 5672 18108
rect 6454 18096 6460 18108
rect 6512 18096 6518 18148
rect 3835 18040 5672 18068
rect 6748 18068 6776 18176
rect 6822 18164 6828 18216
rect 6880 18204 6886 18216
rect 7282 18204 7288 18216
rect 6880 18176 7288 18204
rect 6880 18164 6886 18176
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 7561 18207 7619 18213
rect 7561 18173 7573 18207
rect 7607 18204 7619 18207
rect 7650 18204 7656 18216
rect 7607 18176 7656 18204
rect 7607 18173 7619 18176
rect 7561 18167 7619 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 9309 18207 9367 18213
rect 9309 18173 9321 18207
rect 9355 18204 9367 18207
rect 10042 18204 10048 18216
rect 9355 18176 10048 18204
rect 9355 18173 9367 18176
rect 9309 18167 9367 18173
rect 10042 18164 10048 18176
rect 10100 18164 10106 18216
rect 10152 18204 10180 18244
rect 11701 18241 11713 18275
rect 11747 18272 11759 18275
rect 12618 18272 12624 18284
rect 11747 18244 12624 18272
rect 11747 18241 11759 18244
rect 11701 18235 11759 18241
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 13556 18281 13584 18312
rect 14090 18300 14096 18312
rect 14148 18300 14154 18352
rect 14200 18340 14228 18380
rect 15286 18368 15292 18380
rect 15344 18368 15350 18420
rect 18598 18408 18604 18420
rect 18559 18380 18604 18408
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 18966 18368 18972 18420
rect 19024 18408 19030 18420
rect 22649 18411 22707 18417
rect 19024 18380 20668 18408
rect 19024 18368 19030 18380
rect 17129 18343 17187 18349
rect 14200 18312 14306 18340
rect 17129 18309 17141 18343
rect 17175 18340 17187 18343
rect 17218 18340 17224 18352
rect 17175 18312 17224 18340
rect 17175 18309 17187 18312
rect 17129 18303 17187 18309
rect 17218 18300 17224 18312
rect 17276 18300 17282 18352
rect 18414 18340 18420 18352
rect 18354 18312 18420 18340
rect 18414 18300 18420 18312
rect 18472 18300 18478 18352
rect 18616 18340 18644 18368
rect 18616 18312 20576 18340
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 20548 18281 20576 18312
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16632 18244 16865 18272
rect 16632 18232 16638 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 19797 18275 19855 18281
rect 19797 18241 19809 18275
rect 19843 18241 19855 18275
rect 19797 18235 19855 18241
rect 20533 18275 20591 18281
rect 20533 18241 20545 18275
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 13814 18204 13820 18216
rect 10152 18176 13676 18204
rect 13775 18176 13820 18204
rect 11146 18068 11152 18080
rect 6748 18040 11152 18068
rect 3835 18037 3847 18040
rect 3789 18031 3847 18037
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 11330 18028 11336 18080
rect 11388 18068 11394 18080
rect 13538 18068 13544 18080
rect 11388 18040 13544 18068
rect 11388 18028 11394 18040
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 13648 18068 13676 18176
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 19812 18136 19840 18235
rect 20640 18204 20668 18380
rect 22649 18377 22661 18411
rect 22695 18408 22707 18411
rect 22738 18408 22744 18420
rect 22695 18380 22744 18408
rect 22695 18377 22707 18380
rect 22649 18371 22707 18377
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 23109 18411 23167 18417
rect 23109 18377 23121 18411
rect 23155 18408 23167 18411
rect 24026 18408 24032 18420
rect 23155 18380 24032 18408
rect 23155 18377 23167 18380
rect 23109 18371 23167 18377
rect 24026 18368 24032 18380
rect 24084 18368 24090 18420
rect 36630 18368 36636 18420
rect 36688 18408 36694 18420
rect 38105 18411 38163 18417
rect 38105 18408 38117 18411
rect 36688 18380 38117 18408
rect 36688 18368 36694 18380
rect 38105 18377 38117 18380
rect 38151 18377 38163 18411
rect 38105 18371 38163 18377
rect 20806 18300 20812 18352
rect 20864 18340 20870 18352
rect 21726 18340 21732 18352
rect 20864 18312 21732 18340
rect 20864 18300 20870 18312
rect 21726 18300 21732 18312
rect 21784 18340 21790 18352
rect 21784 18312 23336 18340
rect 21784 18300 21790 18312
rect 21910 18232 21916 18284
rect 21968 18272 21974 18284
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 21968 18244 22017 18272
rect 21968 18232 21974 18244
rect 22005 18241 22017 18244
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 23308 18281 23336 18312
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 22152 18244 22201 18272
rect 22152 18232 22158 18244
rect 22189 18241 22201 18244
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18241 23351 18275
rect 24486 18272 24492 18284
rect 24447 18244 24492 18272
rect 23293 18235 23351 18241
rect 24486 18232 24492 18244
rect 24544 18232 24550 18284
rect 38286 18272 38292 18284
rect 38247 18244 38292 18272
rect 38286 18232 38292 18244
rect 38344 18232 38350 18284
rect 24673 18207 24731 18213
rect 20640 18176 22094 18204
rect 14844 18108 15411 18136
rect 14844 18068 14872 18108
rect 13648 18040 14872 18068
rect 15383 18068 15411 18108
rect 18156 18108 19840 18136
rect 22066 18136 22094 18176
rect 24673 18173 24685 18207
rect 24719 18173 24731 18207
rect 24673 18167 24731 18173
rect 24688 18136 24716 18167
rect 22066 18108 24716 18136
rect 18156 18068 18184 18108
rect 15383 18040 18184 18068
rect 19794 18028 19800 18080
rect 19852 18068 19858 18080
rect 19889 18071 19947 18077
rect 19889 18068 19901 18071
rect 19852 18040 19901 18068
rect 19852 18028 19858 18040
rect 19889 18037 19901 18040
rect 19935 18037 19947 18071
rect 19889 18031 19947 18037
rect 20625 18071 20683 18077
rect 20625 18037 20637 18071
rect 20671 18068 20683 18071
rect 21358 18068 21364 18080
rect 20671 18040 21364 18068
rect 20671 18037 20683 18040
rect 20625 18031 20683 18037
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 4246 17824 4252 17876
rect 4304 17864 4310 17876
rect 4798 17864 4804 17876
rect 4304 17836 4804 17864
rect 4304 17824 4310 17836
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 5721 17867 5779 17873
rect 5721 17833 5733 17867
rect 5767 17864 5779 17867
rect 7006 17864 7012 17876
rect 5767 17836 7012 17864
rect 5767 17833 5779 17836
rect 5721 17827 5779 17833
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10778 17864 10784 17876
rect 9732 17836 10784 17864
rect 9732 17824 9738 17836
rect 10778 17824 10784 17836
rect 10836 17864 10842 17876
rect 11517 17867 11575 17873
rect 10836 17836 11100 17864
rect 10836 17824 10842 17836
rect 3970 17728 3976 17740
rect 3931 17700 3976 17728
rect 3970 17688 3976 17700
rect 4028 17688 4034 17740
rect 4249 17731 4307 17737
rect 4249 17697 4261 17731
rect 4295 17728 4307 17731
rect 4614 17728 4620 17740
rect 4295 17700 4620 17728
rect 4295 17697 4307 17700
rect 4249 17691 4307 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 6365 17731 6423 17737
rect 6365 17697 6377 17731
rect 6411 17728 6423 17731
rect 7282 17728 7288 17740
rect 6411 17700 7288 17728
rect 6411 17697 6423 17700
rect 6365 17691 6423 17697
rect 7282 17688 7288 17700
rect 7340 17728 7346 17740
rect 9769 17731 9827 17737
rect 9769 17728 9781 17731
rect 7340 17700 9781 17728
rect 7340 17688 7346 17700
rect 9769 17697 9781 17700
rect 9815 17697 9827 17731
rect 10042 17728 10048 17740
rect 10003 17700 10048 17728
rect 9769 17691 9827 17697
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 11072 17728 11100 17836
rect 11517 17833 11529 17867
rect 11563 17864 11575 17867
rect 15010 17864 15016 17876
rect 11563 17836 15016 17864
rect 11563 17833 11575 17836
rect 11517 17827 11575 17833
rect 15010 17824 15016 17836
rect 15068 17824 15074 17876
rect 17034 17864 17040 17876
rect 15120 17836 17040 17864
rect 12253 17731 12311 17737
rect 12253 17728 12265 17731
rect 11072 17700 12265 17728
rect 12253 17697 12265 17700
rect 12299 17697 12311 17731
rect 12253 17691 12311 17697
rect 1762 17660 1768 17672
rect 1723 17632 1768 17660
rect 1762 17620 1768 17632
rect 1820 17620 1826 17672
rect 2222 17660 2228 17672
rect 2183 17632 2228 17660
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 11974 17660 11980 17672
rect 11935 17632 11980 17660
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 1596 17564 4292 17592
rect 1596 17533 1624 17564
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17493 1639 17527
rect 1581 17487 1639 17493
rect 1762 17484 1768 17536
rect 1820 17524 1826 17536
rect 2038 17524 2044 17536
rect 1820 17496 2044 17524
rect 1820 17484 1826 17496
rect 2038 17484 2044 17496
rect 2096 17484 2102 17536
rect 2317 17527 2375 17533
rect 2317 17493 2329 17527
rect 2363 17524 2375 17527
rect 4154 17524 4160 17536
rect 2363 17496 4160 17524
rect 2363 17493 2375 17496
rect 2317 17487 2375 17493
rect 4154 17484 4160 17496
rect 4212 17484 4218 17536
rect 4264 17524 4292 17564
rect 4890 17552 4896 17604
rect 4948 17552 4954 17604
rect 5810 17592 5816 17604
rect 5552 17564 5816 17592
rect 5552 17524 5580 17564
rect 5810 17552 5816 17564
rect 5868 17552 5874 17604
rect 6641 17595 6699 17601
rect 6641 17561 6653 17595
rect 6687 17561 6699 17595
rect 6641 17555 6699 17561
rect 4264 17496 5580 17524
rect 6454 17484 6460 17536
rect 6512 17524 6518 17536
rect 6656 17524 6684 17555
rect 7098 17552 7104 17604
rect 7156 17552 7162 17604
rect 10502 17552 10508 17604
rect 10560 17552 10566 17604
rect 12710 17552 12716 17604
rect 12768 17552 12774 17604
rect 15120 17592 15148 17836
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 22557 17867 22615 17873
rect 22557 17833 22569 17867
rect 22603 17864 22615 17867
rect 22738 17864 22744 17876
rect 22603 17836 22744 17864
rect 22603 17833 22615 17836
rect 22557 17827 22615 17833
rect 22738 17824 22744 17836
rect 22796 17824 22802 17876
rect 17586 17756 17592 17808
rect 17644 17796 17650 17808
rect 24854 17796 24860 17808
rect 17644 17768 24860 17796
rect 17644 17756 17650 17768
rect 24854 17756 24860 17768
rect 24912 17756 24918 17808
rect 16301 17731 16359 17737
rect 16301 17697 16313 17731
rect 16347 17728 16359 17731
rect 16574 17728 16580 17740
rect 16347 17700 16580 17728
rect 16347 17697 16359 17700
rect 16301 17691 16359 17697
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 19794 17728 19800 17740
rect 19755 17700 19800 17728
rect 19794 17688 19800 17700
rect 19852 17688 19858 17740
rect 20806 17728 20812 17740
rect 20767 17700 20812 17728
rect 20806 17688 20812 17700
rect 20864 17688 20870 17740
rect 21358 17688 21364 17740
rect 21416 17728 21422 17740
rect 22097 17731 22155 17737
rect 22097 17728 22109 17731
rect 21416 17700 22109 17728
rect 21416 17688 21422 17700
rect 22097 17697 22109 17700
rect 22143 17697 22155 17731
rect 22097 17691 22155 17697
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 18104 17632 18521 17660
rect 18104 17620 18110 17632
rect 18509 17629 18521 17632
rect 18555 17660 18567 17663
rect 19334 17660 19340 17672
rect 18555 17632 19340 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 19334 17620 19340 17632
rect 19392 17620 19398 17672
rect 19426 17620 19432 17672
rect 19484 17660 19490 17672
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 19484 17632 19625 17660
rect 19484 17620 19490 17632
rect 19613 17629 19625 17632
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 21913 17663 21971 17669
rect 21913 17629 21925 17663
rect 21959 17660 21971 17663
rect 23014 17660 23020 17672
rect 21959 17632 23020 17660
rect 21959 17629 21971 17632
rect 21913 17623 21971 17629
rect 23014 17620 23020 17632
rect 23072 17620 23078 17672
rect 13648 17564 15148 17592
rect 16577 17595 16635 17601
rect 6512 17496 6684 17524
rect 6512 17484 6518 17496
rect 7558 17484 7564 17536
rect 7616 17524 7622 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7616 17496 8125 17524
rect 7616 17484 7622 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8113 17487 8171 17493
rect 10686 17484 10692 17536
rect 10744 17524 10750 17536
rect 13648 17524 13676 17564
rect 16577 17561 16589 17595
rect 16623 17592 16635 17595
rect 16666 17592 16672 17604
rect 16623 17564 16672 17592
rect 16623 17561 16635 17564
rect 16577 17555 16635 17561
rect 16666 17552 16672 17564
rect 16724 17552 16730 17604
rect 18601 17595 18659 17601
rect 18601 17592 18613 17595
rect 17802 17564 18613 17592
rect 18601 17561 18613 17564
rect 18647 17561 18659 17595
rect 18601 17555 18659 17561
rect 20806 17552 20812 17604
rect 20864 17592 20870 17604
rect 24026 17592 24032 17604
rect 20864 17564 24032 17592
rect 20864 17552 20870 17564
rect 24026 17552 24032 17564
rect 24084 17592 24090 17604
rect 37274 17592 37280 17604
rect 24084 17564 37280 17592
rect 24084 17552 24090 17564
rect 37274 17552 37280 17564
rect 37332 17552 37338 17604
rect 10744 17496 13676 17524
rect 13725 17527 13783 17533
rect 10744 17484 10750 17496
rect 13725 17493 13737 17527
rect 13771 17524 13783 17527
rect 13814 17524 13820 17536
rect 13771 17496 13820 17524
rect 13771 17493 13783 17496
rect 13725 17487 13783 17493
rect 13814 17484 13820 17496
rect 13872 17524 13878 17536
rect 14826 17524 14832 17536
rect 13872 17496 14832 17524
rect 13872 17484 13878 17496
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 15194 17484 15200 17536
rect 15252 17524 15258 17536
rect 18049 17527 18107 17533
rect 18049 17524 18061 17527
rect 15252 17496 18061 17524
rect 15252 17484 15258 17496
rect 18049 17493 18061 17496
rect 18095 17493 18107 17527
rect 18049 17487 18107 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1578 17280 1584 17332
rect 1636 17320 1642 17332
rect 2317 17323 2375 17329
rect 2317 17320 2329 17323
rect 1636 17292 2329 17320
rect 1636 17280 1642 17292
rect 2317 17289 2329 17292
rect 2363 17289 2375 17323
rect 2317 17283 2375 17289
rect 3145 17323 3203 17329
rect 3145 17289 3157 17323
rect 3191 17320 3203 17323
rect 7098 17320 7104 17332
rect 3191 17292 7104 17320
rect 3191 17289 3203 17292
rect 3145 17283 3203 17289
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 11054 17320 11060 17332
rect 9416 17292 11060 17320
rect 3786 17252 3792 17264
rect 3068 17224 3792 17252
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 2516 17116 2544 17147
rect 2958 17144 2964 17196
rect 3016 17184 3022 17196
rect 3068 17193 3096 17224
rect 3786 17212 3792 17224
rect 3844 17212 3850 17264
rect 4062 17212 4068 17264
rect 4120 17252 4126 17264
rect 4433 17255 4491 17261
rect 4433 17252 4445 17255
rect 4120 17224 4445 17252
rect 4120 17212 4126 17224
rect 4433 17221 4445 17224
rect 4479 17221 4491 17255
rect 5350 17252 5356 17264
rect 5263 17224 5356 17252
rect 4433 17215 4491 17221
rect 3053 17187 3111 17193
rect 3053 17184 3065 17187
rect 3016 17156 3065 17184
rect 3016 17144 3022 17156
rect 3053 17153 3065 17156
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 3418 17144 3424 17196
rect 3476 17184 3482 17196
rect 3697 17187 3755 17193
rect 3476 17156 3648 17184
rect 3476 17144 3482 17156
rect 3510 17116 3516 17128
rect 2516 17088 3516 17116
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 3620 17116 3648 17156
rect 3697 17153 3709 17187
rect 3743 17184 3755 17187
rect 4246 17184 4252 17196
rect 3743 17156 4252 17184
rect 3743 17153 3755 17156
rect 3697 17147 3755 17153
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 5276 17184 5304 17224
rect 5350 17212 5356 17224
rect 5408 17252 5414 17264
rect 6546 17252 6552 17264
rect 5408 17224 6552 17252
rect 5408 17212 5414 17224
rect 6546 17212 6552 17224
rect 6604 17212 6610 17264
rect 5442 17184 5448 17196
rect 4387 17156 5304 17184
rect 5403 17156 5448 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 5534 17144 5540 17196
rect 5592 17184 5598 17196
rect 7926 17184 7932 17196
rect 5592 17156 7932 17184
rect 5592 17144 5598 17156
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 9416 17193 9444 17292
rect 11054 17280 11060 17292
rect 11112 17320 11118 17332
rect 11974 17320 11980 17332
rect 11112 17292 11980 17320
rect 11112 17280 11118 17292
rect 11974 17280 11980 17292
rect 12032 17280 12038 17332
rect 14001 17323 14059 17329
rect 14001 17289 14013 17323
rect 14047 17320 14059 17323
rect 14182 17320 14188 17332
rect 14047 17292 14188 17320
rect 14047 17289 14059 17292
rect 14001 17283 14059 17289
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 17770 17320 17776 17332
rect 17731 17292 17776 17320
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 18414 17320 18420 17332
rect 18375 17292 18420 17320
rect 18414 17280 18420 17292
rect 18472 17280 18478 17332
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 19705 17323 19763 17329
rect 19705 17320 19717 17323
rect 19484 17292 19717 17320
rect 19484 17280 19490 17292
rect 19705 17289 19717 17292
rect 19751 17289 19763 17323
rect 19705 17283 19763 17289
rect 20717 17323 20775 17329
rect 20717 17289 20729 17323
rect 20763 17320 20775 17323
rect 23106 17320 23112 17332
rect 20763 17292 23112 17320
rect 20763 17289 20775 17292
rect 20717 17283 20775 17289
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 28902 17280 28908 17332
rect 28960 17320 28966 17332
rect 29181 17323 29239 17329
rect 29181 17320 29193 17323
rect 28960 17292 29193 17320
rect 28960 17280 28966 17292
rect 29181 17289 29193 17292
rect 29227 17289 29239 17323
rect 29181 17283 29239 17289
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 11882 17252 11888 17264
rect 9732 17224 10166 17252
rect 11843 17224 11888 17252
rect 9732 17212 9738 17224
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 18432 17224 20668 17252
rect 18432 17196 18460 17224
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17153 9459 17187
rect 9401 17147 9459 17153
rect 10962 17144 10968 17196
rect 11020 17184 11026 17196
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 11020 17156 12633 17184
rect 11020 17144 11026 17156
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 13909 17187 13967 17193
rect 13909 17153 13921 17187
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 8386 17116 8392 17128
rect 3620 17088 8392 17116
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17116 9735 17119
rect 9766 17116 9772 17128
rect 9723 17088 9772 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 9766 17076 9772 17088
rect 9824 17116 9830 17128
rect 10870 17116 10876 17128
rect 9824 17088 10876 17116
rect 9824 17076 9830 17088
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 13170 17116 13176 17128
rect 11112 17088 13176 17116
rect 11112 17076 11118 17088
rect 13170 17076 13176 17088
rect 13228 17116 13234 17128
rect 13924 17116 13952 17147
rect 15930 17144 15936 17196
rect 15988 17184 15994 17196
rect 16025 17187 16083 17193
rect 16025 17184 16037 17187
rect 15988 17156 16037 17184
rect 15988 17144 15994 17156
rect 16025 17153 16037 17156
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 16540 17156 17693 17184
rect 16540 17144 16546 17156
rect 17681 17153 17693 17156
rect 17727 17184 17739 17187
rect 18046 17184 18052 17196
rect 17727 17156 18052 17184
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 18138 17144 18144 17196
rect 18196 17184 18202 17196
rect 18325 17187 18383 17193
rect 18325 17184 18337 17187
rect 18196 17156 18337 17184
rect 18196 17144 18202 17156
rect 18325 17153 18337 17156
rect 18371 17153 18383 17187
rect 18325 17147 18383 17153
rect 18414 17144 18420 17196
rect 18472 17144 18478 17196
rect 20640 17193 20668 17224
rect 37550 17212 37556 17264
rect 37608 17252 37614 17264
rect 37608 17224 37872 17252
rect 37608 17212 37614 17224
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17153 19027 17187
rect 18969 17147 19027 17153
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 29089 17187 29147 17193
rect 29089 17153 29101 17187
rect 29135 17184 29147 17187
rect 37734 17184 37740 17196
rect 29135 17156 37740 17184
rect 29135 17153 29147 17156
rect 29089 17147 29147 17153
rect 13228 17088 13952 17116
rect 13228 17076 13234 17088
rect 15286 17076 15292 17128
rect 15344 17116 15350 17128
rect 18984 17116 19012 17147
rect 37734 17144 37740 17156
rect 37792 17144 37798 17196
rect 37844 17193 37872 17224
rect 37829 17187 37887 17193
rect 37829 17153 37841 17187
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 15344 17088 19012 17116
rect 15344 17076 15350 17088
rect 1857 17051 1915 17057
rect 1857 17017 1869 17051
rect 1903 17048 1915 17051
rect 2590 17048 2596 17060
rect 1903 17020 2596 17048
rect 1903 17017 1915 17020
rect 1857 17011 1915 17017
rect 2590 17008 2596 17020
rect 2648 17008 2654 17060
rect 8478 17048 8484 17060
rect 2700 17020 8484 17048
rect 1486 16940 1492 16992
rect 1544 16980 1550 16992
rect 2700 16980 2728 17020
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 11072 17020 12434 17048
rect 3786 16980 3792 16992
rect 1544 16952 2728 16980
rect 3747 16952 3792 16980
rect 1544 16940 1550 16952
rect 3786 16940 3792 16952
rect 3844 16940 3850 16992
rect 5537 16983 5595 16989
rect 5537 16949 5549 16983
rect 5583 16980 5595 16983
rect 6638 16980 6644 16992
rect 5583 16952 6644 16980
rect 5583 16949 5595 16952
rect 5537 16943 5595 16949
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 11072 16980 11100 17020
rect 10192 16952 11100 16980
rect 10192 16940 10198 16952
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 12406 16980 12434 17020
rect 15010 17008 15016 17060
rect 15068 17048 15074 17060
rect 22370 17048 22376 17060
rect 15068 17020 22376 17048
rect 15068 17008 15074 17020
rect 22370 17008 22376 17020
rect 22428 17008 22434 17060
rect 15194 16980 15200 16992
rect 11204 16952 11249 16980
rect 12406 16952 15200 16980
rect 11204 16940 11210 16952
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 16117 16983 16175 16989
rect 16117 16949 16129 16983
rect 16163 16980 16175 16983
rect 17034 16980 17040 16992
rect 16163 16952 17040 16980
rect 16163 16949 16175 16952
rect 16117 16943 16175 16949
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 19061 16983 19119 16989
rect 19061 16949 19073 16983
rect 19107 16980 19119 16983
rect 19150 16980 19156 16992
rect 19107 16952 19156 16980
rect 19107 16949 19119 16952
rect 19061 16943 19119 16949
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 37645 16983 37703 16989
rect 37645 16949 37657 16983
rect 37691 16980 37703 16983
rect 37826 16980 37832 16992
rect 37691 16952 37832 16980
rect 37691 16949 37703 16952
rect 37645 16943 37703 16949
rect 37826 16940 37832 16952
rect 37884 16940 37890 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 3510 16736 3516 16788
rect 3568 16776 3574 16788
rect 6178 16776 6184 16788
rect 3568 16748 6184 16776
rect 3568 16736 3574 16748
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 6546 16736 6552 16788
rect 6604 16776 6610 16788
rect 9582 16776 9588 16788
rect 6604 16748 9588 16776
rect 6604 16736 6610 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 17586 16776 17592 16788
rect 9784 16748 17592 16776
rect 6086 16708 6092 16720
rect 4080 16680 6092 16708
rect 2958 16640 2964 16652
rect 2608 16612 2964 16640
rect 1670 16532 1676 16584
rect 1728 16572 1734 16584
rect 2608 16581 2636 16612
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 1949 16575 2007 16581
rect 1949 16572 1961 16575
rect 1728 16544 1961 16572
rect 1728 16532 1734 16544
rect 1949 16541 1961 16544
rect 1995 16572 2007 16575
rect 2593 16575 2651 16581
rect 1995 16544 2544 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 1762 16464 1768 16516
rect 1820 16504 1826 16516
rect 2041 16507 2099 16513
rect 2041 16504 2053 16507
rect 1820 16476 2053 16504
rect 1820 16464 1826 16476
rect 2041 16473 2053 16476
rect 2087 16473 2099 16507
rect 2516 16504 2544 16544
rect 2593 16541 2605 16575
rect 2639 16574 2651 16575
rect 3237 16575 3295 16581
rect 2639 16546 2673 16574
rect 2639 16541 2651 16546
rect 2593 16535 2651 16541
rect 3237 16541 3249 16575
rect 3283 16572 3295 16575
rect 3970 16572 3976 16584
rect 3283 16544 3976 16572
rect 3283 16541 3295 16544
rect 3237 16535 3295 16541
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4080 16581 4108 16680
rect 6086 16668 6092 16680
rect 6144 16668 6150 16720
rect 6270 16668 6276 16720
rect 6328 16708 6334 16720
rect 6328 16680 7328 16708
rect 6328 16668 6334 16680
rect 5626 16640 5632 16652
rect 4356 16612 5632 16640
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 3418 16504 3424 16516
rect 2516 16476 3424 16504
rect 2041 16467 2099 16473
rect 3418 16464 3424 16476
rect 3476 16464 3482 16516
rect 3694 16464 3700 16516
rect 3752 16504 3758 16516
rect 4157 16507 4215 16513
rect 4157 16504 4169 16507
rect 3752 16476 4169 16504
rect 3752 16464 3758 16476
rect 4157 16473 4169 16476
rect 4203 16473 4215 16507
rect 4157 16467 4215 16473
rect 1946 16396 1952 16448
rect 2004 16436 2010 16448
rect 2685 16439 2743 16445
rect 2685 16436 2697 16439
rect 2004 16408 2697 16436
rect 2004 16396 2010 16408
rect 2685 16405 2697 16408
rect 2731 16405 2743 16439
rect 2685 16399 2743 16405
rect 3329 16439 3387 16445
rect 3329 16405 3341 16439
rect 3375 16436 3387 16439
rect 4356 16436 4384 16612
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 5166 16532 5172 16584
rect 5224 16572 5230 16584
rect 5224 16544 5269 16572
rect 5224 16532 5230 16544
rect 5534 16532 5540 16584
rect 5592 16572 5598 16584
rect 5813 16575 5871 16581
rect 5813 16572 5825 16575
rect 5592 16544 5825 16572
rect 5592 16532 5598 16544
rect 5813 16541 5825 16544
rect 5859 16541 5871 16575
rect 5813 16535 5871 16541
rect 5902 16532 5908 16584
rect 5960 16532 5966 16584
rect 6086 16532 6092 16584
rect 6144 16572 6150 16584
rect 7300 16581 7328 16680
rect 8110 16640 8116 16652
rect 8036 16612 8116 16640
rect 8036 16581 8064 16612
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 9784 16640 9812 16748
rect 17586 16736 17592 16748
rect 17644 16736 17650 16788
rect 25130 16776 25136 16788
rect 19352 16748 25136 16776
rect 12526 16708 12532 16720
rect 11716 16680 12532 16708
rect 8444 16612 9904 16640
rect 8444 16600 8450 16612
rect 9876 16581 9904 16612
rect 9968 16612 11560 16640
rect 6457 16575 6515 16581
rect 6457 16572 6469 16575
rect 6144 16544 6469 16572
rect 6144 16532 6150 16544
rect 6457 16541 6469 16544
rect 6503 16541 6515 16575
rect 6457 16535 6515 16541
rect 6549 16575 6607 16581
rect 6549 16541 6561 16575
rect 6595 16541 6607 16575
rect 6549 16535 6607 16541
rect 7285 16575 7343 16581
rect 7285 16541 7297 16575
rect 7331 16541 7343 16575
rect 7285 16535 7343 16541
rect 8021 16575 8079 16581
rect 8021 16541 8033 16575
rect 8067 16541 8079 16575
rect 8021 16535 8079 16541
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 5920 16504 5948 16532
rect 6564 16504 6592 16535
rect 5920 16476 6592 16504
rect 8754 16464 8760 16516
rect 8812 16504 8818 16516
rect 9968 16504 9996 16612
rect 10686 16572 10692 16584
rect 10647 16544 10692 16572
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 8812 16476 9996 16504
rect 11532 16504 11560 16612
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 11716 16572 11744 16680
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 12618 16668 12624 16720
rect 12676 16708 12682 16720
rect 12676 16680 14780 16708
rect 12676 16668 12682 16680
rect 12342 16640 12348 16652
rect 11655 16544 11744 16572
rect 11808 16612 12348 16640
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 11808 16504 11836 16612
rect 12342 16600 12348 16612
rect 12400 16640 12406 16652
rect 12400 16600 12434 16640
rect 11532 16476 11836 16504
rect 12406 16504 12434 16600
rect 12544 16612 13584 16640
rect 12544 16504 12572 16612
rect 13556 16581 13584 16612
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 14752 16581 14780 16680
rect 14826 16668 14832 16720
rect 14884 16708 14890 16720
rect 19352 16708 19380 16748
rect 25130 16736 25136 16748
rect 25188 16736 25194 16788
rect 14884 16680 17080 16708
rect 14884 16668 14890 16680
rect 16942 16640 16948 16652
rect 16684 16612 16948 16640
rect 14737 16575 14795 16581
rect 13688 16544 13733 16572
rect 13688 16532 13694 16544
rect 14737 16541 14749 16575
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 14829 16575 14887 16581
rect 14829 16541 14841 16575
rect 14875 16572 14887 16575
rect 15102 16572 15108 16584
rect 14875 16544 15108 16572
rect 14875 16541 14887 16544
rect 14829 16535 14887 16541
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 16684 16581 16712 16612
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17052 16640 17080 16680
rect 19306 16680 19380 16708
rect 22756 16680 23888 16708
rect 19306 16640 19334 16680
rect 17052 16612 19334 16640
rect 19444 16612 21312 16640
rect 15565 16575 15623 16581
rect 15565 16572 15577 16575
rect 15344 16544 15577 16572
rect 15344 16532 15350 16544
rect 15565 16541 15577 16544
rect 15611 16541 15623 16575
rect 15565 16535 15623 16541
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 16669 16535 16727 16541
rect 18690 16532 18696 16584
rect 18748 16572 18754 16584
rect 19444 16572 19472 16612
rect 21284 16581 21312 16612
rect 18748 16544 19472 16572
rect 21269 16575 21327 16581
rect 18748 16532 18754 16544
rect 21269 16541 21281 16575
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 22094 16532 22100 16584
rect 22152 16572 22158 16584
rect 22756 16572 22784 16680
rect 23293 16643 23351 16649
rect 23293 16640 23305 16643
rect 22152 16544 22784 16572
rect 22848 16612 23305 16640
rect 22152 16532 22158 16544
rect 12406 16476 12572 16504
rect 8812 16464 8818 16476
rect 16850 16464 16856 16516
rect 16908 16504 16914 16516
rect 17405 16507 17463 16513
rect 17405 16504 17417 16507
rect 16908 16476 17417 16504
rect 16908 16464 16914 16476
rect 17405 16473 17417 16476
rect 17451 16473 17463 16507
rect 17405 16467 17463 16473
rect 17494 16464 17500 16516
rect 17552 16504 17558 16516
rect 18049 16507 18107 16513
rect 17552 16476 17597 16504
rect 17552 16464 17558 16476
rect 18049 16473 18061 16507
rect 18095 16504 18107 16507
rect 19334 16504 19340 16516
rect 18095 16476 19340 16504
rect 18095 16473 18107 16476
rect 18049 16467 18107 16473
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 20070 16464 20076 16516
rect 20128 16504 20134 16516
rect 22848 16504 22876 16612
rect 23293 16609 23305 16612
rect 23339 16609 23351 16643
rect 23293 16603 23351 16609
rect 23860 16572 23888 16680
rect 26510 16572 26516 16584
rect 23860 16544 26516 16572
rect 26510 16532 26516 16544
rect 26568 16532 26574 16584
rect 37553 16575 37611 16581
rect 37553 16541 37565 16575
rect 37599 16572 37611 16575
rect 37918 16572 37924 16584
rect 37599 16544 37924 16572
rect 37599 16541 37611 16544
rect 37553 16535 37611 16541
rect 37918 16532 37924 16544
rect 37976 16532 37982 16584
rect 20128 16476 22876 16504
rect 23017 16507 23075 16513
rect 20128 16464 20134 16476
rect 23017 16473 23029 16507
rect 23063 16473 23075 16507
rect 23017 16467 23075 16473
rect 23109 16507 23167 16513
rect 23109 16473 23121 16507
rect 23155 16504 23167 16507
rect 23198 16504 23204 16516
rect 23155 16476 23204 16504
rect 23155 16473 23167 16476
rect 23109 16467 23167 16473
rect 3375 16408 4384 16436
rect 5261 16439 5319 16445
rect 3375 16405 3387 16408
rect 3329 16399 3387 16405
rect 5261 16405 5273 16439
rect 5307 16436 5319 16439
rect 5718 16436 5724 16448
rect 5307 16408 5724 16436
rect 5307 16405 5319 16408
rect 5261 16399 5319 16405
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 5902 16436 5908 16448
rect 5863 16408 5908 16436
rect 5902 16396 5908 16408
rect 5960 16396 5966 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7377 16439 7435 16445
rect 7377 16436 7389 16439
rect 6972 16408 7389 16436
rect 6972 16396 6978 16408
rect 7377 16405 7389 16408
rect 7423 16405 7435 16439
rect 7377 16399 7435 16405
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 8113 16439 8171 16445
rect 8113 16436 8125 16439
rect 7708 16408 8125 16436
rect 7708 16396 7714 16408
rect 8113 16405 8125 16408
rect 8159 16405 8171 16439
rect 8113 16399 8171 16405
rect 9953 16439 10011 16445
rect 9953 16405 9965 16439
rect 9999 16436 10011 16439
rect 10134 16436 10140 16448
rect 9999 16408 10140 16436
rect 9999 16405 10011 16408
rect 9953 16399 10011 16405
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 10781 16439 10839 16445
rect 10781 16405 10793 16439
rect 10827 16436 10839 16439
rect 11514 16436 11520 16448
rect 10827 16408 11520 16436
rect 10827 16405 10839 16408
rect 10781 16399 10839 16405
rect 11514 16396 11520 16408
rect 11572 16396 11578 16448
rect 11698 16436 11704 16448
rect 11659 16408 11704 16436
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 15381 16439 15439 16445
rect 15381 16405 15393 16439
rect 15427 16436 15439 16439
rect 16298 16436 16304 16448
rect 15427 16408 16304 16436
rect 15427 16405 15439 16408
rect 15381 16399 15439 16405
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16758 16436 16764 16448
rect 16719 16408 16764 16436
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 21361 16439 21419 16445
rect 21361 16405 21373 16439
rect 21407 16436 21419 16439
rect 22646 16436 22652 16448
rect 21407 16408 22652 16436
rect 21407 16405 21419 16408
rect 21361 16399 21419 16405
rect 22646 16396 22652 16408
rect 22704 16396 22710 16448
rect 22738 16396 22744 16448
rect 22796 16436 22802 16448
rect 23032 16436 23060 16467
rect 23198 16464 23204 16476
rect 23256 16464 23262 16516
rect 38102 16504 38108 16516
rect 38063 16476 38108 16504
rect 38102 16464 38108 16476
rect 38160 16464 38166 16516
rect 22796 16408 23060 16436
rect 37369 16439 37427 16445
rect 22796 16396 22802 16408
rect 37369 16405 37381 16439
rect 37415 16436 37427 16439
rect 37918 16436 37924 16448
rect 37415 16408 37924 16436
rect 37415 16405 37427 16408
rect 37369 16399 37427 16405
rect 37918 16396 37924 16408
rect 37976 16396 37982 16448
rect 38194 16436 38200 16448
rect 38155 16408 38200 16436
rect 38194 16396 38200 16408
rect 38252 16396 38258 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 3326 16232 3332 16244
rect 3287 16204 3332 16232
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 3418 16192 3424 16244
rect 3476 16232 3482 16244
rect 6917 16235 6975 16241
rect 3476 16204 6040 16232
rect 3476 16192 3482 16204
rect 4154 16164 4160 16176
rect 4115 16136 4160 16164
rect 4154 16124 4160 16136
rect 4212 16124 4218 16176
rect 4249 16167 4307 16173
rect 4249 16133 4261 16167
rect 4295 16164 4307 16167
rect 5902 16164 5908 16176
rect 4295 16136 5908 16164
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 5902 16124 5908 16136
rect 5960 16124 5966 16176
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16065 1639 16099
rect 2590 16096 2596 16108
rect 2551 16068 2596 16096
rect 1581 16059 1639 16065
rect 1596 15960 1624 16059
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 2958 16056 2964 16108
rect 3016 16096 3022 16108
rect 3237 16099 3295 16105
rect 3237 16096 3249 16099
rect 3016 16068 3249 16096
rect 3016 16056 3022 16068
rect 3237 16065 3249 16068
rect 3283 16065 3295 16099
rect 3237 16059 3295 16065
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6012 16096 6040 16204
rect 6917 16201 6929 16235
rect 6963 16232 6975 16235
rect 7190 16232 7196 16244
rect 6963 16204 7196 16232
rect 6963 16201 6975 16204
rect 6917 16195 6975 16201
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 8202 16232 8208 16244
rect 8163 16204 8208 16232
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 8849 16235 8907 16241
rect 8849 16201 8861 16235
rect 8895 16232 8907 16235
rect 9674 16232 9680 16244
rect 8895 16204 9680 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10410 16232 10416 16244
rect 10371 16204 10416 16232
rect 10410 16192 10416 16204
rect 10468 16192 10474 16244
rect 11057 16235 11115 16241
rect 11057 16201 11069 16235
rect 11103 16232 11115 16235
rect 11238 16232 11244 16244
rect 11103 16204 11244 16232
rect 11103 16201 11115 16204
rect 11057 16195 11115 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 13722 16232 13728 16244
rect 13683 16204 13728 16232
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 17494 16232 17500 16244
rect 16163 16204 17500 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 19334 16192 19340 16244
rect 19392 16232 19398 16244
rect 22094 16232 22100 16244
rect 19392 16204 22100 16232
rect 19392 16192 19398 16204
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 22554 16192 22560 16244
rect 22612 16232 22618 16244
rect 24578 16232 24584 16244
rect 22612 16204 24584 16232
rect 22612 16192 22618 16204
rect 24578 16192 24584 16204
rect 24636 16192 24642 16244
rect 37734 16192 37740 16244
rect 37792 16232 37798 16244
rect 38105 16235 38163 16241
rect 38105 16232 38117 16235
rect 37792 16204 38117 16232
rect 37792 16192 37798 16204
rect 38105 16201 38117 16204
rect 38151 16201 38163 16235
rect 38105 16195 38163 16201
rect 11882 16164 11888 16176
rect 8128 16136 10364 16164
rect 11843 16136 11888 16164
rect 6086 16096 6092 16108
rect 5859 16068 6092 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 8128 16105 8156 16136
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16096 6883 16099
rect 8113 16099 8171 16105
rect 8113 16096 8125 16099
rect 6871 16068 8125 16096
rect 6871 16065 6883 16068
rect 6825 16059 6883 16065
rect 8113 16065 8125 16068
rect 8159 16065 8171 16099
rect 8754 16096 8760 16108
rect 8715 16068 8760 16096
rect 8113 16059 8171 16065
rect 8754 16056 8760 16068
rect 8812 16056 8818 16108
rect 9674 16096 9680 16108
rect 9635 16068 9680 16096
rect 9674 16056 9680 16068
rect 9732 16056 9738 16108
rect 10336 16105 10364 16136
rect 11882 16124 11888 16136
rect 11940 16124 11946 16176
rect 12618 16164 12624 16176
rect 12579 16136 12624 16164
rect 12618 16124 12624 16136
rect 12676 16124 12682 16176
rect 17034 16164 17040 16176
rect 16995 16136 17040 16164
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 19150 16164 19156 16176
rect 19111 16136 19156 16164
rect 19150 16124 19156 16136
rect 19208 16124 19214 16176
rect 20533 16167 20591 16173
rect 20533 16133 20545 16167
rect 20579 16164 20591 16167
rect 20622 16164 20628 16176
rect 20579 16136 20628 16164
rect 20579 16133 20591 16136
rect 20533 16127 20591 16133
rect 20622 16124 20628 16136
rect 20680 16124 20686 16176
rect 22462 16124 22468 16176
rect 22520 16164 22526 16176
rect 22833 16167 22891 16173
rect 22833 16164 22845 16167
rect 22520 16136 22845 16164
rect 22520 16124 22526 16136
rect 22833 16133 22845 16136
rect 22879 16133 22891 16167
rect 22833 16127 22891 16133
rect 22922 16124 22928 16176
rect 22980 16164 22986 16176
rect 23290 16164 23296 16176
rect 22980 16136 23296 16164
rect 22980 16124 22986 16136
rect 23290 16124 23296 16136
rect 23348 16124 23354 16176
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16096 10379 16099
rect 10965 16099 11023 16105
rect 10965 16096 10977 16099
rect 10367 16068 10977 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 10965 16065 10977 16068
rect 11011 16096 11023 16099
rect 11054 16096 11060 16108
rect 11011 16068 11060 16096
rect 11011 16065 11023 16068
rect 10965 16059 11023 16065
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 11606 16056 11612 16108
rect 11664 16056 11670 16108
rect 13170 16056 13176 16108
rect 13228 16096 13234 16108
rect 13633 16099 13691 16105
rect 13633 16096 13645 16099
rect 13228 16068 13645 16096
rect 13228 16056 13234 16068
rect 13633 16065 13645 16068
rect 13679 16065 13691 16099
rect 16298 16096 16304 16108
rect 16259 16068 16304 16096
rect 13633 16059 13691 16065
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 27433 16099 27491 16105
rect 27433 16065 27445 16099
rect 27479 16096 27491 16099
rect 33505 16099 33563 16105
rect 27479 16068 31754 16096
rect 27479 16065 27491 16068
rect 27433 16059 27491 16065
rect 2685 16031 2743 16037
rect 2685 15997 2697 16031
rect 2731 16028 2743 16031
rect 4706 16028 4712 16040
rect 2731 16000 4712 16028
rect 2731 15997 2743 16000
rect 2685 15991 2743 15997
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 16028 5227 16031
rect 5442 16028 5448 16040
rect 5215 16000 5448 16028
rect 5215 15997 5227 16000
rect 5169 15991 5227 15997
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 8294 16028 8300 16040
rect 5951 16000 8300 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 11624 16028 11652 16056
rect 8444 16000 11652 16028
rect 16945 16031 17003 16037
rect 8444 15988 8450 16000
rect 16945 15997 16957 16031
rect 16991 15997 17003 16031
rect 16945 15991 17003 15997
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 15997 18015 16031
rect 17957 15991 18015 15997
rect 7190 15960 7196 15972
rect 1596 15932 7196 15960
rect 7190 15920 7196 15932
rect 7248 15920 7254 15972
rect 10686 15960 10692 15972
rect 9692 15932 10692 15960
rect 9692 15904 9720 15932
rect 10686 15920 10692 15932
rect 10744 15920 10750 15972
rect 11606 15920 11612 15972
rect 11664 15960 11670 15972
rect 16960 15960 16988 15991
rect 11664 15932 16988 15960
rect 17972 15960 18000 15991
rect 18322 15988 18328 16040
rect 18380 16028 18386 16040
rect 18874 16028 18880 16040
rect 18380 16000 18880 16028
rect 18380 15988 18386 16000
rect 18874 15988 18880 16000
rect 18932 16028 18938 16040
rect 19061 16031 19119 16037
rect 19061 16028 19073 16031
rect 18932 16000 19073 16028
rect 18932 15988 18938 16000
rect 19061 15997 19073 16000
rect 19107 15997 19119 16031
rect 19334 16028 19340 16040
rect 19295 16000 19340 16028
rect 19061 15991 19119 15997
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 20441 16031 20499 16037
rect 20441 15997 20453 16031
rect 20487 15997 20499 16031
rect 20441 15991 20499 15997
rect 20070 15960 20076 15972
rect 17972 15932 20076 15960
rect 11664 15920 11670 15932
rect 20070 15920 20076 15932
rect 20128 15920 20134 15972
rect 20456 15960 20484 15991
rect 20622 15988 20628 16040
rect 20680 16028 20686 16040
rect 20717 16031 20775 16037
rect 20717 16028 20729 16031
rect 20680 16000 20729 16028
rect 20680 15988 20686 16000
rect 20717 15997 20729 16000
rect 20763 15997 20775 16031
rect 20717 15991 20775 15997
rect 22741 16031 22799 16037
rect 22741 15997 22753 16031
rect 22787 16028 22799 16031
rect 23566 16028 23572 16040
rect 22787 16000 23152 16028
rect 23527 16000 23572 16028
rect 22787 15997 22799 16000
rect 22741 15991 22799 15997
rect 21910 15960 21916 15972
rect 20456 15932 21916 15960
rect 21910 15920 21916 15932
rect 21968 15920 21974 15972
rect 23124 15960 23152 16000
rect 23566 15988 23572 16000
rect 23624 15988 23630 16040
rect 26142 15988 26148 16040
rect 26200 16028 26206 16040
rect 26237 16031 26295 16037
rect 26237 16028 26249 16031
rect 26200 16000 26249 16028
rect 26200 15988 26206 16000
rect 26237 15997 26249 16000
rect 26283 15997 26295 16031
rect 31726 16028 31754 16068
rect 33505 16065 33517 16099
rect 33551 16096 33563 16099
rect 37642 16096 37648 16108
rect 33551 16068 37648 16096
rect 33551 16065 33563 16068
rect 33505 16059 33563 16065
rect 37642 16056 37648 16068
rect 37700 16056 37706 16108
rect 38286 16096 38292 16108
rect 38247 16068 38292 16096
rect 38286 16056 38292 16068
rect 38344 16056 38350 16108
rect 36538 16028 36544 16040
rect 31726 16000 36544 16028
rect 26237 15991 26295 15997
rect 36538 15988 36544 16000
rect 36596 15988 36602 16040
rect 23474 15960 23480 15972
rect 23124 15932 23480 15960
rect 23474 15920 23480 15932
rect 23532 15920 23538 15972
rect 26418 15960 26424 15972
rect 23584 15932 26424 15960
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 2590 15852 2596 15904
rect 2648 15892 2654 15904
rect 5350 15892 5356 15904
rect 2648 15864 5356 15892
rect 2648 15852 2654 15864
rect 5350 15852 5356 15864
rect 5408 15892 5414 15904
rect 5534 15892 5540 15904
rect 5408 15864 5540 15892
rect 5408 15852 5414 15864
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6086 15852 6092 15904
rect 6144 15892 6150 15904
rect 9674 15892 9680 15904
rect 6144 15864 9680 15892
rect 6144 15852 6150 15864
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 9769 15895 9827 15901
rect 9769 15861 9781 15895
rect 9815 15892 9827 15895
rect 10226 15892 10232 15904
rect 9815 15864 10232 15892
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 10226 15852 10232 15864
rect 10284 15852 10290 15904
rect 12066 15852 12072 15904
rect 12124 15892 12130 15904
rect 18782 15892 18788 15904
rect 12124 15864 18788 15892
rect 12124 15852 12130 15864
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 20622 15892 20628 15904
rect 19392 15864 20628 15892
rect 19392 15852 19398 15864
rect 20622 15852 20628 15864
rect 20680 15852 20686 15904
rect 22097 15895 22155 15901
rect 22097 15861 22109 15895
rect 22143 15892 22155 15895
rect 22922 15892 22928 15904
rect 22143 15864 22928 15892
rect 22143 15861 22155 15864
rect 22097 15855 22155 15861
rect 22922 15852 22928 15864
rect 22980 15852 22986 15904
rect 23106 15852 23112 15904
rect 23164 15892 23170 15904
rect 23584 15892 23612 15932
rect 26418 15920 26424 15932
rect 26476 15920 26482 15972
rect 23164 15864 23612 15892
rect 23164 15852 23170 15864
rect 24854 15852 24860 15904
rect 24912 15892 24918 15904
rect 27525 15895 27583 15901
rect 27525 15892 27537 15895
rect 24912 15864 27537 15892
rect 24912 15852 24918 15864
rect 27525 15861 27537 15864
rect 27571 15861 27583 15895
rect 33318 15892 33324 15904
rect 33279 15864 33324 15892
rect 27525 15855 27583 15861
rect 33318 15852 33324 15864
rect 33376 15852 33382 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 6641 15691 6699 15697
rect 6641 15657 6653 15691
rect 6687 15688 6699 15691
rect 8386 15688 8392 15700
rect 6687 15660 8392 15688
rect 6687 15657 6699 15660
rect 6641 15651 6699 15657
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 9401 15691 9459 15697
rect 9401 15657 9413 15691
rect 9447 15688 9459 15691
rect 10502 15688 10508 15700
rect 9447 15660 10508 15688
rect 9447 15657 9459 15660
rect 9401 15651 9459 15657
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 16574 15688 16580 15700
rect 10612 15660 16580 15688
rect 3142 15620 3148 15632
rect 3103 15592 3148 15620
rect 3142 15580 3148 15592
rect 3200 15580 3206 15632
rect 5905 15623 5963 15629
rect 5905 15589 5917 15623
rect 5951 15620 5963 15623
rect 10612 15620 10640 15660
rect 16574 15648 16580 15660
rect 16632 15648 16638 15700
rect 18782 15648 18788 15700
rect 18840 15688 18846 15700
rect 22002 15688 22008 15700
rect 18840 15660 22008 15688
rect 18840 15648 18846 15660
rect 22002 15648 22008 15660
rect 22060 15688 22066 15700
rect 22554 15688 22560 15700
rect 22060 15660 22560 15688
rect 22060 15648 22066 15660
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 22646 15648 22652 15700
rect 22704 15688 22710 15700
rect 22704 15660 26372 15688
rect 22704 15648 22710 15660
rect 5951 15592 10640 15620
rect 5951 15589 5963 15592
rect 5905 15583 5963 15589
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 12250 15620 12256 15632
rect 10744 15592 12256 15620
rect 10744 15580 10750 15592
rect 12250 15580 12256 15592
rect 12308 15620 12314 15632
rect 13170 15620 13176 15632
rect 12308 15592 13176 15620
rect 12308 15580 12314 15592
rect 13170 15580 13176 15592
rect 13228 15580 13234 15632
rect 20622 15580 20628 15632
rect 20680 15620 20686 15632
rect 20680 15592 23520 15620
rect 20680 15580 20686 15592
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 2823 15524 10333 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 10321 15521 10333 15524
rect 10367 15552 10379 15555
rect 23106 15552 23112 15564
rect 10367 15524 23112 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 23492 15561 23520 15592
rect 23477 15555 23535 15561
rect 23477 15521 23489 15555
rect 23523 15521 23535 15555
rect 26142 15552 26148 15564
rect 26103 15524 26148 15552
rect 23477 15515 23535 15521
rect 26142 15512 26148 15524
rect 26200 15512 26206 15564
rect 26344 15561 26372 15660
rect 30009 15623 30067 15629
rect 30009 15589 30021 15623
rect 30055 15620 30067 15623
rect 34790 15620 34796 15632
rect 30055 15592 34796 15620
rect 30055 15589 30067 15592
rect 30009 15583 30067 15589
rect 34790 15580 34796 15592
rect 34848 15580 34854 15632
rect 26329 15555 26387 15561
rect 26329 15521 26341 15555
rect 26375 15521 26387 15555
rect 27890 15552 27896 15564
rect 27851 15524 27896 15552
rect 26329 15515 26387 15521
rect 27890 15512 27896 15524
rect 27948 15512 27954 15564
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15453 1639 15487
rect 2958 15484 2964 15496
rect 2919 15456 2964 15484
rect 1581 15447 1639 15453
rect 1596 15416 1624 15447
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 5810 15484 5816 15496
rect 5771 15456 5816 15484
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 6546 15484 6552 15496
rect 6507 15456 6552 15484
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 9674 15484 9680 15496
rect 9355 15456 9680 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 12897 15487 12955 15493
rect 12897 15484 12909 15487
rect 12268 15456 12909 15484
rect 1596 15388 2774 15416
rect 1762 15348 1768 15360
rect 1723 15320 1768 15348
rect 1762 15308 1768 15320
rect 1820 15308 1826 15360
rect 2746 15348 2774 15388
rect 4154 15376 4160 15428
rect 4212 15416 4218 15428
rect 4341 15419 4399 15425
rect 4341 15416 4353 15419
rect 4212 15388 4353 15416
rect 4212 15376 4218 15388
rect 4341 15385 4353 15388
rect 4387 15385 4399 15419
rect 4341 15379 4399 15385
rect 4433 15419 4491 15425
rect 4433 15385 4445 15419
rect 4479 15416 4491 15419
rect 5258 15416 5264 15428
rect 4479 15388 5264 15416
rect 4479 15385 4491 15388
rect 4433 15379 4491 15385
rect 5258 15376 5264 15388
rect 5316 15376 5322 15428
rect 5350 15376 5356 15428
rect 5408 15416 5414 15428
rect 5408 15388 5453 15416
rect 6564 15388 6960 15416
rect 5408 15376 5414 15388
rect 6564 15348 6592 15388
rect 2746 15320 6592 15348
rect 6932 15348 6960 15388
rect 7006 15376 7012 15428
rect 7064 15416 7070 15428
rect 7561 15419 7619 15425
rect 7561 15416 7573 15419
rect 7064 15388 7573 15416
rect 7064 15376 7070 15388
rect 7561 15385 7573 15388
rect 7607 15385 7619 15419
rect 7561 15379 7619 15385
rect 7650 15376 7656 15428
rect 7708 15416 7714 15428
rect 8570 15416 8576 15428
rect 7708 15388 7753 15416
rect 8531 15388 8576 15416
rect 7708 15376 7714 15388
rect 8570 15376 8576 15388
rect 8628 15376 8634 15428
rect 10042 15416 10048 15428
rect 10003 15388 10048 15416
rect 10042 15376 10048 15388
rect 10100 15376 10106 15428
rect 10134 15376 10140 15428
rect 10192 15416 10198 15428
rect 11425 15419 11483 15425
rect 10192 15388 10237 15416
rect 10192 15376 10198 15388
rect 11425 15385 11437 15419
rect 11471 15385 11483 15419
rect 11425 15379 11483 15385
rect 8018 15348 8024 15360
rect 6932 15320 8024 15348
rect 8018 15308 8024 15320
rect 8076 15308 8082 15360
rect 9858 15308 9864 15360
rect 9916 15348 9922 15360
rect 10410 15348 10416 15360
rect 9916 15320 10416 15348
rect 9916 15308 9922 15320
rect 10410 15308 10416 15320
rect 10468 15308 10474 15360
rect 11440 15348 11468 15379
rect 11514 15376 11520 15428
rect 11572 15416 11578 15428
rect 11572 15388 11617 15416
rect 11572 15376 11578 15388
rect 11882 15376 11888 15428
rect 11940 15416 11946 15428
rect 12268 15416 12296 15456
rect 12897 15453 12909 15456
rect 12943 15453 12955 15487
rect 13170 15484 13176 15496
rect 13131 15456 13176 15484
rect 12897 15447 12955 15453
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18104 15456 18705 15484
rect 18104 15444 18110 15456
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15484 19487 15487
rect 20254 15484 20260 15496
rect 19475 15456 20260 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 11940 15388 12296 15416
rect 11940 15376 11946 15388
rect 12342 15376 12348 15428
rect 12400 15416 12406 15428
rect 12437 15419 12495 15425
rect 12437 15416 12449 15419
rect 12400 15388 12449 15416
rect 12400 15376 12406 15388
rect 12437 15385 12449 15388
rect 12483 15416 12495 15419
rect 15654 15416 15660 15428
rect 12483 15388 15660 15416
rect 12483 15385 12495 15388
rect 12437 15379 12495 15385
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 16850 15416 16856 15428
rect 16811 15388 16856 15416
rect 16850 15376 16856 15388
rect 16908 15376 16914 15428
rect 16945 15419 17003 15425
rect 16945 15385 16957 15419
rect 16991 15385 17003 15419
rect 17862 15416 17868 15428
rect 17823 15388 17868 15416
rect 16945 15379 17003 15385
rect 11606 15348 11612 15360
rect 11440 15320 11612 15348
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 16960 15348 16988 15379
rect 17862 15376 17868 15388
rect 17920 15376 17926 15428
rect 18708 15416 18736 15447
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20990 15444 20996 15496
rect 21048 15484 21054 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 21048 15456 21097 15484
rect 21048 15444 21054 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 21177 15487 21235 15493
rect 21177 15453 21189 15487
rect 21223 15484 21235 15487
rect 22462 15484 22468 15496
rect 21223 15456 22468 15484
rect 21223 15453 21235 15456
rect 21177 15447 21235 15453
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 21358 15416 21364 15428
rect 18708 15388 21364 15416
rect 21358 15376 21364 15388
rect 21416 15376 21422 15428
rect 22833 15419 22891 15425
rect 22833 15385 22845 15419
rect 22879 15385 22891 15419
rect 22833 15379 22891 15385
rect 11756 15320 16988 15348
rect 18785 15351 18843 15357
rect 11756 15308 11762 15320
rect 18785 15317 18797 15351
rect 18831 15348 18843 15351
rect 19426 15348 19432 15360
rect 18831 15320 19432 15348
rect 18831 15317 18843 15320
rect 18785 15311 18843 15317
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 19521 15351 19579 15357
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 22002 15348 22008 15360
rect 19567 15320 22008 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 22848 15348 22876 15379
rect 22922 15376 22928 15428
rect 22980 15416 22986 15428
rect 22980 15388 23025 15416
rect 22980 15376 22986 15388
rect 23106 15376 23112 15428
rect 23164 15416 23170 15428
rect 24673 15419 24731 15425
rect 24673 15416 24685 15419
rect 23164 15388 24685 15416
rect 23164 15376 23170 15388
rect 24673 15385 24685 15388
rect 24719 15385 24731 15419
rect 24673 15379 24731 15385
rect 24765 15419 24823 15425
rect 24765 15385 24777 15419
rect 24811 15416 24823 15419
rect 25038 15416 25044 15428
rect 24811 15388 25044 15416
rect 24811 15385 24823 15388
rect 24765 15379 24823 15385
rect 25038 15376 25044 15388
rect 25096 15376 25102 15428
rect 25685 15419 25743 15425
rect 25685 15385 25697 15419
rect 25731 15416 25743 15419
rect 26050 15416 26056 15428
rect 25731 15388 26056 15416
rect 25731 15385 25743 15388
rect 25685 15379 25743 15385
rect 26050 15376 26056 15388
rect 26108 15376 26114 15428
rect 29822 15416 29828 15428
rect 29783 15388 29828 15416
rect 29822 15376 29828 15388
rect 29880 15376 29886 15428
rect 23474 15348 23480 15360
rect 22848 15320 23480 15348
rect 23474 15308 23480 15320
rect 23532 15308 23538 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 5408 15116 11008 15144
rect 5408 15104 5414 15116
rect 2041 15079 2099 15085
rect 2041 15045 2053 15079
rect 2087 15076 2099 15079
rect 3786 15076 3792 15088
rect 2087 15048 3792 15076
rect 2087 15045 2099 15048
rect 2041 15039 2099 15045
rect 3786 15036 3792 15048
rect 3844 15036 3850 15088
rect 5718 15036 5724 15088
rect 5776 15076 5782 15088
rect 6733 15079 6791 15085
rect 6733 15076 6745 15079
rect 5776 15048 6745 15076
rect 5776 15036 5782 15048
rect 6733 15045 6745 15048
rect 6779 15045 6791 15079
rect 6733 15039 6791 15045
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 8294 15076 8300 15088
rect 6880 15048 8300 15076
rect 6880 15036 6886 15048
rect 8294 15036 8300 15048
rect 8352 15036 8358 15088
rect 10226 15076 10232 15088
rect 10187 15048 10232 15076
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 7282 14966 7288 15018
rect 7340 15006 7346 15018
rect 7340 14978 7383 15006
rect 7340 14966 7346 14978
rect 7650 14968 7656 15020
rect 7708 15008 7714 15020
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7708 14980 7757 15008
rect 7708 14968 7714 14980
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 9125 15011 9183 15017
rect 9125 14977 9137 15011
rect 9171 15008 9183 15011
rect 9766 15008 9772 15020
rect 9171 14980 9772 15008
rect 9171 14977 9183 14980
rect 9125 14971 9183 14977
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 3326 14940 3332 14952
rect 1903 14912 3332 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 3694 14940 3700 14952
rect 3655 14912 3700 14940
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14909 4215 14943
rect 4157 14903 4215 14909
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14940 4399 14943
rect 5902 14940 5908 14952
rect 4387 14912 5908 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 1946 14832 1952 14884
rect 2004 14872 2010 14884
rect 4172 14872 4200 14903
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 5997 14943 6055 14949
rect 5997 14909 6009 14943
rect 6043 14909 6055 14943
rect 5997 14903 6055 14909
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 7929 14943 7987 14949
rect 6687 14912 7144 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 2004 14844 4200 14872
rect 6012 14872 6040 14903
rect 6822 14872 6828 14884
rect 6012 14844 6828 14872
rect 2004 14832 2010 14844
rect 6822 14832 6828 14844
rect 6880 14832 6886 14884
rect 7116 14804 7144 14912
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 8202 14940 8208 14952
rect 7975 14912 8208 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8478 14900 8484 14952
rect 8536 14940 8542 14952
rect 10138 14943 10196 14949
rect 8536 14912 10088 14940
rect 8536 14900 8542 14912
rect 9858 14872 9864 14884
rect 7944 14844 9864 14872
rect 7944 14804 7972 14844
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 10060 14872 10088 14912
rect 10138 14909 10150 14943
rect 10184 14940 10196 14943
rect 10226 14940 10232 14952
rect 10184 14912 10232 14940
rect 10184 14909 10196 14912
rect 10138 14903 10196 14909
rect 10226 14900 10232 14912
rect 10284 14900 10290 14952
rect 10980 14940 11008 15116
rect 11698 15104 11704 15156
rect 11756 15104 11762 15156
rect 12437 15147 12495 15153
rect 12437 15113 12449 15147
rect 12483 15144 12495 15147
rect 12710 15144 12716 15156
rect 12483 15116 12716 15144
rect 12483 15113 12495 15116
rect 12437 15107 12495 15113
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 16574 15104 16580 15156
rect 16632 15144 16638 15156
rect 16632 15116 17908 15144
rect 16632 15104 16638 15116
rect 11149 15079 11207 15085
rect 11149 15045 11161 15079
rect 11195 15076 11207 15079
rect 11422 15076 11428 15088
rect 11195 15048 11428 15076
rect 11195 15045 11207 15048
rect 11149 15039 11207 15045
rect 11422 15036 11428 15048
rect 11480 15036 11486 15088
rect 11716 15076 11744 15104
rect 16206 15076 16212 15088
rect 11716 15048 16212 15076
rect 16206 15036 16212 15048
rect 16264 15036 16270 15088
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 17037 15079 17095 15085
rect 17037 15076 17049 15079
rect 16816 15048 17049 15076
rect 16816 15036 16822 15048
rect 17037 15045 17049 15048
rect 17083 15045 17095 15079
rect 17880 15076 17908 15116
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18012 15116 23152 15144
rect 18012 15104 18018 15116
rect 21818 15076 21824 15088
rect 17880 15048 21824 15076
rect 17037 15039 17095 15045
rect 21818 15036 21824 15048
rect 21876 15036 21882 15088
rect 22094 15036 22100 15088
rect 22152 15076 22158 15088
rect 23124 15085 23152 15116
rect 22189 15079 22247 15085
rect 22189 15076 22201 15079
rect 22152 15048 22201 15076
rect 22152 15036 22158 15048
rect 22189 15045 22201 15048
rect 22235 15045 22247 15079
rect 22189 15039 22247 15045
rect 23109 15079 23167 15085
rect 23109 15045 23121 15079
rect 23155 15076 23167 15079
rect 23566 15076 23572 15088
rect 23155 15048 23572 15076
rect 23155 15045 23167 15048
rect 23109 15039 23167 15045
rect 23566 15036 23572 15048
rect 23624 15036 23630 15088
rect 23845 15079 23903 15085
rect 23845 15045 23857 15079
rect 23891 15076 23903 15079
rect 24578 15076 24584 15088
rect 23891 15048 24584 15076
rect 23891 15045 23903 15048
rect 23845 15039 23903 15045
rect 24578 15036 24584 15048
rect 24636 15036 24642 15088
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 11882 15008 11888 15020
rect 11747 14980 11888 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 12250 14968 12256 15020
rect 12308 15008 12314 15020
rect 12345 15011 12403 15017
rect 12345 15008 12357 15011
rect 12308 14980 12357 15008
rect 12308 14968 12314 14980
rect 12345 14977 12357 14980
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 16666 15008 16672 15020
rect 14056 14980 16672 15008
rect 14056 14968 14062 14980
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 18414 15008 18420 15020
rect 18375 14980 18420 15008
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 18782 14968 18788 15020
rect 18840 15008 18846 15020
rect 19061 15011 19119 15017
rect 19061 15008 19073 15011
rect 18840 14980 19073 15008
rect 18840 14968 18846 14980
rect 19061 14977 19073 14980
rect 19107 14977 19119 15011
rect 19061 14971 19119 14977
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 15008 21327 15011
rect 21358 15008 21364 15020
rect 21315 14980 21364 15008
rect 21315 14977 21327 14980
rect 21269 14971 21327 14977
rect 21358 14968 21364 14980
rect 21416 14968 21422 15020
rect 11974 14940 11980 14952
rect 10980 14912 11980 14940
rect 11974 14900 11980 14912
rect 12032 14900 12038 14952
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 16945 14943 17003 14949
rect 16945 14940 16957 14943
rect 16632 14912 16957 14940
rect 16632 14900 16638 14912
rect 16945 14909 16957 14912
rect 16991 14909 17003 14943
rect 17218 14940 17224 14952
rect 17179 14912 17224 14940
rect 16945 14903 17003 14909
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 17586 14900 17592 14952
rect 17644 14940 17650 14952
rect 20898 14940 20904 14952
rect 17644 14912 20904 14940
rect 17644 14900 17650 14912
rect 20898 14900 20904 14912
rect 20956 14900 20962 14952
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 22097 14943 22155 14949
rect 22097 14940 22109 14943
rect 21968 14912 22109 14940
rect 21968 14900 21974 14912
rect 22097 14909 22109 14912
rect 22143 14909 22155 14943
rect 22097 14903 22155 14909
rect 11882 14872 11888 14884
rect 10060 14844 11888 14872
rect 11882 14832 11888 14844
rect 11940 14832 11946 14884
rect 15010 14832 15016 14884
rect 15068 14872 15074 14884
rect 20990 14872 20996 14884
rect 15068 14844 20996 14872
rect 15068 14832 15074 14844
rect 20990 14832 20996 14844
rect 21048 14832 21054 14884
rect 22112 14872 22140 14903
rect 22922 14900 22928 14952
rect 22980 14940 22986 14952
rect 23753 14943 23811 14949
rect 23753 14940 23765 14943
rect 22980 14912 23765 14940
rect 22980 14900 22986 14912
rect 23753 14909 23765 14912
rect 23799 14909 23811 14943
rect 24854 14940 24860 14952
rect 23753 14903 23811 14909
rect 23860 14912 24860 14940
rect 23860 14872 23888 14912
rect 24854 14900 24860 14912
rect 24912 14900 24918 14952
rect 27706 14900 27712 14952
rect 27764 14940 27770 14952
rect 27982 14940 27988 14952
rect 27764 14912 27988 14940
rect 27764 14900 27770 14912
rect 27982 14900 27988 14912
rect 28040 14900 28046 14952
rect 24302 14872 24308 14884
rect 22112 14844 23888 14872
rect 24263 14844 24308 14872
rect 24302 14832 24308 14844
rect 24360 14832 24366 14884
rect 26878 14832 26884 14884
rect 26936 14872 26942 14884
rect 33594 14872 33600 14884
rect 26936 14844 33600 14872
rect 26936 14832 26942 14844
rect 33594 14832 33600 14844
rect 33652 14832 33658 14884
rect 8110 14804 8116 14816
rect 7116 14776 7972 14804
rect 8071 14776 8116 14804
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 9217 14807 9275 14813
rect 9217 14773 9229 14807
rect 9263 14804 9275 14807
rect 9398 14804 9404 14816
rect 9263 14776 9404 14804
rect 9263 14773 9275 14776
rect 9217 14767 9275 14773
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 11793 14807 11851 14813
rect 11793 14773 11805 14807
rect 11839 14804 11851 14807
rect 18322 14804 18328 14816
rect 11839 14776 18328 14804
rect 11839 14773 11851 14776
rect 11793 14767 11851 14773
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 18509 14807 18567 14813
rect 18509 14804 18521 14807
rect 18472 14776 18521 14804
rect 18472 14764 18478 14776
rect 18509 14773 18521 14776
rect 18555 14773 18567 14807
rect 18509 14767 18567 14773
rect 18690 14764 18696 14816
rect 18748 14804 18754 14816
rect 19153 14807 19211 14813
rect 19153 14804 19165 14807
rect 18748 14776 19165 14804
rect 18748 14764 18754 14776
rect 19153 14773 19165 14776
rect 19199 14773 19211 14807
rect 19153 14767 19211 14773
rect 20162 14764 20168 14816
rect 20220 14804 20226 14816
rect 20622 14804 20628 14816
rect 20220 14776 20628 14804
rect 20220 14764 20226 14776
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 21361 14807 21419 14813
rect 21361 14773 21373 14807
rect 21407 14804 21419 14807
rect 27706 14804 27712 14816
rect 21407 14776 27712 14804
rect 21407 14773 21419 14776
rect 21361 14767 21419 14773
rect 27706 14764 27712 14776
rect 27764 14764 27770 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1857 14603 1915 14609
rect 1857 14569 1869 14603
rect 1903 14600 1915 14603
rect 2866 14600 2872 14612
rect 1903 14572 2872 14600
rect 1903 14569 1915 14572
rect 1857 14563 1915 14569
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 3053 14603 3111 14609
rect 3053 14569 3065 14603
rect 3099 14600 3111 14603
rect 3142 14600 3148 14612
rect 3099 14572 3148 14600
rect 3099 14569 3111 14572
rect 3053 14563 3111 14569
rect 3142 14560 3148 14572
rect 3200 14600 3206 14612
rect 4062 14600 4068 14612
rect 3200 14572 4068 14600
rect 3200 14560 3206 14572
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5353 14603 5411 14609
rect 5353 14600 5365 14603
rect 5316 14572 5365 14600
rect 5316 14560 5322 14572
rect 5353 14569 5365 14572
rect 5399 14569 5411 14603
rect 5353 14563 5411 14569
rect 5902 14560 5908 14612
rect 5960 14600 5966 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5960 14572 6009 14600
rect 5960 14560 5966 14572
rect 5997 14569 6009 14572
rect 6043 14569 6055 14603
rect 5997 14563 6055 14569
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 7926 14600 7932 14612
rect 6604 14572 7932 14600
rect 6604 14560 6610 14572
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8202 14600 8208 14612
rect 8163 14572 8208 14600
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 11241 14603 11299 14609
rect 11241 14569 11253 14603
rect 11287 14600 11299 14603
rect 11790 14600 11796 14612
rect 11287 14572 11796 14600
rect 11287 14569 11299 14572
rect 11241 14563 11299 14569
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 15105 14603 15163 14609
rect 15105 14569 15117 14603
rect 15151 14600 15163 14603
rect 16850 14600 16856 14612
rect 15151 14572 16856 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 17678 14560 17684 14612
rect 17736 14600 17742 14612
rect 24118 14600 24124 14612
rect 17736 14572 24124 14600
rect 17736 14560 17742 14572
rect 24118 14560 24124 14572
rect 24176 14560 24182 14612
rect 24578 14600 24584 14612
rect 24539 14572 24584 14600
rect 24578 14560 24584 14572
rect 24636 14560 24642 14612
rect 36538 14560 36544 14612
rect 36596 14600 36602 14612
rect 38105 14603 38163 14609
rect 38105 14600 38117 14603
rect 36596 14572 38117 14600
rect 36596 14560 36602 14572
rect 38105 14569 38117 14572
rect 38151 14569 38163 14603
rect 38105 14563 38163 14569
rect 3694 14492 3700 14544
rect 3752 14532 3758 14544
rect 3752 14504 13216 14532
rect 3752 14492 3758 14504
rect 7374 14464 7380 14476
rect 5920 14436 7380 14464
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 1728 14368 1777 14396
rect 1728 14356 1734 14368
rect 1765 14365 1777 14368
rect 1811 14365 1823 14399
rect 2406 14396 2412 14408
rect 2367 14368 2412 14396
rect 1765 14359 1823 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 3786 14396 3792 14408
rect 2639 14368 3792 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3936 14368 3985 14396
rect 3936 14356 3942 14368
rect 3973 14365 3985 14368
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14396 4675 14399
rect 5261 14399 5319 14405
rect 4663 14368 5212 14396
rect 4663 14365 4675 14368
rect 4617 14359 4675 14365
rect 4065 14331 4123 14337
rect 4065 14297 4077 14331
rect 4111 14328 4123 14331
rect 4798 14328 4804 14340
rect 4111 14300 4804 14328
rect 4111 14297 4123 14300
rect 4065 14291 4123 14297
rect 4798 14288 4804 14300
rect 4856 14288 4862 14340
rect 5184 14328 5212 14368
rect 5261 14365 5273 14399
rect 5307 14396 5319 14399
rect 5626 14396 5632 14408
rect 5307 14368 5632 14396
rect 5307 14365 5319 14368
rect 5261 14359 5319 14365
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 5920 14405 5948 14436
rect 7374 14424 7380 14436
rect 7432 14424 7438 14476
rect 9309 14467 9367 14473
rect 9309 14433 9321 14467
rect 9355 14464 9367 14467
rect 12526 14464 12532 14476
rect 9355 14436 12532 14464
rect 9355 14433 9367 14436
rect 9309 14427 9367 14433
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 13188 14464 13216 14504
rect 13262 14492 13268 14544
rect 13320 14532 13326 14544
rect 19242 14532 19248 14544
rect 13320 14504 19248 14532
rect 13320 14492 13326 14504
rect 19242 14492 19248 14504
rect 19300 14492 19306 14544
rect 20257 14535 20315 14541
rect 20257 14501 20269 14535
rect 20303 14532 20315 14535
rect 23658 14532 23664 14544
rect 20303 14504 23664 14532
rect 20303 14501 20315 14504
rect 20257 14495 20315 14501
rect 23658 14492 23664 14504
rect 23716 14492 23722 14544
rect 17586 14464 17592 14476
rect 13188 14436 17592 14464
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 17862 14424 17868 14476
rect 17920 14464 17926 14476
rect 18141 14467 18199 14473
rect 18141 14464 18153 14467
rect 17920 14436 18153 14464
rect 17920 14424 17926 14436
rect 18141 14433 18153 14436
rect 18187 14464 18199 14467
rect 18187 14436 20852 14464
rect 18187 14433 18199 14436
rect 18141 14427 18199 14433
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14365 5963 14399
rect 5905 14359 5963 14365
rect 7650 14356 7656 14408
rect 7708 14396 7714 14408
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 7708 14368 8125 14396
rect 7708 14356 7714 14368
rect 8113 14365 8125 14368
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 11112 14368 11161 14396
rect 11112 14356 11118 14368
rect 11149 14365 11161 14368
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 11698 14356 11704 14408
rect 11756 14396 11762 14408
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11756 14368 11805 14396
rect 11756 14356 11762 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 12342 14396 12348 14408
rect 11793 14359 11851 14365
rect 12268 14368 12348 14396
rect 6546 14328 6552 14340
rect 5184 14300 6552 14328
rect 6546 14288 6552 14300
rect 6604 14288 6610 14340
rect 6733 14331 6791 14337
rect 6733 14297 6745 14331
rect 6779 14297 6791 14331
rect 6733 14291 6791 14297
rect 6825 14331 6883 14337
rect 6825 14297 6837 14331
rect 6871 14328 6883 14331
rect 6914 14328 6920 14340
rect 6871 14300 6920 14328
rect 6871 14297 6883 14300
rect 6825 14291 6883 14297
rect 4706 14260 4712 14272
rect 4667 14232 4712 14260
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 6748 14260 6776 14291
rect 6914 14288 6920 14300
rect 6972 14288 6978 14340
rect 7374 14328 7380 14340
rect 7335 14300 7380 14328
rect 7374 14288 7380 14300
rect 7432 14288 7438 14340
rect 9398 14288 9404 14340
rect 9456 14328 9462 14340
rect 9456 14300 9501 14328
rect 9456 14288 9462 14300
rect 10226 14288 10232 14340
rect 10284 14328 10290 14340
rect 10321 14331 10379 14337
rect 10321 14328 10333 14331
rect 10284 14300 10333 14328
rect 10284 14288 10290 14300
rect 10321 14297 10333 14300
rect 10367 14297 10379 14331
rect 12268 14328 12296 14368
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 15010 14396 15016 14408
rect 14971 14368 15016 14396
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15286 14328 15292 14340
rect 10321 14291 10379 14297
rect 11716 14300 12296 14328
rect 12406 14300 15292 14328
rect 11716 14260 11744 14300
rect 11882 14260 11888 14272
rect 6748 14232 11744 14260
rect 11843 14232 11888 14260
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 12406 14260 12434 14300
rect 15286 14288 15292 14300
rect 15344 14288 15350 14340
rect 17678 14288 17684 14340
rect 17736 14328 17742 14340
rect 17865 14331 17923 14337
rect 17865 14328 17877 14331
rect 17736 14300 17877 14328
rect 17736 14288 17742 14300
rect 17865 14297 17877 14300
rect 17911 14297 17923 14331
rect 17865 14291 17923 14297
rect 17957 14331 18015 14337
rect 17957 14297 17969 14331
rect 18003 14328 18015 14331
rect 18690 14328 18696 14340
rect 18003 14300 18696 14328
rect 18003 14297 18015 14300
rect 17957 14291 18015 14297
rect 18690 14288 18696 14300
rect 18748 14288 18754 14340
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 19705 14331 19763 14337
rect 19705 14328 19717 14331
rect 19208 14300 19717 14328
rect 19208 14288 19214 14300
rect 19705 14297 19717 14300
rect 19751 14297 19763 14331
rect 19705 14291 19763 14297
rect 19797 14331 19855 14337
rect 19797 14297 19809 14331
rect 19843 14297 19855 14331
rect 20824 14328 20852 14436
rect 20990 14424 20996 14476
rect 21048 14464 21054 14476
rect 29822 14464 29828 14476
rect 21048 14436 29828 14464
rect 21048 14424 21054 14436
rect 29822 14424 29828 14436
rect 29880 14424 29886 14476
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21634 14396 21640 14408
rect 20956 14368 21640 14396
rect 20956 14356 20962 14368
rect 21634 14356 21640 14368
rect 21692 14396 21698 14408
rect 22462 14396 22468 14408
rect 21692 14368 22468 14396
rect 21692 14356 21698 14368
rect 22462 14356 22468 14368
rect 22520 14356 22526 14408
rect 24394 14356 24400 14408
rect 24452 14396 24458 14408
rect 24765 14399 24823 14405
rect 24765 14396 24777 14399
rect 24452 14368 24777 14396
rect 24452 14356 24458 14368
rect 24765 14365 24777 14368
rect 24811 14365 24823 14399
rect 38286 14396 38292 14408
rect 38247 14368 38292 14396
rect 24765 14359 24823 14365
rect 38286 14356 38292 14368
rect 38344 14356 38350 14408
rect 23566 14328 23572 14340
rect 20824 14300 23572 14328
rect 19797 14291 19855 14297
rect 12032 14232 12434 14260
rect 15304 14260 15332 14288
rect 19334 14260 19340 14272
rect 15304 14232 19340 14260
rect 12032 14220 12038 14232
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 19426 14220 19432 14272
rect 19484 14260 19490 14272
rect 19812 14260 19840 14291
rect 23566 14288 23572 14300
rect 23624 14288 23630 14340
rect 19484 14232 19840 14260
rect 22557 14263 22615 14269
rect 19484 14220 19490 14232
rect 22557 14229 22569 14263
rect 22603 14260 22615 14263
rect 23382 14260 23388 14272
rect 22603 14232 23388 14260
rect 22603 14229 22615 14232
rect 22557 14223 22615 14229
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 27614 14260 27620 14272
rect 27575 14232 27620 14260
rect 27614 14220 27620 14232
rect 27672 14220 27678 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 5350 14056 5356 14068
rect 4212 14028 5356 14056
rect 4212 14016 4218 14028
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 7282 14056 7288 14068
rect 7195 14028 7288 14056
rect 7282 14016 7288 14028
rect 7340 14056 7346 14068
rect 8110 14056 8116 14068
rect 7340 14028 8116 14056
rect 7340 14016 7346 14028
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8389 14059 8447 14065
rect 8389 14025 8401 14059
rect 8435 14056 8447 14059
rect 9858 14056 9864 14068
rect 8435 14028 9864 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10336 14028 12756 14056
rect 2501 13991 2559 13997
rect 2501 13957 2513 13991
rect 2547 13988 2559 13991
rect 4706 13988 4712 14000
rect 2547 13960 4712 13988
rect 2547 13957 2559 13960
rect 2501 13951 2559 13957
rect 4706 13948 4712 13960
rect 4764 13948 4770 14000
rect 6564 13960 10180 13988
rect 1578 13920 1584 13932
rect 1539 13892 1584 13920
rect 1578 13880 1584 13892
rect 1636 13880 1642 13932
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 4120 13892 4445 13920
rect 4120 13880 4126 13892
rect 4433 13889 4445 13892
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 5166 13880 5172 13932
rect 5224 13920 5230 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 5224 13892 5273 13920
rect 5224 13880 5230 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5718 13920 5724 13932
rect 5631 13892 5724 13920
rect 5261 13883 5319 13889
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13852 2467 13855
rect 2590 13852 2596 13864
rect 2455 13824 2596 13852
rect 2455 13821 2467 13824
rect 2409 13815 2467 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3421 13855 3479 13861
rect 3421 13821 3433 13855
rect 3467 13852 3479 13855
rect 4154 13852 4160 13864
rect 3467 13824 4160 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 4706 13852 4712 13864
rect 4571 13824 4712 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 4706 13812 4712 13824
rect 4764 13812 4770 13864
rect 5276 13852 5304 13883
rect 5718 13880 5724 13892
rect 5776 13920 5782 13932
rect 5994 13920 6000 13932
rect 5776 13892 6000 13920
rect 5776 13880 5782 13892
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 6564 13920 6592 13960
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 6564 13892 6653 13920
rect 6641 13889 6653 13892
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 6748 13892 7052 13920
rect 5350 13852 5356 13864
rect 5263 13824 5356 13852
rect 5350 13812 5356 13824
rect 5408 13852 5414 13864
rect 5408 13840 6684 13852
rect 6748 13840 6776 13892
rect 5408 13824 6776 13840
rect 5408 13812 5414 13824
rect 6656 13812 6776 13824
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 7024 13852 7052 13892
rect 7098 13880 7104 13932
rect 7156 13920 7162 13932
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7156 13892 7757 13920
rect 7156 13880 7162 13892
rect 7745 13889 7757 13892
rect 7791 13920 7803 13923
rect 8573 13923 8631 13929
rect 8573 13920 8585 13923
rect 7791 13892 8585 13920
rect 7791 13889 7803 13892
rect 7745 13883 7803 13889
rect 8573 13889 8585 13892
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9950 13920 9956 13932
rect 9723 13892 9956 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 7650 13852 7656 13864
rect 6880 13824 6925 13852
rect 7024 13824 7656 13852
rect 6880 13812 6886 13824
rect 7650 13812 7656 13824
rect 7708 13812 7714 13864
rect 7834 13852 7840 13864
rect 7795 13824 7840 13852
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8018 13812 8024 13864
rect 8076 13852 8082 13864
rect 8076 13824 8340 13852
rect 8076 13812 8082 13824
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 8312 13784 8340 13824
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 9232 13852 9260 13883
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 8444 13824 9260 13852
rect 10152 13852 10180 13960
rect 10336 13929 10364 14028
rect 10413 13991 10471 13997
rect 10413 13957 10425 13991
rect 10459 13988 10471 13991
rect 11885 13991 11943 13997
rect 11885 13988 11897 13991
rect 10459 13960 11897 13988
rect 10459 13957 10471 13960
rect 10413 13951 10471 13957
rect 11885 13957 11897 13960
rect 11931 13957 11943 13991
rect 11885 13951 11943 13957
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 10778 13880 10784 13932
rect 10836 13920 10842 13932
rect 10962 13920 10968 13932
rect 10836 13892 10968 13920
rect 10836 13880 10842 13892
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13920 11115 13923
rect 11330 13920 11336 13932
rect 11103 13892 11336 13920
rect 11103 13889 11115 13892
rect 11057 13883 11115 13889
rect 11330 13880 11336 13892
rect 11388 13880 11394 13932
rect 12728 13920 12756 14028
rect 12820 14028 16160 14056
rect 12820 13997 12848 14028
rect 12805 13991 12863 13997
rect 12805 13957 12817 13991
rect 12851 13957 12863 13991
rect 12805 13951 12863 13957
rect 12912 13960 13400 13988
rect 12912 13920 12940 13960
rect 13262 13920 13268 13932
rect 12728 13892 12940 13920
rect 13223 13892 13268 13920
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 13372 13920 13400 13960
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 15381 13991 15439 13997
rect 15381 13988 15393 13991
rect 13872 13960 15393 13988
rect 13872 13948 13878 13960
rect 15381 13957 15393 13960
rect 15427 13957 15439 13991
rect 16132 13988 16160 14028
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 20714 14056 20720 14068
rect 16264 14028 20024 14056
rect 16264 14016 16270 14028
rect 17126 13988 17132 14000
rect 16132 13960 17132 13988
rect 15381 13951 15439 13957
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 18414 13988 18420 14000
rect 18375 13960 18420 13988
rect 18414 13948 18420 13960
rect 18472 13948 18478 14000
rect 19242 13948 19248 14000
rect 19300 13988 19306 14000
rect 19886 13988 19892 14000
rect 19300 13960 19892 13988
rect 19300 13948 19306 13960
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 19996 13997 20024 14028
rect 20088 14028 20720 14056
rect 19981 13991 20039 13997
rect 19981 13957 19993 13991
rect 20027 13957 20039 13991
rect 19981 13951 20039 13957
rect 13998 13920 14004 13932
rect 13372 13892 14004 13920
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13889 14611 13923
rect 17862 13920 17868 13932
rect 14553 13883 14611 13889
rect 16316 13892 17868 13920
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 10152 13824 10916 13852
rect 8444 13812 8450 13824
rect 9033 13787 9091 13793
rect 9033 13784 9045 13787
rect 5500 13756 8248 13784
rect 8312 13756 9045 13784
rect 5500 13744 5506 13756
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 5074 13716 5080 13728
rect 5035 13688 5080 13716
rect 5074 13676 5080 13688
rect 5132 13676 5138 13728
rect 5813 13719 5871 13725
rect 5813 13685 5825 13719
rect 5859 13716 5871 13719
rect 6822 13716 6828 13728
rect 5859 13688 6828 13716
rect 5859 13685 5871 13688
rect 5813 13679 5871 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 8220 13716 8248 13756
rect 9033 13753 9045 13756
rect 9079 13753 9091 13787
rect 10888 13784 10916 13824
rect 11164 13824 11805 13852
rect 11164 13784 11192 13824
rect 11793 13821 11805 13824
rect 11839 13852 11851 13855
rect 11882 13852 11888 13864
rect 11839 13824 11888 13852
rect 11839 13821 11851 13824
rect 11793 13815 11851 13821
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 13722 13852 13728 13864
rect 12860 13824 13728 13852
rect 12860 13812 12866 13824
rect 13722 13812 13728 13824
rect 13780 13852 13786 13864
rect 14568 13852 14596 13883
rect 13780 13824 14596 13852
rect 14645 13855 14703 13861
rect 13780 13812 13786 13824
rect 14645 13821 14657 13855
rect 14691 13852 14703 13855
rect 15010 13852 15016 13864
rect 14691 13824 15016 13852
rect 14691 13821 14703 13824
rect 14645 13815 14703 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15286 13852 15292 13864
rect 15247 13824 15292 13852
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 16316 13861 16344 13892
rect 17862 13880 17868 13892
rect 17920 13880 17926 13932
rect 18969 13923 19027 13929
rect 18969 13889 18981 13923
rect 19015 13920 19027 13923
rect 20088 13920 20116 14028
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 24394 14056 24400 14068
rect 24355 14028 24400 14056
rect 24394 14016 24400 14028
rect 24452 14016 24458 14068
rect 20165 13991 20223 13997
rect 20165 13957 20177 13991
rect 20211 13988 20223 13991
rect 26878 13988 26884 14000
rect 20211 13960 26884 13988
rect 20211 13957 20223 13960
rect 20165 13951 20223 13957
rect 26878 13948 26884 13960
rect 26936 13948 26942 14000
rect 27614 13988 27620 14000
rect 27575 13960 27620 13988
rect 27614 13948 27620 13960
rect 27672 13948 27678 14000
rect 27706 13948 27712 14000
rect 27764 13988 27770 14000
rect 27764 13960 27809 13988
rect 27764 13948 27770 13960
rect 19015 13910 19288 13920
rect 19015 13892 19334 13910
rect 19015 13889 19027 13892
rect 18969 13883 19027 13889
rect 19260 13882 19334 13892
rect 16301 13855 16359 13861
rect 16301 13821 16313 13855
rect 16347 13821 16359 13855
rect 16301 13815 16359 13821
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 18325 13855 18383 13861
rect 18325 13852 18337 13855
rect 16540 13824 18337 13852
rect 16540 13812 16546 13824
rect 18325 13821 18337 13824
rect 18371 13852 18383 13855
rect 19150 13852 19156 13864
rect 18371 13824 19156 13852
rect 18371 13821 18383 13824
rect 18325 13815 18383 13821
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 19306 13852 19334 13882
rect 19812 13892 20116 13920
rect 20625 13923 20683 13929
rect 19812 13852 19840 13892
rect 20625 13889 20637 13923
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 19306 13824 19840 13852
rect 19886 13812 19892 13864
rect 19944 13852 19950 13864
rect 20640 13852 20668 13883
rect 22462 13880 22468 13932
rect 22520 13920 22526 13932
rect 24578 13920 24584 13932
rect 22520 13892 24584 13920
rect 22520 13880 22526 13892
rect 24578 13880 24584 13892
rect 24636 13880 24642 13932
rect 19944 13824 20668 13852
rect 20717 13855 20775 13861
rect 19944 13812 19950 13824
rect 20717 13821 20729 13855
rect 20763 13852 20775 13855
rect 26142 13852 26148 13864
rect 20763 13824 26148 13852
rect 20763 13821 20775 13824
rect 20717 13815 20775 13821
rect 26142 13812 26148 13824
rect 26200 13812 26206 13864
rect 27706 13812 27712 13864
rect 27764 13852 27770 13864
rect 27982 13852 27988 13864
rect 27764 13824 27988 13852
rect 27764 13812 27770 13824
rect 27982 13812 27988 13824
rect 28040 13812 28046 13864
rect 9033 13747 9091 13753
rect 9140 13756 10824 13784
rect 10888 13756 11192 13784
rect 9140 13716 9168 13756
rect 9766 13716 9772 13728
rect 8220 13688 9168 13716
rect 9727 13688 9772 13716
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 10796 13716 10824 13756
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 12158 13784 12164 13796
rect 11296 13756 12164 13784
rect 11296 13744 11302 13756
rect 12158 13744 12164 13756
rect 12216 13744 12222 13796
rect 17954 13784 17960 13796
rect 12406 13756 17960 13784
rect 12406 13716 12434 13756
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 18046 13744 18052 13796
rect 18104 13784 18110 13796
rect 18104 13756 31754 13784
rect 18104 13744 18110 13756
rect 13354 13716 13360 13728
rect 10796 13688 12434 13716
rect 13315 13688 13360 13716
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 22278 13716 22284 13728
rect 15712 13688 22284 13716
rect 15712 13676 15718 13688
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 31726 13716 31754 13756
rect 38194 13716 38200 13728
rect 31726 13688 38200 13716
rect 38194 13676 38200 13688
rect 38252 13676 38258 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2958 13472 2964 13524
rect 3016 13512 3022 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 3016 13484 4077 13512
rect 3016 13472 3022 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 5353 13515 5411 13521
rect 5353 13481 5365 13515
rect 5399 13512 5411 13515
rect 6730 13512 6736 13524
rect 5399 13484 6736 13512
rect 5399 13481 5411 13484
rect 5353 13475 5411 13481
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 7248 13484 12081 13512
rect 7248 13472 7254 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 12342 13472 12348 13524
rect 12400 13512 12406 13524
rect 12710 13512 12716 13524
rect 12400 13484 12716 13512
rect 12400 13472 12406 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 12805 13515 12863 13521
rect 12805 13481 12817 13515
rect 12851 13512 12863 13515
rect 13814 13512 13820 13524
rect 12851 13484 13820 13512
rect 12851 13481 12863 13484
rect 12805 13475 12863 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 17218 13512 17224 13524
rect 14384 13484 17224 13512
rect 7282 13444 7288 13456
rect 6748 13416 7288 13444
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13376 2099 13379
rect 2406 13376 2412 13388
rect 2087 13348 2412 13376
rect 2087 13345 2099 13348
rect 2041 13339 2099 13345
rect 2406 13336 2412 13348
rect 2464 13336 2470 13388
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 3418 13376 3424 13388
rect 2832 13348 2877 13376
rect 3379 13348 3424 13376
rect 2832 13336 2838 13348
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 6748 13385 6776 13416
rect 7282 13404 7288 13416
rect 7340 13404 7346 13456
rect 14384 13444 14412 13484
rect 17218 13472 17224 13484
rect 17276 13512 17282 13524
rect 30374 13512 30380 13524
rect 17276 13484 30380 13512
rect 17276 13472 17282 13484
rect 30374 13472 30380 13484
rect 30432 13512 30438 13524
rect 30558 13512 30564 13524
rect 30432 13484 30564 13512
rect 30432 13472 30438 13484
rect 30558 13472 30564 13484
rect 30616 13472 30622 13524
rect 17034 13444 17040 13456
rect 9692 13416 14412 13444
rect 14476 13416 17040 13444
rect 6733 13379 6791 13385
rect 6733 13345 6745 13379
rect 6779 13345 6791 13379
rect 7006 13376 7012 13388
rect 6967 13348 7012 13376
rect 6733 13339 6791 13345
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 9692 13385 9720 13416
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13345 9735 13379
rect 10226 13376 10232 13388
rect 10187 13348 10232 13376
rect 9677 13339 9735 13345
rect 10226 13336 10232 13348
rect 10284 13376 10290 13388
rect 10502 13376 10508 13388
rect 10284 13348 10508 13376
rect 10284 13336 10290 13348
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 14476 13376 14504 13416
rect 17034 13404 17040 13416
rect 17092 13444 17098 13456
rect 18046 13444 18052 13456
rect 17092 13416 18052 13444
rect 17092 13404 17098 13416
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 23198 13404 23204 13456
rect 23256 13404 23262 13456
rect 26326 13404 26332 13456
rect 26384 13444 26390 13456
rect 26384 13416 38056 13444
rect 26384 13404 26390 13416
rect 12268 13348 14504 13376
rect 14553 13379 14611 13385
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4614 13308 4620 13320
rect 4019 13280 4620 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4614 13268 4620 13280
rect 4672 13308 4678 13320
rect 4801 13311 4859 13317
rect 4801 13308 4813 13311
rect 4672 13280 4813 13308
rect 4672 13268 4678 13280
rect 4801 13277 4813 13280
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5537 13311 5595 13317
rect 5537 13308 5549 13311
rect 5132 13280 5549 13308
rect 5132 13268 5138 13280
rect 5537 13277 5549 13280
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 5997 13311 6055 13317
rect 5997 13277 6009 13311
rect 6043 13308 6055 13311
rect 8386 13308 8392 13320
rect 6043 13280 6592 13308
rect 8347 13280 8392 13308
rect 6043 13277 6055 13280
rect 5997 13271 6055 13277
rect 2869 13243 2927 13249
rect 2869 13209 2881 13243
rect 2915 13209 2927 13243
rect 2869 13203 2927 13209
rect 2884 13172 2912 13203
rect 2958 13172 2964 13184
rect 2884 13144 2964 13172
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 4614 13172 4620 13184
rect 4575 13144 4620 13172
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 6086 13172 6092 13184
rect 6047 13144 6092 13172
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 6564 13172 6592 13280
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 12158 13308 12164 13320
rect 11563 13280 12164 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 6880 13212 6925 13240
rect 6880 13200 6886 13212
rect 9766 13200 9772 13252
rect 9824 13240 9830 13252
rect 9824 13212 9869 13240
rect 9824 13200 9830 13212
rect 9950 13200 9956 13252
rect 10008 13240 10014 13252
rect 10686 13240 10692 13252
rect 10008 13212 10692 13240
rect 10008 13200 10014 13212
rect 10686 13200 10692 13212
rect 10744 13200 10750 13252
rect 11440 13240 11468 13271
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 12268 13317 12296 13348
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15930 13376 15936 13388
rect 14599 13348 15936 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15930 13336 15936 13348
rect 15988 13376 15994 13388
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 15988 13348 16405 13376
rect 15988 13336 15994 13348
rect 16393 13345 16405 13348
rect 16439 13345 16451 13379
rect 16666 13376 16672 13388
rect 16627 13348 16672 13376
rect 16393 13339 16451 13345
rect 16666 13336 16672 13348
rect 16724 13376 16730 13388
rect 23216 13376 23244 13404
rect 23293 13379 23351 13385
rect 23293 13376 23305 13379
rect 16724 13348 19334 13376
rect 23216 13348 23305 13376
rect 16724 13336 16730 13348
rect 12253 13311 12311 13317
rect 12253 13277 12265 13311
rect 12299 13277 12311 13311
rect 12710 13308 12716 13320
rect 12671 13280 12716 13308
rect 12253 13271 12311 13277
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 13538 13308 13544 13320
rect 13499 13280 13544 13308
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13308 14519 13311
rect 14642 13308 14648 13320
rect 14507 13280 14648 13308
rect 14507 13277 14519 13280
rect 14461 13271 14519 13277
rect 14642 13268 14648 13280
rect 14700 13268 14706 13320
rect 15654 13308 15660 13320
rect 15615 13280 15660 13308
rect 15654 13268 15660 13280
rect 15712 13268 15718 13320
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17489 13313 17547 13319
rect 17489 13310 17501 13313
rect 17420 13308 17501 13310
rect 17092 13282 17501 13308
rect 17092 13280 17448 13282
rect 17092 13268 17098 13280
rect 17489 13279 17501 13282
rect 17535 13279 17547 13313
rect 19306 13308 19334 13348
rect 23293 13345 23305 13348
rect 23339 13345 23351 13379
rect 23293 13339 23351 13345
rect 30101 13379 30159 13385
rect 30101 13345 30113 13379
rect 30147 13376 30159 13379
rect 30466 13376 30472 13388
rect 30147 13348 30472 13376
rect 30147 13345 30159 13348
rect 30101 13339 30159 13345
rect 30466 13336 30472 13348
rect 30524 13336 30530 13388
rect 30558 13336 30564 13388
rect 30616 13376 30622 13388
rect 30616 13348 30661 13376
rect 30616 13336 30622 13348
rect 21450 13308 21456 13320
rect 19306 13280 21456 13308
rect 17489 13273 17547 13279
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 37274 13308 37280 13320
rect 37235 13280 37280 13308
rect 37274 13268 37280 13280
rect 37332 13268 37338 13320
rect 38028 13317 38056 13416
rect 38013 13311 38071 13317
rect 38013 13277 38025 13311
rect 38059 13277 38071 13311
rect 38013 13271 38071 13277
rect 13262 13240 13268 13252
rect 11440 13212 13268 13240
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13633 13243 13691 13249
rect 13633 13209 13645 13243
rect 13679 13240 13691 13243
rect 14734 13240 14740 13252
rect 13679 13212 14740 13240
rect 13679 13209 13691 13212
rect 13633 13203 13691 13209
rect 14734 13200 14740 13212
rect 14792 13200 14798 13252
rect 16485 13243 16543 13249
rect 16485 13209 16497 13243
rect 16531 13209 16543 13243
rect 16485 13203 16543 13209
rect 7466 13172 7472 13184
rect 6564 13144 7472 13172
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 8478 13172 8484 13184
rect 8439 13144 8484 13172
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 8662 13132 8668 13184
rect 8720 13172 8726 13184
rect 12342 13172 12348 13184
rect 8720 13144 12348 13172
rect 8720 13132 8726 13144
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 15749 13175 15807 13181
rect 15749 13141 15761 13175
rect 15795 13172 15807 13175
rect 16500 13172 16528 13203
rect 17310 13200 17316 13252
rect 17368 13240 17374 13252
rect 20346 13240 20352 13252
rect 17368 13212 20352 13240
rect 17368 13200 17374 13212
rect 20346 13200 20352 13212
rect 20404 13240 20410 13252
rect 20404 13212 22094 13240
rect 20404 13200 20410 13212
rect 17586 13172 17592 13184
rect 15795 13144 16528 13172
rect 17547 13144 17592 13172
rect 15795 13141 15807 13144
rect 15749 13135 15807 13141
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 17678 13132 17684 13184
rect 17736 13172 17742 13184
rect 20806 13172 20812 13184
rect 17736 13144 20812 13172
rect 17736 13132 17742 13144
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 22066 13172 22094 13212
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 23937 13243 23995 13249
rect 23440 13212 23485 13240
rect 23440 13200 23446 13212
rect 23937 13209 23949 13243
rect 23983 13240 23995 13243
rect 25314 13240 25320 13252
rect 23983 13212 25320 13240
rect 23983 13209 23995 13212
rect 23937 13203 23995 13209
rect 25314 13200 25320 13212
rect 25372 13200 25378 13252
rect 26142 13200 26148 13252
rect 26200 13240 26206 13252
rect 30193 13243 30251 13249
rect 30193 13240 30205 13243
rect 26200 13212 30205 13240
rect 26200 13200 26206 13212
rect 30193 13209 30205 13212
rect 30239 13209 30251 13243
rect 30193 13203 30251 13209
rect 26602 13172 26608 13184
rect 22066 13144 26608 13172
rect 26602 13132 26608 13144
rect 26660 13132 26666 13184
rect 37366 13172 37372 13184
rect 37327 13144 37372 13172
rect 37366 13132 37372 13144
rect 37424 13132 37430 13184
rect 38194 13172 38200 13184
rect 38155 13144 38200 13172
rect 38194 13132 38200 13144
rect 38252 13132 38258 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 2409 12971 2467 12977
rect 2409 12937 2421 12971
rect 2455 12968 2467 12971
rect 2958 12968 2964 12980
rect 2455 12940 2964 12968
rect 2455 12937 2467 12940
rect 2409 12931 2467 12937
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3145 12971 3203 12977
rect 3145 12968 3157 12971
rect 3108 12940 3157 12968
rect 3108 12928 3114 12940
rect 3145 12937 3157 12940
rect 3191 12937 3203 12971
rect 3145 12931 3203 12937
rect 3789 12971 3847 12977
rect 3789 12937 3801 12971
rect 3835 12968 3847 12971
rect 4890 12968 4896 12980
rect 3835 12940 4896 12968
rect 3835 12937 3847 12940
rect 3789 12931 3847 12937
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 10594 12968 10600 12980
rect 8352 12940 10600 12968
rect 8352 12928 8358 12940
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 13538 12968 13544 12980
rect 10744 12940 13544 12968
rect 10744 12928 10750 12940
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17000 12940 19932 12968
rect 17000 12928 17006 12940
rect 1670 12860 1676 12912
rect 1728 12900 1734 12912
rect 4709 12903 4767 12909
rect 1728 12872 3096 12900
rect 1728 12860 1734 12872
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 2038 12832 2044 12844
rect 1627 12804 2044 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2498 12832 2504 12844
rect 2363 12804 2504 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3068 12841 3096 12872
rect 4709 12869 4721 12903
rect 4755 12900 4767 12903
rect 4798 12900 4804 12912
rect 4755 12872 4804 12900
rect 4755 12869 4767 12872
rect 4709 12863 4767 12869
rect 4798 12860 4804 12872
rect 4856 12860 4862 12912
rect 6638 12860 6644 12912
rect 6696 12900 6702 12912
rect 7561 12903 7619 12909
rect 7561 12900 7573 12903
rect 6696 12872 7573 12900
rect 6696 12860 6702 12872
rect 7561 12869 7573 12872
rect 7607 12869 7619 12903
rect 7561 12863 7619 12869
rect 10134 12860 10140 12912
rect 10192 12900 10198 12912
rect 10229 12903 10287 12909
rect 10229 12900 10241 12903
rect 10192 12872 10241 12900
rect 10192 12860 10198 12872
rect 10229 12869 10241 12872
rect 10275 12869 10287 12903
rect 10229 12863 10287 12869
rect 12345 12903 12403 12909
rect 12345 12869 12357 12903
rect 12391 12900 12403 12903
rect 13354 12900 13360 12912
rect 12391 12872 13360 12900
rect 12391 12869 12403 12872
rect 12345 12863 12403 12869
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 17770 12860 17776 12912
rect 17828 12900 17834 12912
rect 17865 12903 17923 12909
rect 17865 12900 17877 12903
rect 17828 12872 17877 12900
rect 17828 12860 17834 12872
rect 17865 12869 17877 12872
rect 17911 12869 17923 12903
rect 17865 12863 17923 12869
rect 18785 12903 18843 12909
rect 18785 12869 18797 12903
rect 18831 12900 18843 12903
rect 19058 12900 19064 12912
rect 18831 12872 19064 12900
rect 18831 12869 18843 12872
rect 18785 12863 18843 12869
rect 19058 12860 19064 12872
rect 19116 12860 19122 12912
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 3099 12804 3709 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 6604 12804 6745 12832
rect 6604 12792 6610 12804
rect 6733 12801 6745 12804
rect 6779 12801 6791 12835
rect 9950 12832 9956 12844
rect 6733 12795 6791 12801
rect 8772 12804 9956 12832
rect 2590 12724 2596 12776
rect 2648 12764 2654 12776
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 2648 12736 4629 12764
rect 2648 12724 2654 12736
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 5442 12764 5448 12776
rect 5403 12736 5448 12764
rect 4617 12727 4675 12733
rect 5442 12724 5448 12736
rect 5500 12764 5506 12776
rect 7377 12767 7435 12773
rect 7377 12764 7389 12767
rect 5500 12736 7389 12764
rect 5500 12724 5506 12736
rect 7377 12733 7389 12736
rect 7423 12733 7435 12767
rect 8294 12764 8300 12776
rect 8255 12736 8300 12764
rect 7377 12727 7435 12733
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 8772 12696 8800 12804
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 13722 12832 13728 12844
rect 13683 12804 13728 12832
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 17310 12832 17316 12844
rect 15488 12804 17316 12832
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 4948 12668 8800 12696
rect 9968 12736 10149 12764
rect 4948 12656 4954 12668
rect 1762 12628 1768 12640
rect 1723 12600 1768 12628
rect 1762 12588 1768 12600
rect 1820 12588 1826 12640
rect 6825 12631 6883 12637
rect 6825 12597 6837 12631
rect 6871 12628 6883 12631
rect 8110 12628 8116 12640
rect 6871 12600 8116 12628
rect 6871 12597 6883 12600
rect 6825 12591 6883 12597
rect 8110 12588 8116 12600
rect 8168 12588 8174 12640
rect 9968 12628 9996 12736
rect 10137 12733 10149 12736
rect 10183 12733 10195 12767
rect 10502 12764 10508 12776
rect 10463 12736 10508 12764
rect 10137 12727 10195 12733
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 11422 12724 11428 12776
rect 11480 12764 11486 12776
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 11480 12736 12265 12764
rect 11480 12724 11486 12736
rect 12253 12733 12265 12736
rect 12299 12733 12311 12767
rect 12526 12764 12532 12776
rect 12487 12736 12532 12764
rect 12253 12727 12311 12733
rect 12526 12724 12532 12736
rect 12584 12764 12590 12776
rect 15488 12764 15516 12804
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 19904 12841 19932 12940
rect 23106 12928 23112 12980
rect 23164 12968 23170 12980
rect 25869 12971 25927 12977
rect 25869 12968 25881 12971
rect 23164 12940 25881 12968
rect 23164 12928 23170 12940
rect 25869 12937 25881 12940
rect 25915 12937 25927 12971
rect 25869 12931 25927 12937
rect 23290 12860 23296 12912
rect 23348 12900 23354 12912
rect 23385 12903 23443 12909
rect 23385 12900 23397 12903
rect 23348 12872 23397 12900
rect 23348 12860 23354 12872
rect 23385 12869 23397 12872
rect 23431 12869 23443 12903
rect 23385 12863 23443 12869
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 22005 12835 22063 12841
rect 22005 12801 22017 12835
rect 22051 12801 22063 12835
rect 25774 12832 25780 12844
rect 25735 12804 25780 12832
rect 22005 12795 22063 12801
rect 12584 12736 15516 12764
rect 12584 12724 12590 12736
rect 15562 12724 15568 12776
rect 15620 12764 15626 12776
rect 17586 12764 17592 12776
rect 15620 12736 17592 12764
rect 15620 12724 15626 12736
rect 17586 12724 17592 12736
rect 17644 12764 17650 12776
rect 17773 12767 17831 12773
rect 17773 12764 17785 12767
rect 17644 12736 17785 12764
rect 17644 12724 17650 12736
rect 17773 12733 17785 12736
rect 17819 12733 17831 12767
rect 22020 12764 22048 12795
rect 25774 12792 25780 12804
rect 25832 12792 25838 12844
rect 38010 12832 38016 12844
rect 37971 12804 38016 12832
rect 38010 12792 38016 12804
rect 38068 12792 38074 12844
rect 23290 12764 23296 12776
rect 17773 12727 17831 12733
rect 18892 12736 22048 12764
rect 23251 12736 23296 12764
rect 10594 12656 10600 12708
rect 10652 12696 10658 12708
rect 17678 12696 17684 12708
rect 10652 12668 17684 12696
rect 10652 12656 10658 12668
rect 17678 12656 17684 12668
rect 17736 12656 17742 12708
rect 17862 12656 17868 12708
rect 17920 12696 17926 12708
rect 18892 12696 18920 12736
rect 23290 12724 23296 12736
rect 23348 12724 23354 12776
rect 23566 12764 23572 12776
rect 23527 12736 23572 12764
rect 23566 12724 23572 12736
rect 23624 12724 23630 12776
rect 24854 12696 24860 12708
rect 17920 12668 18920 12696
rect 18984 12668 24860 12696
rect 17920 12656 17926 12668
rect 12250 12628 12256 12640
rect 9968 12600 12256 12628
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 13817 12631 13875 12637
rect 13817 12628 13829 12631
rect 12768 12600 13829 12628
rect 12768 12588 12774 12600
rect 13817 12597 13829 12600
rect 13863 12597 13875 12631
rect 13817 12591 13875 12597
rect 14642 12588 14648 12640
rect 14700 12628 14706 12640
rect 18984 12628 19012 12668
rect 24854 12656 24860 12668
rect 24912 12656 24918 12708
rect 14700 12600 19012 12628
rect 19981 12631 20039 12637
rect 14700 12588 14706 12600
rect 19981 12597 19993 12631
rect 20027 12628 20039 12631
rect 20070 12628 20076 12640
rect 20027 12600 20076 12628
rect 20027 12597 20039 12600
rect 19981 12591 20039 12597
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 38194 12628 38200 12640
rect 22152 12600 22197 12628
rect 38155 12600 38200 12628
rect 22152 12588 22158 12600
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 2130 12424 2136 12436
rect 2087 12396 2136 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 3786 12384 3792 12436
rect 3844 12424 3850 12436
rect 3973 12427 4031 12433
rect 3973 12424 3985 12427
rect 3844 12396 3985 12424
rect 3844 12384 3850 12396
rect 3973 12393 3985 12396
rect 4019 12393 4031 12427
rect 3973 12387 4031 12393
rect 6546 12384 6552 12436
rect 6604 12424 6610 12436
rect 7009 12427 7067 12433
rect 7009 12424 7021 12427
rect 6604 12396 7021 12424
rect 6604 12384 6610 12396
rect 7009 12393 7021 12396
rect 7055 12393 7067 12427
rect 16666 12424 16672 12436
rect 7009 12387 7067 12393
rect 7852 12396 16672 12424
rect 2590 12316 2596 12368
rect 2648 12356 2654 12368
rect 4890 12356 4896 12368
rect 2648 12328 4896 12356
rect 2648 12316 2654 12328
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 7558 12356 7564 12368
rect 6012 12328 7564 12356
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 3145 12291 3203 12297
rect 3145 12288 3157 12291
rect 2832 12260 3157 12288
rect 2832 12248 2838 12260
rect 3145 12257 3157 12260
rect 3191 12257 3203 12291
rect 3145 12251 3203 12257
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 5718 12288 5724 12300
rect 3568 12260 5724 12288
rect 3568 12248 3574 12260
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 1670 12180 1676 12232
rect 1728 12220 1734 12232
rect 1949 12223 2007 12229
rect 1949 12220 1961 12223
rect 1728 12192 1961 12220
rect 1728 12180 1734 12192
rect 1949 12189 1961 12192
rect 1995 12189 2007 12223
rect 1949 12183 2007 12189
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4614 12220 4620 12232
rect 4203 12192 4620 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4724 12152 4752 12183
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 6012 12229 6040 12328
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 6086 12248 6092 12300
rect 6144 12288 6150 12300
rect 6825 12291 6883 12297
rect 6825 12288 6837 12291
rect 6144 12260 6837 12288
rect 6144 12248 6150 12260
rect 6825 12257 6837 12260
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 5316 12192 5365 12220
rect 5316 12180 5322 12192
rect 5353 12189 5365 12192
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12189 6055 12223
rect 5997 12183 6055 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 7852 12220 7880 12396
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 17126 12384 17132 12436
rect 17184 12424 17190 12436
rect 26050 12424 26056 12436
rect 17184 12396 26056 12424
rect 17184 12384 17190 12396
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 37829 12427 37887 12433
rect 37829 12393 37841 12427
rect 37875 12424 37887 12427
rect 38010 12424 38016 12436
rect 37875 12396 38016 12424
rect 37875 12393 37887 12396
rect 37829 12387 37887 12393
rect 38010 12384 38016 12396
rect 38068 12384 38074 12436
rect 8294 12356 8300 12368
rect 8255 12328 8300 12356
rect 8294 12316 8300 12328
rect 8352 12316 8358 12368
rect 10318 12316 10324 12368
rect 10376 12356 10382 12368
rect 12158 12356 12164 12368
rect 10376 12328 12164 12356
rect 10376 12316 10382 12328
rect 12158 12316 12164 12328
rect 12216 12316 12222 12368
rect 17494 12356 17500 12368
rect 12406 12328 17500 12356
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8478 12288 8484 12300
rect 7975 12260 8484 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8478 12248 8484 12260
rect 8536 12288 8542 12300
rect 9217 12291 9275 12297
rect 9217 12288 9229 12291
rect 8536 12260 9229 12288
rect 8536 12248 8542 12260
rect 9217 12257 9229 12260
rect 9263 12257 9275 12291
rect 9217 12251 9275 12257
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 9677 12291 9735 12297
rect 9677 12288 9689 12291
rect 9548 12260 9689 12288
rect 9548 12248 9554 12260
rect 9677 12257 9689 12260
rect 9723 12288 9735 12291
rect 12406 12288 12434 12328
rect 17494 12316 17500 12328
rect 17552 12316 17558 12368
rect 18138 12316 18144 12368
rect 18196 12356 18202 12368
rect 20717 12359 20775 12365
rect 20717 12356 20729 12359
rect 18196 12328 20729 12356
rect 18196 12316 18202 12328
rect 20717 12325 20729 12328
rect 20763 12356 20775 12359
rect 24302 12356 24308 12368
rect 20763 12328 24308 12356
rect 20763 12325 20775 12328
rect 20717 12319 20775 12325
rect 24302 12316 24308 12328
rect 24360 12316 24366 12368
rect 15930 12288 15936 12300
rect 9723 12260 12434 12288
rect 15891 12260 15936 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 16945 12291 17003 12297
rect 16945 12257 16957 12291
rect 16991 12288 17003 12291
rect 17126 12288 17132 12300
rect 16991 12260 17132 12288
rect 16991 12257 17003 12260
rect 16945 12251 17003 12257
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 21913 12291 21971 12297
rect 21913 12257 21925 12291
rect 21959 12288 21971 12291
rect 22738 12288 22744 12300
rect 21959 12260 22744 12288
rect 21959 12257 21971 12260
rect 21913 12251 21971 12257
rect 22738 12248 22744 12260
rect 22796 12248 22802 12300
rect 23290 12248 23296 12300
rect 23348 12288 23354 12300
rect 23385 12291 23443 12297
rect 23385 12288 23397 12291
rect 23348 12260 23397 12288
rect 23348 12248 23354 12260
rect 23385 12257 23397 12260
rect 23431 12257 23443 12291
rect 23385 12251 23443 12257
rect 6687 12192 7880 12220
rect 8113 12223 8171 12229
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8846 12220 8852 12232
rect 8159 12192 8852 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12189 10747 12223
rect 14274 12220 14280 12232
rect 14235 12192 14280 12220
rect 10689 12183 10747 12189
rect 5074 12152 5080 12164
rect 4724 12124 5080 12152
rect 5074 12112 5080 12124
rect 5132 12152 5138 12164
rect 7742 12152 7748 12164
rect 5132 12124 7748 12152
rect 5132 12112 5138 12124
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 8202 12112 8208 12164
rect 8260 12152 8266 12164
rect 9309 12155 9367 12161
rect 8260 12124 8708 12152
rect 8260 12112 8266 12124
rect 4798 12084 4804 12096
rect 4759 12056 4804 12084
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 5166 12084 5172 12096
rect 4948 12056 5172 12084
rect 4948 12044 4954 12056
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 5445 12087 5503 12093
rect 5445 12053 5457 12087
rect 5491 12084 5503 12087
rect 5994 12084 6000 12096
rect 5491 12056 6000 12084
rect 5491 12053 5503 12056
rect 5445 12047 5503 12053
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6089 12087 6147 12093
rect 6089 12053 6101 12087
rect 6135 12084 6147 12087
rect 7098 12084 7104 12096
rect 6135 12056 7104 12084
rect 6135 12053 6147 12056
rect 6089 12047 6147 12053
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 8680 12084 8708 12124
rect 9309 12121 9321 12155
rect 9355 12121 9367 12155
rect 9309 12115 9367 12121
rect 9324 12084 9352 12115
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 10704 12152 10732 12183
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15105 12223 15163 12229
rect 15105 12220 15117 12223
rect 14976 12192 15117 12220
rect 14976 12180 14982 12192
rect 15105 12189 15117 12192
rect 15151 12189 15163 12223
rect 15105 12183 15163 12189
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 17276 12192 17785 12220
rect 17276 12180 17282 12192
rect 17773 12189 17785 12192
rect 17819 12220 17831 12223
rect 17862 12220 17868 12232
rect 17819 12192 17868 12220
rect 17819 12189 17831 12192
rect 17773 12183 17831 12189
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 22830 12180 22836 12232
rect 22888 12220 22894 12232
rect 25041 12223 25099 12229
rect 25041 12220 25053 12223
rect 22888 12192 25053 12220
rect 22888 12180 22894 12192
rect 25041 12189 25053 12192
rect 25087 12189 25099 12223
rect 25222 12220 25228 12232
rect 25183 12192 25228 12220
rect 25041 12183 25099 12189
rect 25222 12180 25228 12192
rect 25280 12180 25286 12232
rect 28442 12220 28448 12232
rect 28403 12192 28448 12220
rect 28442 12180 28448 12192
rect 28500 12180 28506 12232
rect 37366 12180 37372 12232
rect 37424 12220 37430 12232
rect 38013 12223 38071 12229
rect 38013 12220 38025 12223
rect 37424 12192 38025 12220
rect 37424 12180 37430 12192
rect 38013 12189 38025 12192
rect 38059 12189 38071 12223
rect 38013 12183 38071 12189
rect 10870 12152 10876 12164
rect 9456 12124 10732 12152
rect 10831 12124 10876 12152
rect 9456 12112 9462 12124
rect 10870 12112 10876 12124
rect 10928 12112 10934 12164
rect 12526 12152 12532 12164
rect 12487 12124 12532 12152
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 13262 12152 13268 12164
rect 13223 12124 13268 12152
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 15010 12112 15016 12164
rect 15068 12152 15074 12164
rect 16025 12155 16083 12161
rect 16025 12152 16037 12155
rect 15068 12124 16037 12152
rect 15068 12112 15074 12124
rect 16025 12121 16037 12124
rect 16071 12121 16083 12155
rect 16025 12115 16083 12121
rect 19334 12112 19340 12164
rect 19392 12152 19398 12164
rect 20165 12155 20223 12161
rect 20165 12152 20177 12155
rect 19392 12124 20177 12152
rect 19392 12112 19398 12124
rect 20165 12121 20177 12124
rect 20211 12121 20223 12155
rect 20165 12115 20223 12121
rect 20254 12112 20260 12164
rect 20312 12152 20318 12164
rect 22005 12155 22063 12161
rect 20312 12124 20357 12152
rect 20312 12112 20318 12124
rect 22005 12121 22017 12155
rect 22051 12152 22063 12155
rect 22094 12152 22100 12164
rect 22051 12124 22100 12152
rect 22051 12121 22063 12124
rect 22005 12115 22063 12121
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 22370 12112 22376 12164
rect 22428 12152 22434 12164
rect 22925 12155 22983 12161
rect 22925 12152 22937 12155
rect 22428 12124 22937 12152
rect 22428 12112 22434 12124
rect 22925 12121 22937 12124
rect 22971 12121 22983 12155
rect 28537 12155 28595 12161
rect 28537 12152 28549 12155
rect 22925 12115 22983 12121
rect 23676 12124 28549 12152
rect 13354 12084 13360 12096
rect 8680 12056 9352 12084
rect 13315 12056 13360 12084
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 14369 12087 14427 12093
rect 14369 12053 14381 12087
rect 14415 12084 14427 12087
rect 14642 12084 14648 12096
rect 14415 12056 14648 12084
rect 14415 12053 14427 12056
rect 14369 12047 14427 12053
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 15197 12087 15255 12093
rect 15197 12053 15209 12087
rect 15243 12084 15255 12087
rect 15286 12084 15292 12096
rect 15243 12056 15292 12084
rect 15243 12053 15255 12056
rect 15197 12047 15255 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 17865 12087 17923 12093
rect 17865 12053 17877 12087
rect 17911 12084 17923 12087
rect 18414 12084 18420 12096
rect 17911 12056 18420 12084
rect 17911 12053 17923 12056
rect 17865 12047 17923 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 19521 12087 19579 12093
rect 19521 12053 19533 12087
rect 19567 12084 19579 12087
rect 19978 12084 19984 12096
rect 19567 12056 19984 12084
rect 19567 12053 19579 12056
rect 19521 12047 19579 12053
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 22738 12044 22744 12096
rect 22796 12084 22802 12096
rect 23676 12084 23704 12124
rect 28537 12121 28549 12124
rect 28583 12121 28595 12155
rect 28537 12115 28595 12121
rect 25682 12084 25688 12096
rect 22796 12056 23704 12084
rect 25643 12056 25688 12084
rect 22796 12044 22802 12056
rect 25682 12044 25688 12056
rect 25740 12044 25746 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 3329 11883 3387 11889
rect 3329 11849 3341 11883
rect 3375 11849 3387 11883
rect 3329 11843 3387 11849
rect 3973 11883 4031 11889
rect 3973 11849 3985 11883
rect 4019 11880 4031 11883
rect 4019 11852 4844 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 3344 11812 3372 11843
rect 4816 11812 4844 11852
rect 5626 11840 5632 11892
rect 5684 11880 5690 11892
rect 7006 11880 7012 11892
rect 5684 11852 7012 11880
rect 5684 11840 5690 11852
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9582 11880 9588 11892
rect 9180 11852 9588 11880
rect 9180 11840 9186 11852
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10226 11880 10232 11892
rect 9815 11852 10232 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 23750 11880 23756 11892
rect 10336 11852 20668 11880
rect 23663 11852 23756 11880
rect 5445 11815 5503 11821
rect 5445 11812 5457 11815
rect 3344 11784 4200 11812
rect 4816 11784 5457 11812
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11744 2099 11747
rect 2590 11744 2596 11756
rect 2087 11716 2596 11744
rect 2087 11713 2099 11716
rect 2041 11707 2099 11713
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11713 2743 11747
rect 3510 11744 3516 11756
rect 3471 11716 3516 11744
rect 2685 11707 2743 11713
rect 2700 11608 2728 11707
rect 3510 11704 3516 11716
rect 3568 11704 3574 11756
rect 4172 11753 4200 11784
rect 5445 11781 5457 11784
rect 5491 11781 5503 11815
rect 5445 11775 5503 11781
rect 6178 11772 6184 11824
rect 6236 11812 6242 11824
rect 8478 11812 8484 11824
rect 6236 11784 8484 11812
rect 6236 11772 6242 11784
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11713 4675 11747
rect 4617 11707 4675 11713
rect 4062 11608 4068 11620
rect 2700 11580 4068 11608
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 4632 11608 4660 11707
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 7208 11753 7236 11784
rect 8478 11772 8484 11784
rect 8536 11772 8542 11824
rect 10336 11812 10364 11852
rect 9324 11784 10364 11812
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 6512 11716 6745 11744
rect 6512 11704 6518 11716
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 8205 11747 8263 11753
rect 8205 11744 8217 11747
rect 7892 11716 8217 11744
rect 7892 11704 7898 11716
rect 8205 11713 8217 11716
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 5166 11636 5172 11688
rect 5224 11676 5230 11688
rect 5353 11679 5411 11685
rect 5353 11676 5365 11679
rect 5224 11648 5365 11676
rect 5224 11636 5230 11648
rect 5353 11645 5365 11648
rect 5399 11645 5411 11679
rect 5626 11676 5632 11688
rect 5587 11648 5632 11676
rect 5353 11639 5411 11645
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 6362 11676 6368 11688
rect 5828 11648 6368 11676
rect 5828 11608 5856 11648
rect 6362 11636 6368 11648
rect 6420 11636 6426 11688
rect 7745 11679 7803 11685
rect 7745 11645 7757 11679
rect 7791 11676 7803 11679
rect 8021 11679 8079 11685
rect 8021 11676 8033 11679
rect 7791 11648 8033 11676
rect 7791 11645 7803 11648
rect 7745 11639 7803 11645
rect 8021 11645 8033 11648
rect 8067 11676 8079 11679
rect 9324 11676 9352 11784
rect 11330 11772 11336 11824
rect 11388 11812 11394 11824
rect 12253 11815 12311 11821
rect 12253 11812 12265 11815
rect 11388 11784 12265 11812
rect 11388 11772 11394 11784
rect 12253 11781 12265 11784
rect 12299 11781 12311 11815
rect 13446 11812 13452 11824
rect 13407 11784 13452 11812
rect 12253 11775 12311 11781
rect 13446 11772 13452 11784
rect 13504 11772 13510 11824
rect 18138 11812 18144 11824
rect 14476 11784 18144 11812
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 8067 11648 9352 11676
rect 9692 11676 9720 11707
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 9824 11716 10333 11744
rect 9824 11704 9830 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 14476 11753 14504 11784
rect 18138 11772 18144 11784
rect 18196 11772 18202 11824
rect 18414 11812 18420 11824
rect 18375 11784 18420 11812
rect 18414 11772 18420 11784
rect 18472 11772 18478 11824
rect 19978 11812 19984 11824
rect 19939 11784 19984 11812
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 20640 11812 20668 11852
rect 23750 11840 23756 11852
rect 23808 11880 23814 11892
rect 24762 11880 24768 11892
rect 23808 11852 24768 11880
rect 23808 11840 23814 11852
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 25041 11883 25099 11889
rect 25041 11849 25053 11883
rect 25087 11880 25099 11883
rect 25222 11880 25228 11892
rect 25087 11852 25228 11880
rect 25087 11849 25099 11852
rect 25041 11843 25099 11849
rect 25222 11840 25228 11852
rect 25280 11840 25286 11892
rect 25682 11840 25688 11892
rect 25740 11880 25746 11892
rect 27801 11883 27859 11889
rect 27801 11880 27813 11883
rect 25740 11852 27813 11880
rect 25740 11840 25746 11852
rect 27801 11849 27813 11852
rect 27847 11849 27859 11883
rect 27801 11843 27859 11849
rect 26234 11812 26240 11824
rect 20640 11784 26240 11812
rect 26234 11772 26240 11784
rect 26292 11772 26298 11824
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10468 11716 10977 11744
rect 10468 11704 10474 11716
rect 10965 11713 10977 11716
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 14461 11747 14519 11753
rect 14461 11713 14473 11747
rect 14507 11713 14519 11747
rect 14642 11744 14648 11756
rect 14603 11716 14648 11744
rect 14461 11707 14519 11713
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 15749 11747 15807 11753
rect 15749 11744 15761 11747
rect 14752 11716 15761 11744
rect 11146 11676 11152 11688
rect 9692 11648 11152 11676
rect 8067 11645 8079 11648
rect 8021 11639 8079 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 12158 11676 12164 11688
rect 12119 11648 12164 11676
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 12250 11636 12256 11688
rect 12308 11676 12314 11688
rect 13357 11679 13415 11685
rect 13357 11676 13369 11679
rect 12308 11648 13369 11676
rect 12308 11636 12314 11648
rect 13357 11645 13369 11648
rect 13403 11645 13415 11679
rect 13357 11639 13415 11645
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14752 11676 14780 11716
rect 15749 11713 15761 11716
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 21726 11704 21732 11756
rect 21784 11744 21790 11756
rect 22465 11747 22523 11753
rect 22465 11744 22477 11747
rect 21784 11716 22477 11744
rect 21784 11704 21790 11716
rect 22465 11713 22477 11716
rect 22511 11713 22523 11747
rect 22465 11707 22523 11713
rect 22557 11747 22615 11753
rect 22557 11713 22569 11747
rect 22603 11744 22615 11747
rect 23293 11747 23351 11753
rect 23293 11744 23305 11747
rect 22603 11716 23305 11744
rect 22603 11713 22615 11716
rect 22557 11707 22615 11713
rect 23293 11713 23305 11716
rect 23339 11713 23351 11747
rect 23293 11707 23351 11713
rect 23566 11704 23572 11756
rect 23624 11744 23630 11756
rect 24949 11747 25007 11753
rect 23624 11716 24900 11744
rect 23624 11704 23630 11716
rect 14332 11648 14780 11676
rect 15105 11679 15163 11685
rect 14332 11636 14338 11648
rect 15105 11645 15117 11679
rect 15151 11676 15163 11679
rect 15378 11676 15384 11688
rect 15151 11648 15384 11676
rect 15151 11645 15163 11648
rect 15105 11639 15163 11645
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 18322 11676 18328 11688
rect 18283 11648 18328 11676
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 18966 11676 18972 11688
rect 18927 11648 18972 11676
rect 18966 11636 18972 11648
rect 19024 11636 19030 11688
rect 19889 11679 19947 11685
rect 19889 11645 19901 11679
rect 19935 11676 19947 11679
rect 20162 11676 20168 11688
rect 19935 11648 20168 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 20533 11679 20591 11685
rect 20533 11645 20545 11679
rect 20579 11676 20591 11679
rect 20579 11648 20668 11676
rect 20579 11645 20591 11648
rect 20533 11639 20591 11645
rect 20640 11620 20668 11648
rect 21266 11636 21272 11688
rect 21324 11676 21330 11688
rect 23014 11676 23020 11688
rect 21324 11648 23020 11676
rect 21324 11636 21330 11648
rect 23014 11636 23020 11648
rect 23072 11676 23078 11688
rect 23109 11679 23167 11685
rect 23109 11676 23121 11679
rect 23072 11648 23121 11676
rect 23072 11636 23078 11648
rect 23109 11645 23121 11648
rect 23155 11645 23167 11679
rect 23109 11639 23167 11645
rect 24305 11679 24363 11685
rect 24305 11645 24317 11679
rect 24351 11676 24363 11679
rect 24670 11676 24676 11688
rect 24351 11648 24676 11676
rect 24351 11645 24363 11648
rect 24305 11639 24363 11645
rect 7282 11608 7288 11620
rect 4632 11580 5856 11608
rect 7195 11580 7288 11608
rect 7282 11568 7288 11580
rect 7340 11608 7346 11620
rect 9398 11608 9404 11620
rect 7340 11580 9404 11608
rect 7340 11568 7346 11580
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 10413 11611 10471 11617
rect 10413 11577 10425 11611
rect 10459 11608 10471 11611
rect 11882 11608 11888 11620
rect 10459 11580 11888 11608
rect 10459 11577 10471 11580
rect 10413 11571 10471 11577
rect 11882 11568 11888 11580
rect 11940 11568 11946 11620
rect 12713 11611 12771 11617
rect 12713 11577 12725 11611
rect 12759 11608 12771 11611
rect 13909 11611 13967 11617
rect 13909 11608 13921 11611
rect 12759 11580 13921 11608
rect 12759 11577 12771 11580
rect 12713 11571 12771 11577
rect 13909 11577 13921 11580
rect 13955 11608 13967 11611
rect 13955 11580 16574 11608
rect 13955 11577 13967 11580
rect 13909 11571 13967 11577
rect 2130 11540 2136 11552
rect 2091 11512 2136 11540
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 2222 11500 2228 11552
rect 2280 11540 2286 11552
rect 2777 11543 2835 11549
rect 2777 11540 2789 11543
rect 2280 11512 2789 11540
rect 2280 11500 2286 11512
rect 2777 11509 2789 11512
rect 2823 11509 2835 11543
rect 2777 11503 2835 11509
rect 4709 11543 4767 11549
rect 4709 11509 4721 11543
rect 4755 11540 4767 11543
rect 5442 11540 5448 11552
rect 4755 11512 5448 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 7190 11540 7196 11552
rect 6871 11512 7196 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 8352 11512 8401 11540
rect 8352 11500 8358 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 10962 11540 10968 11552
rect 8536 11512 10968 11540
rect 8536 11500 8542 11512
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 11146 11540 11152 11552
rect 11103 11512 11152 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15565 11543 15623 11549
rect 15565 11540 15577 11543
rect 15252 11512 15577 11540
rect 15252 11500 15258 11512
rect 15565 11509 15577 11512
rect 15611 11509 15623 11543
rect 16546 11540 16574 11580
rect 20622 11568 20628 11620
rect 20680 11568 20686 11620
rect 22830 11540 22836 11552
rect 16546 11512 22836 11540
rect 15565 11503 15623 11509
rect 22830 11500 22836 11512
rect 22888 11500 22894 11552
rect 23124 11540 23152 11639
rect 24670 11636 24676 11648
rect 24728 11636 24734 11688
rect 24872 11676 24900 11716
rect 24949 11713 24961 11747
rect 24995 11744 25007 11747
rect 25130 11744 25136 11756
rect 24995 11716 25136 11744
rect 24995 11713 25007 11716
rect 24949 11707 25007 11713
rect 25130 11704 25136 11716
rect 25188 11744 25194 11756
rect 25777 11747 25835 11753
rect 25777 11744 25789 11747
rect 25188 11716 25789 11744
rect 25188 11704 25194 11716
rect 25777 11713 25789 11716
rect 25823 11713 25835 11747
rect 25777 11707 25835 11713
rect 25866 11704 25872 11756
rect 25924 11744 25930 11756
rect 27706 11744 27712 11756
rect 25924 11716 27712 11744
rect 25924 11704 25930 11716
rect 27706 11704 27712 11716
rect 27764 11704 27770 11756
rect 27816 11744 27844 11843
rect 28261 11747 28319 11753
rect 28261 11744 28273 11747
rect 27816 11716 28273 11744
rect 28261 11713 28273 11716
rect 28307 11713 28319 11747
rect 28261 11707 28319 11713
rect 24872 11648 26004 11676
rect 23198 11568 23204 11620
rect 23256 11608 23262 11620
rect 25866 11608 25872 11620
rect 23256 11580 25872 11608
rect 23256 11568 23262 11580
rect 25866 11568 25872 11580
rect 25924 11568 25930 11620
rect 25976 11608 26004 11648
rect 26050 11636 26056 11688
rect 26108 11676 26114 11688
rect 26326 11676 26332 11688
rect 26108 11648 26332 11676
rect 26108 11636 26114 11648
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 26970 11636 26976 11688
rect 27028 11676 27034 11688
rect 27157 11679 27215 11685
rect 27157 11676 27169 11679
rect 27028 11648 27169 11676
rect 27028 11636 27034 11648
rect 27157 11645 27169 11648
rect 27203 11645 27215 11679
rect 27338 11676 27344 11688
rect 27299 11648 27344 11676
rect 27157 11639 27215 11645
rect 27338 11636 27344 11648
rect 27396 11636 27402 11688
rect 31846 11608 31852 11620
rect 25976 11580 31852 11608
rect 31846 11568 31852 11580
rect 31904 11568 31910 11620
rect 24946 11540 24952 11552
rect 23124 11512 24952 11540
rect 24946 11500 24952 11512
rect 25004 11500 25010 11552
rect 25593 11543 25651 11549
rect 25593 11509 25605 11543
rect 25639 11540 25651 11543
rect 26510 11540 26516 11552
rect 25639 11512 26516 11540
rect 25639 11509 25651 11512
rect 25593 11503 25651 11509
rect 26510 11500 26516 11512
rect 26568 11500 26574 11552
rect 28353 11543 28411 11549
rect 28353 11509 28365 11543
rect 28399 11540 28411 11543
rect 34422 11540 34428 11552
rect 28399 11512 34428 11540
rect 28399 11509 28411 11512
rect 28353 11503 28411 11509
rect 34422 11500 34428 11512
rect 34480 11500 34486 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1578 11296 1584 11348
rect 1636 11336 1642 11348
rect 1765 11339 1823 11345
rect 1765 11336 1777 11339
rect 1636 11308 1777 11336
rect 1636 11296 1642 11308
rect 1765 11305 1777 11308
rect 1811 11305 1823 11339
rect 1765 11299 1823 11305
rect 2038 11296 2044 11348
rect 2096 11336 2102 11348
rect 3973 11339 4031 11345
rect 3973 11336 3985 11339
rect 2096 11308 3985 11336
rect 2096 11296 2102 11308
rect 3973 11305 3985 11308
rect 4019 11305 4031 11339
rect 3973 11299 4031 11305
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 5626 11336 5632 11348
rect 4120 11308 5632 11336
rect 4120 11296 4126 11308
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 6604 11308 9689 11336
rect 6604 11296 6610 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 9677 11299 9735 11305
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11974 11336 11980 11348
rect 11112 11308 11980 11336
rect 11112 11296 11118 11308
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 12584 11308 23980 11336
rect 12584 11296 12590 11308
rect 3329 11271 3387 11277
rect 3329 11237 3341 11271
rect 3375 11268 3387 11271
rect 4982 11268 4988 11280
rect 3375 11240 4988 11268
rect 3375 11237 3387 11240
rect 3329 11231 3387 11237
rect 4982 11228 4988 11240
rect 5040 11228 5046 11280
rect 6825 11271 6883 11277
rect 6825 11237 6837 11271
rect 6871 11268 6883 11271
rect 7834 11268 7840 11280
rect 6871 11240 7840 11268
rect 6871 11237 6883 11240
rect 6825 11231 6883 11237
rect 7834 11228 7840 11240
rect 7892 11228 7898 11280
rect 10042 11268 10048 11280
rect 8496 11240 10048 11268
rect 4706 11200 4712 11212
rect 4172 11172 4712 11200
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11132 2007 11135
rect 2222 11132 2228 11144
rect 1995 11104 2228 11132
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11132 2467 11135
rect 2682 11132 2688 11144
rect 2455 11104 2688 11132
rect 2455 11101 2467 11104
rect 2409 11095 2467 11101
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 4062 11132 4068 11144
rect 3283 11104 4068 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4172 11141 4200 11172
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5350 11200 5356 11212
rect 4816 11172 5356 11200
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4304 11104 4629 11132
rect 4304 11092 4310 11104
rect 4617 11101 4629 11104
rect 4663 11132 4675 11135
rect 4816 11132 4844 11172
rect 5350 11160 5356 11172
rect 5408 11160 5414 11212
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5629 11203 5687 11209
rect 5629 11200 5641 11203
rect 5592 11172 5641 11200
rect 5592 11160 5598 11172
rect 5629 11169 5641 11172
rect 5675 11200 5687 11203
rect 8496 11200 8524 11240
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 14734 11228 14740 11280
rect 14792 11268 14798 11280
rect 15654 11268 15660 11280
rect 14792 11240 15660 11268
rect 14792 11228 14798 11240
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 23198 11268 23204 11280
rect 16546 11240 23204 11268
rect 5675 11172 8524 11200
rect 8573 11203 8631 11209
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 8573 11169 8585 11203
rect 8619 11200 8631 11203
rect 9490 11200 9496 11212
rect 8619 11172 9496 11200
rect 8619 11169 8631 11172
rect 8573 11163 8631 11169
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 11330 11200 11336 11212
rect 11291 11172 11336 11200
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 16546 11200 16574 11240
rect 23198 11228 23204 11240
rect 23256 11228 23262 11280
rect 13679 11172 16574 11200
rect 19521 11203 19579 11209
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 19521 11169 19533 11203
rect 19567 11200 19579 11203
rect 19978 11200 19984 11212
rect 19567 11172 19984 11200
rect 19567 11169 19579 11172
rect 19521 11163 19579 11169
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 20346 11200 20352 11212
rect 20307 11172 20352 11200
rect 20346 11160 20352 11172
rect 20404 11160 20410 11212
rect 22649 11203 22707 11209
rect 22649 11169 22661 11203
rect 22695 11200 22707 11203
rect 23385 11203 23443 11209
rect 23385 11200 23397 11203
rect 22695 11172 23397 11200
rect 22695 11169 22707 11172
rect 22649 11163 22707 11169
rect 23385 11169 23397 11172
rect 23431 11169 23443 11203
rect 23385 11163 23443 11169
rect 4663 11104 4844 11132
rect 7009 11135 7067 11141
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7374 11132 7380 11144
rect 7055 11104 7380 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 9122 11132 9128 11144
rect 9083 11104 9128 11132
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9306 11132 9312 11144
rect 9267 11104 9312 11132
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 9640 11104 10333 11132
rect 9640 11092 9646 11104
rect 10321 11101 10333 11104
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 15013 11135 15071 11141
rect 15013 11101 15025 11135
rect 15059 11132 15071 11135
rect 15194 11132 15200 11144
rect 15059 11104 15200 11132
rect 15059 11101 15071 11104
rect 15013 11095 15071 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 20990 11092 20996 11144
rect 21048 11132 21054 11144
rect 21085 11135 21143 11141
rect 21085 11132 21097 11135
rect 21048 11104 21097 11132
rect 21048 11092 21054 11104
rect 21085 11101 21097 11104
rect 21131 11132 21143 11135
rect 21726 11132 21732 11144
rect 21131 11104 21732 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 21726 11092 21732 11104
rect 21784 11092 21790 11144
rect 22462 11092 22468 11144
rect 22520 11132 22526 11144
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 22520 11104 22569 11132
rect 22520 11092 22526 11104
rect 22557 11101 22569 11104
rect 22603 11101 22615 11135
rect 22557 11095 22615 11101
rect 23201 11135 23259 11141
rect 23201 11101 23213 11135
rect 23247 11132 23259 11135
rect 23750 11132 23756 11144
rect 23247 11104 23756 11132
rect 23247 11101 23259 11104
rect 23201 11095 23259 11101
rect 23750 11092 23756 11104
rect 23808 11092 23814 11144
rect 5350 11064 5356 11076
rect 5311 11036 5356 11064
rect 5350 11024 5356 11036
rect 5408 11024 5414 11076
rect 5442 11024 5448 11076
rect 5500 11064 5506 11076
rect 5500 11036 5545 11064
rect 5500 11024 5506 11036
rect 6454 11024 6460 11076
rect 6512 11064 6518 11076
rect 7561 11067 7619 11073
rect 7561 11064 7573 11067
rect 6512 11036 7573 11064
rect 6512 11024 6518 11036
rect 7561 11033 7573 11036
rect 7607 11033 7619 11067
rect 7561 11027 7619 11033
rect 7653 11067 7711 11073
rect 7653 11033 7665 11067
rect 7699 11064 7711 11067
rect 8202 11064 8208 11076
rect 7699 11036 8208 11064
rect 7699 11033 7711 11036
rect 7653 11027 7711 11033
rect 8202 11024 8208 11036
rect 8260 11024 8266 11076
rect 10410 11064 10416 11076
rect 10371 11036 10416 11064
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 11054 11064 11060 11076
rect 11015 11036 11060 11064
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11204 11036 11249 11064
rect 11204 11024 11210 11036
rect 11698 11024 11704 11076
rect 11756 11064 11762 11076
rect 12158 11064 12164 11076
rect 11756 11036 12164 11064
rect 11756 11024 11762 11036
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 12618 11064 12624 11076
rect 12579 11036 12624 11064
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 12710 11024 12716 11076
rect 12768 11064 12774 11076
rect 15562 11064 15568 11076
rect 12768 11036 12813 11064
rect 15523 11036 15568 11064
rect 12768 11024 12774 11036
rect 15562 11024 15568 11036
rect 15620 11024 15626 11076
rect 15654 11024 15660 11076
rect 15712 11064 15718 11076
rect 16206 11064 16212 11076
rect 15712 11036 15757 11064
rect 16167 11036 16212 11064
rect 15712 11024 15718 11036
rect 16206 11024 16212 11036
rect 16264 11024 16270 11076
rect 19613 11067 19671 11073
rect 19613 11033 19625 11067
rect 19659 11064 19671 11067
rect 20070 11064 20076 11076
rect 19659 11036 20076 11064
rect 19659 11033 19671 11036
rect 19613 11027 19671 11033
rect 20070 11024 20076 11036
rect 20128 11024 20134 11076
rect 23842 11064 23848 11076
rect 23803 11036 23848 11064
rect 23842 11024 23848 11036
rect 23900 11024 23906 11076
rect 23952 11064 23980 11308
rect 24946 11296 24952 11348
rect 25004 11336 25010 11348
rect 26050 11336 26056 11348
rect 25004 11308 26056 11336
rect 25004 11296 25010 11308
rect 26050 11296 26056 11308
rect 26108 11296 26114 11348
rect 26329 11339 26387 11345
rect 26329 11305 26341 11339
rect 26375 11336 26387 11339
rect 27338 11336 27344 11348
rect 26375 11308 27344 11336
rect 26375 11305 26387 11308
rect 26329 11299 26387 11305
rect 27338 11296 27344 11308
rect 27396 11296 27402 11348
rect 24210 11228 24216 11280
rect 24268 11268 24274 11280
rect 28077 11271 28135 11277
rect 28077 11268 28089 11271
rect 24268 11240 28089 11268
rect 24268 11228 24274 11240
rect 28077 11237 28089 11240
rect 28123 11237 28135 11271
rect 28077 11231 28135 11237
rect 37458 11228 37464 11280
rect 37516 11228 37522 11280
rect 24670 11200 24676 11212
rect 24631 11172 24676 11200
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 26970 11200 26976 11212
rect 26931 11172 26976 11200
rect 26970 11160 26976 11172
rect 27028 11160 27034 11212
rect 37476 11200 37504 11228
rect 37737 11203 37795 11209
rect 37737 11200 37749 11203
rect 37476 11172 37749 11200
rect 37737 11169 37749 11172
rect 37783 11169 37795 11203
rect 37737 11163 37795 11169
rect 26510 11132 26516 11144
rect 26471 11104 26516 11132
rect 26510 11092 26516 11104
rect 26568 11092 26574 11144
rect 27982 11132 27988 11144
rect 27943 11104 27988 11132
rect 27982 11092 27988 11104
rect 28040 11092 28046 11144
rect 31846 11132 31852 11144
rect 31807 11104 31852 11132
rect 31846 11092 31852 11104
rect 31904 11092 31910 11144
rect 37182 11092 37188 11144
rect 37240 11132 37246 11144
rect 37461 11135 37519 11141
rect 37461 11132 37473 11135
rect 37240 11104 37473 11132
rect 37240 11092 37246 11104
rect 37461 11101 37473 11104
rect 37507 11101 37519 11135
rect 37461 11095 37519 11101
rect 24765 11067 24823 11073
rect 23952 11036 24716 11064
rect 2314 10956 2320 11008
rect 2372 10996 2378 11008
rect 2501 10999 2559 11005
rect 2501 10996 2513 10999
rect 2372 10968 2513 10996
rect 2372 10956 2378 10968
rect 2501 10965 2513 10968
rect 2547 10965 2559 10999
rect 2501 10959 2559 10965
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 4709 10999 4767 11005
rect 4709 10996 4721 10999
rect 3292 10968 4721 10996
rect 3292 10956 3298 10968
rect 4709 10965 4721 10968
rect 4755 10965 4767 10999
rect 4709 10959 4767 10965
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 9674 10996 9680 11008
rect 7248 10968 9680 10996
rect 7248 10956 7254 10968
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 14366 10996 14372 11008
rect 10836 10968 14372 10996
rect 10836 10956 10842 10968
rect 14366 10956 14372 10968
rect 14424 10956 14430 11008
rect 14826 10996 14832 11008
rect 14787 10968 14832 10996
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 14918 10956 14924 11008
rect 14976 10996 14982 11008
rect 17218 10996 17224 11008
rect 14976 10968 17224 10996
rect 14976 10956 14982 10968
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 17310 10956 17316 11008
rect 17368 10996 17374 11008
rect 19426 10996 19432 11008
rect 17368 10968 19432 10996
rect 17368 10956 17374 10968
rect 19426 10956 19432 10968
rect 19484 10956 19490 11008
rect 21174 10996 21180 11008
rect 21135 10968 21180 10996
rect 21174 10956 21180 10968
rect 21232 10956 21238 11008
rect 24688 10996 24716 11036
rect 24765 11033 24777 11067
rect 24811 11064 24823 11067
rect 25038 11064 25044 11076
rect 24811 11036 25044 11064
rect 24811 11033 24823 11036
rect 24765 11027 24823 11033
rect 25038 11024 25044 11036
rect 25096 11024 25102 11076
rect 25314 11064 25320 11076
rect 25275 11036 25320 11064
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 28074 11064 28080 11076
rect 25424 11036 28080 11064
rect 25424 10996 25452 11036
rect 28074 11024 28080 11036
rect 28132 11064 28138 11076
rect 31941 11067 31999 11073
rect 28132 11036 29316 11064
rect 28132 11024 28138 11036
rect 24688 10968 25452 10996
rect 29288 10996 29316 11036
rect 31941 11033 31953 11067
rect 31987 11064 31999 11067
rect 32582 11064 32588 11076
rect 31987 11036 32588 11064
rect 31987 11033 31999 11036
rect 31941 11027 31999 11033
rect 32582 11024 32588 11036
rect 32640 11024 32646 11076
rect 33134 10996 33140 11008
rect 29288 10968 33140 10996
rect 33134 10956 33140 10968
rect 33192 10956 33198 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 3418 10792 3424 10804
rect 1780 10764 3424 10792
rect 1780 10665 1808 10764
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 5350 10792 5356 10804
rect 5311 10764 5356 10792
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 7653 10795 7711 10801
rect 7653 10761 7665 10795
rect 7699 10792 7711 10795
rect 9306 10792 9312 10804
rect 7699 10764 9312 10792
rect 7699 10761 7711 10764
rect 7653 10755 7711 10761
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 9600 10764 10272 10792
rect 2590 10724 2596 10736
rect 2551 10696 2596 10724
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 3510 10724 3516 10736
rect 3423 10696 3516 10724
rect 3510 10684 3516 10696
rect 3568 10724 3574 10736
rect 7006 10724 7012 10736
rect 3568 10696 7012 10724
rect 3568 10684 3574 10696
rect 7006 10684 7012 10696
rect 7064 10684 7070 10736
rect 7098 10684 7104 10736
rect 7156 10724 7162 10736
rect 8481 10727 8539 10733
rect 8481 10724 8493 10727
rect 7156 10696 8493 10724
rect 7156 10684 7162 10696
rect 8481 10693 8493 10696
rect 8527 10693 8539 10727
rect 8481 10687 8539 10693
rect 9033 10727 9091 10733
rect 9033 10693 9045 10727
rect 9079 10724 9091 10727
rect 9600 10724 9628 10764
rect 9079 10696 9628 10724
rect 9079 10693 9091 10696
rect 9033 10687 9091 10693
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 10244 10733 10272 10764
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10928 10764 10977 10792
rect 10928 10752 10934 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 11072 10764 12480 10792
rect 10229 10727 10287 10733
rect 9732 10696 9777 10724
rect 9732 10684 9738 10696
rect 10229 10693 10241 10727
rect 10275 10724 10287 10727
rect 11072 10724 11100 10764
rect 11882 10724 11888 10736
rect 10275 10696 11100 10724
rect 11843 10696 11888 10724
rect 10275 10693 10287 10696
rect 10229 10687 10287 10693
rect 11882 10684 11888 10696
rect 11940 10684 11946 10736
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4798 10656 4804 10668
rect 4295 10628 4804 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 6052 10628 6745 10656
rect 6052 10616 6058 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 7834 10656 7840 10668
rect 7795 10628 7840 10656
rect 6733 10619 6791 10625
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10656 10931 10659
rect 11238 10656 11244 10668
rect 10919 10628 11244 10656
rect 10919 10625 10931 10628
rect 10873 10619 10931 10625
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10557 2559 10591
rect 2501 10551 2559 10557
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10557 4123 10591
rect 4065 10551 4123 10557
rect 6549 10591 6607 10597
rect 6549 10557 6561 10591
rect 6595 10588 6607 10591
rect 7282 10588 7288 10600
rect 6595 10560 7288 10588
rect 6595 10557 6607 10560
rect 6549 10551 6607 10557
rect 2406 10480 2412 10532
rect 2464 10520 2470 10532
rect 2516 10520 2544 10551
rect 2464 10492 2544 10520
rect 4080 10520 4108 10551
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8478 10588 8484 10600
rect 8435 10560 8484 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8478 10548 8484 10560
rect 8536 10548 8542 10600
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10588 9643 10591
rect 11790 10588 11796 10600
rect 9631 10560 11468 10588
rect 11751 10560 11796 10588
rect 9631 10557 9643 10560
rect 9585 10551 9643 10557
rect 8294 10520 8300 10532
rect 4080 10492 8300 10520
rect 2464 10480 2470 10492
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 11440 10520 11468 10560
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10557 12127 10591
rect 12452 10588 12480 10764
rect 13446 10752 13452 10804
rect 13504 10792 13510 10804
rect 13541 10795 13599 10801
rect 13541 10792 13553 10795
rect 13504 10764 13553 10792
rect 13504 10752 13510 10764
rect 13541 10761 13553 10764
rect 13587 10761 13599 10795
rect 13541 10755 13599 10761
rect 14185 10795 14243 10801
rect 14185 10761 14197 10795
rect 14231 10761 14243 10795
rect 14185 10755 14243 10761
rect 14090 10724 14096 10736
rect 12912 10696 14096 10724
rect 12912 10668 12940 10696
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 12894 10656 12900 10668
rect 12855 10628 12900 10656
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 14200 10656 14228 10755
rect 17218 10752 17224 10804
rect 17276 10792 17282 10804
rect 17276 10764 18276 10792
rect 17276 10752 17282 10764
rect 17954 10724 17960 10736
rect 17915 10696 17960 10724
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18248 10724 18276 10764
rect 18322 10752 18328 10804
rect 18380 10792 18386 10804
rect 19061 10795 19119 10801
rect 19061 10792 19073 10795
rect 18380 10764 19073 10792
rect 18380 10752 18386 10764
rect 19061 10761 19073 10764
rect 19107 10761 19119 10795
rect 19061 10755 19119 10761
rect 19889 10795 19947 10801
rect 19889 10761 19901 10795
rect 19935 10792 19947 10795
rect 20254 10792 20260 10804
rect 19935 10764 20260 10792
rect 19935 10761 19947 10764
rect 19889 10755 19947 10761
rect 20254 10752 20260 10764
rect 20312 10752 20318 10804
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 23845 10795 23903 10801
rect 23845 10792 23857 10795
rect 23532 10764 23857 10792
rect 23532 10752 23538 10764
rect 23845 10761 23857 10764
rect 23891 10761 23903 10795
rect 23845 10755 23903 10761
rect 25314 10724 25320 10736
rect 18248 10696 25320 10724
rect 25314 10684 25320 10696
rect 25372 10684 25378 10736
rect 14366 10656 14372 10668
rect 13771 10628 14228 10656
rect 14327 10628 14372 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14884 10628 15117 10656
rect 14884 10616 14890 10628
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10656 17187 10659
rect 17310 10656 17316 10668
rect 17175 10628 17316 10656
rect 17175 10625 17187 10628
rect 17129 10619 17187 10625
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 18969 10659 19027 10665
rect 18969 10625 18981 10659
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10656 19855 10659
rect 20898 10656 20904 10668
rect 19843 10628 20904 10656
rect 19843 10625 19855 10628
rect 19797 10619 19855 10625
rect 14550 10588 14556 10600
rect 12452 10560 14556 10588
rect 12069 10551 12127 10557
rect 12084 10520 12112 10551
rect 14550 10548 14556 10560
rect 14608 10548 14614 10600
rect 14918 10588 14924 10600
rect 14879 10560 14924 10588
rect 14918 10548 14924 10560
rect 14976 10548 14982 10600
rect 17862 10588 17868 10600
rect 17823 10560 17868 10588
rect 17862 10548 17868 10560
rect 17920 10548 17926 10600
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 16206 10520 16212 10532
rect 11440 10492 16212 10520
rect 16206 10480 16212 10492
rect 16264 10520 16270 10532
rect 16264 10492 17540 10520
rect 16264 10480 16270 10492
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 1857 10455 1915 10461
rect 1857 10452 1869 10455
rect 1820 10424 1869 10452
rect 1820 10412 1826 10424
rect 1857 10421 1869 10424
rect 1903 10421 1915 10455
rect 1857 10415 1915 10421
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 4433 10455 4491 10461
rect 4433 10452 4445 10455
rect 3568 10424 4445 10452
rect 3568 10412 3574 10424
rect 4433 10421 4445 10424
rect 4479 10421 4491 10455
rect 4433 10415 4491 10421
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 6917 10455 6975 10461
rect 6917 10452 6929 10455
rect 5224 10424 6929 10452
rect 5224 10412 5230 10424
rect 6917 10421 6929 10424
rect 6963 10421 6975 10455
rect 6917 10415 6975 10421
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 11330 10452 11336 10464
rect 7064 10424 11336 10452
rect 7064 10412 7070 10424
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12989 10455 13047 10461
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 14734 10452 14740 10464
rect 13035 10424 14740 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 15289 10455 15347 10461
rect 15289 10452 15301 10455
rect 15252 10424 15301 10452
rect 15252 10412 15258 10424
rect 15289 10421 15301 10424
rect 15335 10452 15347 10455
rect 15378 10452 15384 10464
rect 15335 10424 15384 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 17221 10455 17279 10461
rect 17221 10421 17233 10455
rect 17267 10452 17279 10455
rect 17402 10452 17408 10464
rect 17267 10424 17408 10452
rect 17267 10421 17279 10424
rect 17221 10415 17279 10421
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 17512 10452 17540 10492
rect 18156 10452 18184 10551
rect 18230 10548 18236 10600
rect 18288 10588 18294 10600
rect 18984 10588 19012 10619
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 20993 10659 21051 10665
rect 20993 10625 21005 10659
rect 21039 10656 21051 10659
rect 21174 10656 21180 10668
rect 21039 10628 21180 10656
rect 21039 10625 21051 10628
rect 20993 10619 21051 10625
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 22462 10616 22468 10668
rect 22520 10656 22526 10668
rect 23293 10659 23351 10665
rect 23293 10656 23305 10659
rect 22520 10628 23305 10656
rect 22520 10616 22526 10628
rect 23293 10625 23305 10628
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 23753 10659 23811 10665
rect 23753 10625 23765 10659
rect 23799 10656 23811 10659
rect 24670 10656 24676 10668
rect 23799 10628 24676 10656
rect 23799 10625 23811 10628
rect 23753 10619 23811 10625
rect 24670 10616 24676 10628
rect 24728 10616 24734 10668
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 25041 10659 25099 10665
rect 25041 10656 25053 10659
rect 24912 10628 25053 10656
rect 24912 10616 24918 10628
rect 25041 10625 25053 10628
rect 25087 10625 25099 10659
rect 25041 10619 25099 10625
rect 18288 10560 19012 10588
rect 18288 10548 18294 10560
rect 20162 10548 20168 10600
rect 20220 10588 20226 10600
rect 20622 10588 20628 10600
rect 20220 10560 20628 10588
rect 20220 10548 20226 10560
rect 20622 10548 20628 10560
rect 20680 10588 20686 10600
rect 20809 10591 20867 10597
rect 20809 10588 20821 10591
rect 20680 10560 20821 10588
rect 20680 10548 20686 10560
rect 20809 10557 20821 10560
rect 20855 10557 20867 10591
rect 22005 10591 22063 10597
rect 22005 10588 22017 10591
rect 20809 10551 20867 10557
rect 21192 10560 22017 10588
rect 21192 10464 21220 10560
rect 22005 10557 22017 10560
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 22189 10591 22247 10597
rect 22189 10557 22201 10591
rect 22235 10588 22247 10591
rect 22278 10588 22284 10600
rect 22235 10560 22284 10588
rect 22235 10557 22247 10560
rect 22189 10551 22247 10557
rect 22278 10548 22284 10560
rect 22336 10548 22342 10600
rect 22649 10591 22707 10597
rect 22649 10557 22661 10591
rect 22695 10588 22707 10591
rect 23842 10588 23848 10600
rect 22695 10560 23848 10588
rect 22695 10557 22707 10560
rect 22649 10551 22707 10557
rect 23842 10548 23848 10560
rect 23900 10548 23906 10600
rect 21174 10452 21180 10464
rect 17512 10424 18184 10452
rect 21135 10424 21180 10452
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 23106 10452 23112 10464
rect 23067 10424 23112 10452
rect 23106 10412 23112 10424
rect 23164 10412 23170 10464
rect 24854 10452 24860 10464
rect 24815 10424 24860 10452
rect 24854 10412 24860 10424
rect 24912 10412 24918 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 8846 10208 8852 10260
rect 8904 10248 8910 10260
rect 9585 10251 9643 10257
rect 9585 10248 9597 10251
rect 8904 10220 9597 10248
rect 8904 10208 8910 10220
rect 9585 10217 9597 10220
rect 9631 10217 9643 10251
rect 9585 10211 9643 10217
rect 12618 10208 12624 10260
rect 12676 10248 12682 10260
rect 13357 10251 13415 10257
rect 13357 10248 13369 10251
rect 12676 10220 13369 10248
rect 12676 10208 12682 10220
rect 13357 10217 13369 10220
rect 13403 10217 13415 10251
rect 13357 10211 13415 10217
rect 17862 10208 17868 10260
rect 17920 10248 17926 10260
rect 19889 10251 19947 10257
rect 17920 10220 19840 10248
rect 17920 10208 17926 10220
rect 2869 10183 2927 10189
rect 2869 10149 2881 10183
rect 2915 10180 2927 10183
rect 8478 10180 8484 10192
rect 2915 10152 8484 10180
rect 2915 10149 2927 10152
rect 2869 10143 2927 10149
rect 8478 10140 8484 10152
rect 8536 10140 8542 10192
rect 12437 10183 12495 10189
rect 12437 10149 12449 10183
rect 12483 10180 12495 10183
rect 17954 10180 17960 10192
rect 12483 10152 17960 10180
rect 12483 10149 12495 10152
rect 12437 10143 12495 10149
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 19334 10180 19340 10192
rect 18248 10152 19340 10180
rect 2314 10112 2320 10124
rect 2275 10084 2320 10112
rect 2314 10072 2320 10084
rect 2372 10072 2378 10124
rect 2958 10072 2964 10124
rect 3016 10112 3022 10124
rect 3418 10112 3424 10124
rect 3016 10084 3424 10112
rect 3016 10072 3022 10084
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 4890 10072 4896 10124
rect 4948 10112 4954 10124
rect 7653 10115 7711 10121
rect 4948 10084 7604 10112
rect 4948 10072 4954 10084
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 5169 10047 5227 10053
rect 5169 10044 5181 10047
rect 5132 10016 5181 10044
rect 5132 10004 5138 10016
rect 5169 10013 5181 10016
rect 5215 10013 5227 10047
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 5169 10007 5227 10013
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7576 10044 7604 10084
rect 7653 10081 7665 10115
rect 7699 10112 7711 10115
rect 9122 10112 9128 10124
rect 7699 10084 9128 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 18248 10112 18276 10152
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 19812 10180 19840 10220
rect 19889 10217 19901 10251
rect 19935 10248 19947 10251
rect 19978 10248 19984 10260
rect 19935 10220 19984 10248
rect 19935 10217 19947 10220
rect 19889 10211 19947 10217
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 22278 10248 22284 10260
rect 22239 10220 22284 10248
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 25038 10208 25044 10260
rect 25096 10248 25102 10260
rect 25225 10251 25283 10257
rect 25225 10248 25237 10251
rect 25096 10220 25237 10248
rect 25096 10208 25102 10220
rect 25225 10217 25237 10220
rect 25271 10217 25283 10251
rect 25225 10211 25283 10217
rect 23014 10180 23020 10192
rect 19812 10152 23020 10180
rect 23014 10140 23020 10152
rect 23072 10140 23078 10192
rect 9692 10084 12388 10112
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 7576 10016 8401 10044
rect 8389 10013 8401 10016
rect 8435 10044 8447 10047
rect 9692 10044 9720 10084
rect 8435 10016 9720 10044
rect 9769 10047 9827 10053
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 9769 10013 9781 10047
rect 9815 10044 9827 10047
rect 9858 10044 9864 10056
rect 9815 10016 9864 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10044 11115 10047
rect 11146 10044 11152 10056
rect 11103 10016 11152 10044
rect 11103 10013 11115 10016
rect 11057 10007 11115 10013
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 12360 10053 12388 10084
rect 12452 10084 18276 10112
rect 18325 10115 18383 10121
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 2130 9936 2136 9988
rect 2188 9976 2194 9988
rect 2409 9979 2467 9985
rect 2409 9976 2421 9979
rect 2188 9948 2421 9976
rect 2188 9936 2194 9948
rect 2409 9945 2421 9948
rect 2455 9945 2467 9979
rect 2409 9939 2467 9945
rect 6917 9979 6975 9985
rect 6917 9945 6929 9979
rect 6963 9976 6975 9979
rect 11422 9976 11428 9988
rect 6963 9948 11428 9976
rect 6963 9945 6975 9948
rect 6917 9939 6975 9945
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 11790 9936 11796 9988
rect 11848 9976 11854 9988
rect 12452 9976 12480 10084
rect 18325 10081 18337 10115
rect 18371 10112 18383 10115
rect 20438 10112 20444 10124
rect 18371 10084 20444 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 20438 10072 20444 10084
rect 20496 10072 20502 10124
rect 12986 10004 12992 10056
rect 13044 10044 13050 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 13044 10016 13277 10044
rect 13044 10004 13050 10016
rect 13265 10013 13277 10016
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 19797 10047 19855 10053
rect 19797 10013 19809 10047
rect 19843 10044 19855 10047
rect 22002 10044 22008 10056
rect 19843 10016 22008 10044
rect 19843 10013 19855 10016
rect 19797 10007 19855 10013
rect 22002 10004 22008 10016
rect 22060 10004 22066 10056
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10044 22523 10047
rect 23106 10044 23112 10056
rect 22511 10016 23112 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 23106 10004 23112 10016
rect 23164 10004 23170 10056
rect 24578 10004 24584 10056
rect 24636 10044 24642 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 24636 10016 24777 10044
rect 24636 10004 24642 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 25409 10047 25467 10053
rect 25409 10013 25421 10047
rect 25455 10013 25467 10047
rect 25409 10007 25467 10013
rect 11848 9948 12480 9976
rect 11848 9936 11854 9948
rect 14826 9936 14832 9988
rect 14884 9976 14890 9988
rect 17313 9979 17371 9985
rect 17313 9976 17325 9979
rect 14884 9948 17325 9976
rect 14884 9936 14890 9948
rect 17313 9945 17325 9948
rect 17359 9945 17371 9979
rect 17313 9939 17371 9945
rect 17402 9936 17408 9988
rect 17460 9976 17466 9988
rect 25424 9976 25452 10007
rect 36446 10004 36452 10056
rect 36504 10044 36510 10056
rect 38013 10047 38071 10053
rect 38013 10044 38025 10047
rect 36504 10016 38025 10044
rect 36504 10004 36510 10016
rect 38013 10013 38025 10016
rect 38059 10013 38071 10047
rect 38013 10007 38071 10013
rect 17460 9948 17505 9976
rect 24596 9948 25452 9976
rect 17460 9936 17466 9948
rect 1486 9868 1492 9920
rect 1544 9908 1550 9920
rect 1581 9911 1639 9917
rect 1581 9908 1593 9911
rect 1544 9880 1593 9908
rect 1544 9868 1550 9880
rect 1581 9877 1593 9880
rect 1627 9877 1639 9911
rect 4982 9908 4988 9920
rect 4943 9880 4988 9908
rect 1581 9871 1639 9877
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 8481 9911 8539 9917
rect 8481 9877 8493 9911
rect 8527 9908 8539 9911
rect 9214 9908 9220 9920
rect 8527 9880 9220 9908
rect 8527 9877 8539 9880
rect 8481 9871 8539 9877
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 11149 9911 11207 9917
rect 11149 9877 11161 9911
rect 11195 9908 11207 9911
rect 16482 9908 16488 9920
rect 11195 9880 16488 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 24596 9917 24624 9948
rect 24581 9911 24639 9917
rect 24581 9877 24593 9911
rect 24627 9877 24639 9911
rect 38194 9908 38200 9920
rect 38155 9880 38200 9908
rect 24581 9871 24639 9877
rect 38194 9868 38200 9880
rect 38252 9868 38258 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9704 2099 9707
rect 2590 9704 2596 9716
rect 2087 9676 2596 9704
rect 2087 9673 2099 9676
rect 2041 9667 2099 9673
rect 2590 9664 2596 9676
rect 2648 9664 2654 9716
rect 14734 9664 14740 9716
rect 14792 9704 14798 9716
rect 20622 9704 20628 9716
rect 14792 9676 20628 9704
rect 14792 9664 14798 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 20993 9707 21051 9713
rect 20993 9673 21005 9707
rect 21039 9704 21051 9707
rect 21174 9704 21180 9716
rect 21039 9676 21180 9704
rect 21039 9673 21051 9676
rect 20993 9667 21051 9673
rect 21174 9664 21180 9676
rect 21232 9664 21238 9716
rect 8202 9636 8208 9648
rect 3896 9608 7236 9636
rect 8163 9608 8208 9636
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2590 9568 2596 9580
rect 1995 9540 2596 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 2832 9540 2877 9568
rect 2832 9528 2838 9540
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 3896 9432 3924 9608
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9568 4031 9571
rect 4617 9571 4675 9577
rect 4019 9540 4476 9568
rect 4019 9537 4031 9540
rect 3973 9531 4031 9537
rect 4448 9441 4476 9540
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 5258 9568 5264 9580
rect 4663 9540 5264 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 6454 9568 6460 9580
rect 5951 9540 6460 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 5828 9500 5856 9531
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 6546 9528 6552 9580
rect 6604 9568 6610 9580
rect 7208 9577 7236 9608
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 9214 9636 9220 9648
rect 9175 9608 9220 9636
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 10410 9596 10416 9648
rect 10468 9636 10474 9648
rect 11885 9639 11943 9645
rect 11885 9636 11897 9639
rect 10468 9608 11897 9636
rect 10468 9596 10474 9608
rect 11885 9605 11897 9608
rect 11931 9605 11943 9639
rect 11885 9599 11943 9605
rect 30374 9596 30380 9648
rect 30432 9636 30438 9648
rect 32401 9639 32459 9645
rect 32401 9636 32413 9639
rect 30432 9608 32413 9636
rect 30432 9596 30438 9608
rect 32401 9605 32413 9608
rect 32447 9605 32459 9639
rect 32401 9599 32459 9605
rect 7193 9571 7251 9577
rect 6604 9540 6649 9568
rect 6604 9528 6610 9540
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9537 8171 9571
rect 10226 9568 10232 9580
rect 10187 9540 10232 9568
rect 8113 9531 8171 9537
rect 7098 9500 7104 9512
rect 5828 9472 7104 9500
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 2639 9404 3924 9432
rect 4433 9435 4491 9441
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 4433 9401 4445 9435
rect 4479 9401 4491 9435
rect 4433 9395 4491 9401
rect 5810 9392 5816 9444
rect 5868 9432 5874 9444
rect 8128 9432 8156 9531
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9568 19763 9571
rect 24118 9568 24124 9580
rect 19751 9540 24124 9568
rect 19751 9537 19763 9540
rect 19705 9531 19763 9537
rect 24118 9528 24124 9540
rect 24176 9528 24182 9580
rect 32309 9571 32367 9577
rect 32309 9537 32321 9571
rect 32355 9568 32367 9571
rect 34238 9568 34244 9580
rect 32355 9540 34244 9568
rect 32355 9537 32367 9540
rect 32309 9531 32367 9537
rect 34238 9528 34244 9540
rect 34296 9528 34302 9580
rect 34885 9571 34943 9577
rect 34885 9568 34897 9571
rect 34348 9540 34897 9568
rect 34348 9512 34376 9540
rect 34885 9537 34897 9540
rect 34931 9537 34943 9571
rect 34885 9531 34943 9537
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9500 9183 9503
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 9171 9472 10517 9500
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 11793 9503 11851 9509
rect 11793 9500 11805 9503
rect 11112 9472 11805 9500
rect 11112 9460 11118 9472
rect 11793 9469 11805 9472
rect 11839 9500 11851 9503
rect 12066 9500 12072 9512
rect 11839 9472 12072 9500
rect 11839 9469 11851 9472
rect 11793 9463 11851 9469
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 20349 9503 20407 9509
rect 20349 9469 20361 9503
rect 20395 9500 20407 9503
rect 20438 9500 20444 9512
rect 20395 9472 20444 9500
rect 20395 9469 20407 9472
rect 20349 9463 20407 9469
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 20533 9503 20591 9509
rect 20533 9469 20545 9503
rect 20579 9500 20591 9503
rect 20806 9500 20812 9512
rect 20579 9472 20812 9500
rect 20579 9469 20591 9472
rect 20533 9463 20591 9469
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 34330 9500 34336 9512
rect 34291 9472 34336 9500
rect 34330 9460 34336 9472
rect 34388 9460 34394 9512
rect 5868 9404 8156 9432
rect 5868 9392 5874 9404
rect 8478 9392 8484 9444
rect 8536 9432 8542 9444
rect 9677 9435 9735 9441
rect 9677 9432 9689 9435
rect 8536 9404 9689 9432
rect 8536 9392 8542 9404
rect 9677 9401 9689 9404
rect 9723 9432 9735 9435
rect 12345 9435 12403 9441
rect 12345 9432 12357 9435
rect 9723 9404 12357 9432
rect 9723 9401 9735 9404
rect 9677 9395 9735 9401
rect 12345 9401 12357 9404
rect 12391 9401 12403 9435
rect 12345 9395 12403 9401
rect 34701 9435 34759 9441
rect 34701 9401 34713 9435
rect 34747 9432 34759 9435
rect 36446 9432 36452 9444
rect 34747 9404 36452 9432
rect 34747 9401 34759 9404
rect 34701 9395 34759 9401
rect 36446 9392 36452 9404
rect 36504 9392 36510 9444
rect 3786 9364 3792 9376
rect 3747 9336 3792 9364
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 6638 9364 6644 9376
rect 6599 9336 6644 9364
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 11790 9364 11796 9376
rect 7331 9336 11796 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 19797 9367 19855 9373
rect 19797 9364 19809 9367
rect 19392 9336 19809 9364
rect 19392 9324 19398 9336
rect 19797 9333 19809 9336
rect 19843 9333 19855 9367
rect 19797 9327 19855 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 6822 9160 6828 9172
rect 1627 9132 6828 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 9217 9163 9275 9169
rect 9217 9129 9229 9163
rect 9263 9160 9275 9163
rect 10134 9160 10140 9172
rect 9263 9132 10140 9160
rect 9263 9129 9275 9132
rect 9217 9123 9275 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 11425 9163 11483 9169
rect 11425 9129 11437 9163
rect 11471 9160 11483 9163
rect 11606 9160 11612 9172
rect 11471 9132 11612 9160
rect 11471 9129 11483 9132
rect 11425 9123 11483 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 12066 9160 12072 9172
rect 12027 9132 12072 9160
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 26326 9160 26332 9172
rect 26287 9132 26332 9160
rect 26326 9120 26332 9132
rect 26384 9120 26390 9172
rect 2317 9095 2375 9101
rect 2317 9061 2329 9095
rect 2363 9092 2375 9095
rect 2498 9092 2504 9104
rect 2363 9064 2504 9092
rect 2363 9061 2375 9064
rect 2317 9055 2375 9061
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 3418 9052 3424 9104
rect 3476 9092 3482 9104
rect 5445 9095 5503 9101
rect 5445 9092 5457 9095
rect 3476 9064 5457 9092
rect 3476 9052 3482 9064
rect 5445 9061 5457 9064
rect 5491 9061 5503 9095
rect 5445 9055 5503 9061
rect 2866 9024 2872 9036
rect 1780 8996 2872 9024
rect 1780 8965 1808 8996
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 20438 9024 20444 9036
rect 20399 8996 20444 9024
rect 20438 8984 20444 8996
rect 20496 8984 20502 9036
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 2222 8956 2228 8968
rect 2183 8928 2228 8956
rect 1765 8919 1823 8925
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4982 8956 4988 8968
rect 4203 8928 4988 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8956 5687 8959
rect 6638 8956 6644 8968
rect 5675 8928 6644 8956
rect 5675 8925 5687 8928
rect 5629 8919 5687 8925
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 9122 8956 9128 8968
rect 9083 8928 9128 8956
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 11330 8956 11336 8968
rect 11291 8928 11336 8956
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 13170 8956 13176 8968
rect 12023 8928 13176 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 23842 8916 23848 8968
rect 23900 8956 23906 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 23900 8928 24593 8956
rect 23900 8916 23906 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 26326 8956 26332 8968
rect 26287 8928 26332 8956
rect 24581 8919 24639 8925
rect 26326 8916 26332 8928
rect 26384 8916 26390 8968
rect 32582 8956 32588 8968
rect 32543 8928 32588 8956
rect 32582 8916 32588 8928
rect 32640 8916 32646 8968
rect 2866 8820 2872 8832
rect 2827 8792 2872 8820
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3973 8823 4031 8829
rect 3973 8820 3985 8823
rect 3108 8792 3985 8820
rect 3108 8780 3114 8792
rect 3973 8789 3985 8792
rect 4019 8789 4031 8823
rect 4614 8820 4620 8832
rect 4575 8792 4620 8820
rect 3973 8783 4031 8789
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 24673 8823 24731 8829
rect 24673 8789 24685 8823
rect 24719 8820 24731 8823
rect 24762 8820 24768 8832
rect 24719 8792 24768 8820
rect 24719 8789 24731 8792
rect 24673 8783 24731 8789
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 32401 8823 32459 8829
rect 32401 8789 32413 8823
rect 32447 8820 32459 8823
rect 34146 8820 34152 8832
rect 32447 8792 34152 8820
rect 32447 8789 32459 8792
rect 32401 8783 32459 8789
rect 34146 8780 34152 8792
rect 34204 8780 34210 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1946 8576 1952 8628
rect 2004 8616 2010 8628
rect 2225 8619 2283 8625
rect 2225 8616 2237 8619
rect 2004 8588 2237 8616
rect 2004 8576 2010 8588
rect 2225 8585 2237 8588
rect 2271 8585 2283 8619
rect 3510 8616 3516 8628
rect 3471 8588 3516 8616
rect 2225 8579 2283 8585
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 5166 8616 5172 8628
rect 4663 8588 5172 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 2866 8480 2872 8492
rect 2827 8452 2872 8480
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3050 8480 3056 8492
rect 3011 8452 3056 8480
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8480 4031 8483
rect 4614 8480 4620 8492
rect 4019 8452 4620 8480
rect 4019 8449 4031 8452
rect 3973 8443 4031 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8480 14611 8483
rect 15194 8480 15200 8492
rect 14599 8452 15200 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 20990 8480 20996 8492
rect 20951 8452 20996 8480
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 27062 8440 27068 8492
rect 27120 8480 27126 8492
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 27120 8452 27169 8480
rect 27120 8440 27126 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 38102 8480 38108 8492
rect 38063 8452 38108 8480
rect 27157 8443 27215 8449
rect 38102 8440 38108 8452
rect 38160 8440 38166 8492
rect 3786 8372 3792 8424
rect 3844 8412 3850 8424
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 3844 8384 4169 8412
rect 3844 8372 3850 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 38289 8415 38347 8421
rect 38289 8412 38301 8415
rect 13320 8384 38301 8412
rect 13320 8372 13326 8384
rect 38289 8381 38301 8384
rect 38335 8381 38347 8415
rect 38289 8375 38347 8381
rect 12434 8304 12440 8356
rect 12492 8344 12498 8356
rect 14645 8347 14703 8353
rect 14645 8344 14657 8347
rect 12492 8316 14657 8344
rect 12492 8304 12498 8316
rect 14645 8313 14657 8316
rect 14691 8313 14703 8347
rect 14645 8307 14703 8313
rect 27249 8347 27307 8353
rect 27249 8313 27261 8347
rect 27295 8344 27307 8347
rect 28902 8344 28908 8356
rect 27295 8316 28908 8344
rect 27295 8313 27307 8316
rect 27249 8307 27307 8313
rect 28902 8304 28908 8316
rect 28960 8304 28966 8356
rect 20809 8279 20867 8285
rect 20809 8245 20821 8279
rect 20855 8276 20867 8279
rect 20990 8276 20996 8288
rect 20855 8248 20996 8276
rect 20855 8245 20867 8248
rect 20809 8239 20867 8245
rect 20990 8236 20996 8248
rect 21048 8236 21054 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 3326 8032 3332 8084
rect 3384 8072 3390 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3384 8044 4077 8072
rect 3384 8032 3390 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 14826 8072 14832 8084
rect 14787 8044 14832 8072
rect 4065 8035 4123 8041
rect 14826 8032 14832 8044
rect 14884 8032 14890 8084
rect 20806 8072 20812 8084
rect 20767 8044 20812 8072
rect 20806 8032 20812 8044
rect 20864 8032 20870 8084
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 9122 7936 9128 7948
rect 1903 7908 9128 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 9122 7896 9128 7908
rect 9180 7896 9186 7948
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7868 3203 7871
rect 3510 7868 3516 7880
rect 3191 7840 3516 7868
rect 3191 7837 3203 7840
rect 3145 7831 3203 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 3970 7868 3976 7880
rect 3931 7840 3976 7868
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 12434 7868 12440 7880
rect 11103 7840 12440 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 12434 7828 12440 7840
rect 12492 7828 12498 7880
rect 14734 7868 14740 7880
rect 14695 7840 14740 7868
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19334 7868 19340 7880
rect 18923 7840 19340 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 20990 7868 20996 7880
rect 20951 7840 20996 7868
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 24762 7868 24768 7880
rect 24723 7840 24768 7868
rect 24762 7828 24768 7840
rect 24820 7828 24826 7880
rect 28902 7828 28908 7880
rect 28960 7868 28966 7880
rect 29181 7871 29239 7877
rect 29181 7868 29193 7871
rect 28960 7840 29193 7868
rect 28960 7828 28966 7840
rect 29181 7837 29193 7840
rect 29227 7837 29239 7871
rect 29181 7831 29239 7837
rect 33134 7828 33140 7880
rect 33192 7868 33198 7880
rect 33781 7871 33839 7877
rect 33781 7868 33793 7871
rect 33192 7840 33793 7868
rect 33192 7828 33198 7840
rect 33781 7837 33793 7840
rect 33827 7837 33839 7871
rect 33781 7831 33839 7837
rect 34146 7828 34152 7880
rect 34204 7868 34210 7880
rect 38013 7871 38071 7877
rect 38013 7868 38025 7871
rect 34204 7840 38025 7868
rect 34204 7828 34210 7840
rect 38013 7837 38025 7840
rect 38059 7837 38071 7871
rect 38013 7831 38071 7837
rect 3234 7732 3240 7744
rect 3195 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 6822 7692 6828 7744
rect 6880 7732 6886 7744
rect 10873 7735 10931 7741
rect 10873 7732 10885 7735
rect 6880 7704 10885 7732
rect 6880 7692 6886 7704
rect 10873 7701 10885 7704
rect 10919 7701 10931 7735
rect 10873 7695 10931 7701
rect 17494 7692 17500 7744
rect 17552 7732 17558 7744
rect 18693 7735 18751 7741
rect 18693 7732 18705 7735
rect 17552 7704 18705 7732
rect 17552 7692 17558 7704
rect 18693 7701 18705 7704
rect 18739 7701 18751 7735
rect 18693 7695 18751 7701
rect 24581 7735 24639 7741
rect 24581 7701 24593 7735
rect 24627 7732 24639 7735
rect 25958 7732 25964 7744
rect 24627 7704 25964 7732
rect 24627 7701 24639 7704
rect 24581 7695 24639 7701
rect 25958 7692 25964 7704
rect 26016 7692 26022 7744
rect 28997 7735 29055 7741
rect 28997 7701 29009 7735
rect 29043 7732 29055 7735
rect 31662 7732 31668 7744
rect 29043 7704 31668 7732
rect 29043 7701 29055 7704
rect 28997 7695 29055 7701
rect 31662 7692 31668 7704
rect 31720 7692 31726 7744
rect 33873 7735 33931 7741
rect 33873 7701 33885 7735
rect 33919 7732 33931 7735
rect 34790 7732 34796 7744
rect 33919 7704 34796 7732
rect 33919 7701 33931 7704
rect 33873 7695 33931 7701
rect 34790 7692 34796 7704
rect 34848 7692 34854 7744
rect 38194 7732 38200 7744
rect 38155 7704 38200 7732
rect 38194 7692 38200 7704
rect 38252 7692 38258 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1854 7420 1860 7472
rect 1912 7460 1918 7472
rect 2409 7463 2467 7469
rect 2409 7460 2421 7463
rect 1912 7432 2421 7460
rect 1912 7420 1918 7432
rect 2409 7429 2421 7432
rect 2455 7429 2467 7463
rect 2409 7423 2467 7429
rect 2501 7463 2559 7469
rect 2501 7429 2513 7463
rect 2547 7460 2559 7463
rect 2866 7460 2872 7472
rect 2547 7432 2872 7460
rect 2547 7429 2559 7432
rect 2501 7423 2559 7429
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 3292 7364 4629 7392
rect 3292 7352 3298 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 9122 7352 9128 7404
rect 9180 7392 9186 7404
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 9180 7364 14197 7392
rect 9180 7352 9186 7364
rect 14185 7361 14197 7364
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7392 16911 7395
rect 21082 7392 21088 7404
rect 16899 7364 21088 7392
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 34422 7352 34428 7404
rect 34480 7392 34486 7404
rect 35069 7395 35127 7401
rect 35069 7392 35081 7395
rect 34480 7364 35081 7392
rect 34480 7352 34486 7364
rect 35069 7361 35081 7364
rect 35115 7361 35127 7395
rect 35069 7355 35127 7361
rect 2958 7256 2964 7268
rect 2919 7228 2964 7256
rect 2958 7216 2964 7228
rect 3016 7216 3022 7268
rect 12894 7256 12900 7268
rect 4356 7228 12900 7256
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7188 1823 7191
rect 4356 7188 4384 7228
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 14001 7259 14059 7265
rect 14001 7225 14013 7259
rect 14047 7256 14059 7259
rect 19978 7256 19984 7268
rect 14047 7228 19984 7256
rect 14047 7225 14059 7228
rect 14001 7219 14059 7225
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 1811 7160 4384 7188
rect 4433 7191 4491 7197
rect 1811 7157 1823 7160
rect 1765 7151 1823 7157
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4614 7188 4620 7200
rect 4479 7160 4620 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 16945 7191 17003 7197
rect 16945 7157 16957 7191
rect 16991 7188 17003 7191
rect 17034 7188 17040 7200
rect 16991 7160 17040 7188
rect 16991 7157 17003 7160
rect 16945 7151 17003 7157
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 34885 7191 34943 7197
rect 34885 7157 34897 7191
rect 34931 7188 34943 7191
rect 37734 7188 37740 7200
rect 34931 7160 37740 7188
rect 34931 7157 34943 7160
rect 34885 7151 34943 7157
rect 37734 7148 37740 7160
rect 37792 7148 37798 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 2314 6848 2320 6860
rect 2275 6820 2320 6848
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6749 1823 6783
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 1765 6743 1823 6749
rect 1780 6712 1808 6743
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 34790 6740 34796 6792
rect 34848 6780 34854 6792
rect 35069 6783 35127 6789
rect 35069 6780 35081 6783
rect 34848 6752 35081 6780
rect 34848 6740 34854 6752
rect 35069 6749 35081 6752
rect 35115 6749 35127 6783
rect 35069 6743 35127 6749
rect 2774 6712 2780 6724
rect 1780 6684 2780 6712
rect 2774 6672 2780 6684
rect 2832 6672 2838 6724
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2130 6644 2136 6656
rect 1627 6616 2136 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 34885 6647 34943 6653
rect 34885 6613 34897 6647
rect 34931 6644 34943 6647
rect 38010 6644 38016 6656
rect 34931 6616 38016 6644
rect 34931 6613 34943 6616
rect 34885 6607 34943 6613
rect 38010 6604 38016 6616
rect 38068 6604 38074 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 37737 6307 37795 6313
rect 37737 6304 37749 6307
rect 26206 6276 37749 6304
rect 15194 6236 15200 6248
rect 15155 6208 15200 6236
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 24486 6196 24492 6248
rect 24544 6236 24550 6248
rect 26206 6236 26234 6276
rect 37737 6273 37749 6276
rect 37783 6273 37795 6307
rect 37737 6267 37795 6273
rect 37458 6236 37464 6248
rect 24544 6208 26234 6236
rect 37419 6208 37464 6236
rect 24544 6196 24550 6208
rect 37458 6196 37464 6208
rect 37516 6196 37522 6248
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 2866 5896 2872 5908
rect 2827 5868 2872 5896
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 14550 5788 14556 5840
rect 14608 5828 14614 5840
rect 14608 5800 15516 5828
rect 14608 5788 14614 5800
rect 15194 5760 15200 5772
rect 15155 5732 15200 5760
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 15488 5769 15516 5800
rect 15473 5763 15531 5769
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 15519 5732 16574 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1544 5664 1593 5692
rect 1544 5652 1550 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 3602 5692 3608 5704
rect 2823 5664 3608 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 5442 5692 5448 5704
rect 4479 5664 5448 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 16546 5692 16574 5732
rect 23845 5695 23903 5701
rect 23845 5692 23857 5695
rect 16546 5664 23857 5692
rect 23845 5661 23857 5664
rect 23891 5661 23903 5695
rect 23845 5655 23903 5661
rect 15286 5584 15292 5636
rect 15344 5624 15350 5636
rect 15344 5596 15389 5624
rect 15344 5584 15350 5596
rect 1762 5556 1768 5568
rect 1723 5528 1768 5556
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 4525 5559 4583 5565
rect 4525 5525 4537 5559
rect 4571 5556 4583 5559
rect 4706 5556 4712 5568
rect 4571 5528 4712 5556
rect 4571 5525 4583 5528
rect 4525 5519 4583 5525
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 23937 5559 23995 5565
rect 23937 5525 23949 5559
rect 23983 5556 23995 5559
rect 24762 5556 24768 5568
rect 23983 5528 24768 5556
rect 23983 5525 23995 5528
rect 23937 5519 23995 5525
rect 24762 5516 24768 5528
rect 24820 5516 24826 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 4706 5216 4712 5228
rect 4667 5188 4712 5216
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 11698 5216 11704 5228
rect 9539 5188 11704 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 24762 5216 24768 5228
rect 24723 5188 24768 5216
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 38010 5216 38016 5228
rect 37971 5188 38016 5216
rect 38010 5176 38016 5188
rect 38068 5176 38074 5228
rect 4525 5015 4583 5021
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 4614 5012 4620 5024
rect 4571 4984 4620 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 9309 5015 9367 5021
rect 9309 4981 9321 5015
rect 9355 5012 9367 5015
rect 11698 5012 11704 5024
rect 9355 4984 11704 5012
rect 9355 4981 9367 4984
rect 9309 4975 9367 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 24581 5015 24639 5021
rect 24581 4981 24593 5015
rect 24627 5012 24639 5015
rect 30466 5012 30472 5024
rect 24627 4984 30472 5012
rect 24627 4981 24639 4984
rect 24581 4975 24639 4981
rect 30466 4972 30472 4984
rect 30524 4972 30530 5024
rect 38194 5012 38200 5024
rect 38155 4984 38200 5012
rect 38194 4972 38200 4984
rect 38252 4972 38258 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 32122 4564 32128 4616
rect 32180 4604 32186 4616
rect 33137 4607 33195 4613
rect 33137 4604 33149 4607
rect 32180 4576 33149 4604
rect 32180 4564 32186 4576
rect 33137 4573 33149 4576
rect 33183 4573 33195 4607
rect 33137 4567 33195 4573
rect 33229 4607 33287 4613
rect 33229 4573 33241 4607
rect 33275 4604 33287 4607
rect 35529 4607 35587 4613
rect 35529 4604 35541 4607
rect 33275 4576 35541 4604
rect 33275 4573 33287 4576
rect 33229 4567 33287 4573
rect 35529 4573 35541 4576
rect 35575 4573 35587 4607
rect 35529 4567 35587 4573
rect 37734 4564 37740 4616
rect 37792 4604 37798 4616
rect 38013 4607 38071 4613
rect 38013 4604 38025 4607
rect 37792 4576 38025 4604
rect 37792 4564 37798 4576
rect 38013 4573 38025 4576
rect 38059 4573 38071 4607
rect 38013 4567 38071 4573
rect 1670 4536 1676 4548
rect 1631 4508 1676 4536
rect 1670 4496 1676 4508
rect 1728 4496 1734 4548
rect 1765 4471 1823 4477
rect 1765 4437 1777 4471
rect 1811 4468 1823 4471
rect 12158 4468 12164 4480
rect 1811 4440 12164 4468
rect 1811 4437 1823 4440
rect 1765 4431 1823 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 35342 4468 35348 4480
rect 35303 4440 35348 4468
rect 35342 4428 35348 4440
rect 35400 4428 35406 4480
rect 38194 4468 38200 4480
rect 38155 4440 38200 4468
rect 38194 4428 38200 4440
rect 38252 4428 38258 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 37918 4088 37924 4140
rect 37976 4128 37982 4140
rect 38013 4131 38071 4137
rect 38013 4128 38025 4131
rect 37976 4100 38025 4128
rect 37976 4088 37982 4100
rect 38013 4097 38025 4100
rect 38059 4097 38071 4131
rect 38013 4091 38071 4097
rect 38197 3927 38255 3933
rect 38197 3893 38209 3927
rect 38243 3924 38255 3927
rect 39298 3924 39304 3936
rect 38243 3896 39304 3924
rect 38243 3893 38255 3896
rect 38197 3887 38255 3893
rect 39298 3884 39304 3896
rect 39356 3884 39362 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 2222 3720 2228 3732
rect 1627 3692 2228 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 37826 3544 37832 3596
rect 37884 3584 37890 3596
rect 37884 3556 38056 3584
rect 37884 3544 37890 3556
rect 1762 3516 1768 3528
rect 1723 3488 1768 3516
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 37553 3519 37611 3525
rect 37553 3485 37565 3519
rect 37599 3516 37611 3519
rect 37918 3516 37924 3528
rect 37599 3488 37924 3516
rect 37599 3485 37611 3488
rect 37553 3479 37611 3485
rect 37918 3476 37924 3488
rect 37976 3476 37982 3528
rect 38028 3525 38056 3556
rect 38013 3519 38071 3525
rect 38013 3485 38025 3519
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 27982 3340 27988 3392
rect 28040 3380 28046 3392
rect 37369 3383 37427 3389
rect 37369 3380 37381 3383
rect 28040 3352 37381 3380
rect 28040 3340 28046 3352
rect 37369 3349 37381 3352
rect 37415 3349 37427 3383
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 37369 3343 37427 3349
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3176 2375 3179
rect 3970 3176 3976 3188
rect 2363 3148 3976 3176
rect 2363 3145 2375 3148
rect 2317 3139 2375 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 34238 3136 34244 3188
rect 34296 3176 34302 3188
rect 36725 3179 36783 3185
rect 36725 3176 36737 3179
rect 34296 3148 36737 3176
rect 34296 3136 34302 3148
rect 36725 3145 36737 3148
rect 36771 3145 36783 3179
rect 36725 3139 36783 3145
rect 4614 3108 4620 3120
rect 1596 3080 4620 3108
rect 1596 3049 1624 3080
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 13170 3068 13176 3120
rect 13228 3108 13234 3120
rect 37274 3108 37280 3120
rect 13228 3080 18920 3108
rect 13228 3068 13234 3080
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 1946 3000 1952 3052
rect 2004 3040 2010 3052
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2004 3012 2513 3040
rect 2004 3000 2010 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 3234 3000 3240 3052
rect 3292 3040 3298 3052
rect 3513 3043 3571 3049
rect 3513 3040 3525 3043
rect 3292 3012 3525 3040
rect 3292 3000 3298 3012
rect 3513 3009 3525 3012
rect 3559 3009 3571 3043
rect 11974 3040 11980 3052
rect 11935 3012 11980 3040
rect 3513 3003 3571 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 18892 3049 18920 3080
rect 26206 3080 37280 3108
rect 18877 3043 18935 3049
rect 18877 3009 18889 3043
rect 18923 3009 18935 3043
rect 25774 3040 25780 3052
rect 25735 3012 25780 3040
rect 18877 3003 18935 3009
rect 25774 3000 25780 3012
rect 25832 3040 25838 3052
rect 26206 3040 26234 3080
rect 37274 3068 37280 3080
rect 37332 3068 37338 3120
rect 25832 3012 26234 3040
rect 25832 3000 25838 3012
rect 36722 3000 36728 3052
rect 36780 3040 36786 3052
rect 36909 3043 36967 3049
rect 36909 3040 36921 3043
rect 36780 3012 36921 3040
rect 36780 3000 36786 3012
rect 36909 3009 36921 3012
rect 36955 3009 36967 3043
rect 37737 3043 37795 3049
rect 37737 3040 37749 3043
rect 36909 3003 36967 3009
rect 37016 3012 37749 3040
rect 11606 2932 11612 2984
rect 11664 2972 11670 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 11664 2944 11713 2972
rect 11664 2932 11670 2944
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 28442 2932 28448 2984
rect 28500 2972 28506 2984
rect 37016 2972 37044 3012
rect 37737 3009 37749 3012
rect 37783 3009 37795 3043
rect 37737 3003 37795 3009
rect 37458 2972 37464 2984
rect 28500 2944 37044 2972
rect 37419 2944 37464 2972
rect 28500 2932 28506 2944
rect 37458 2932 37464 2944
rect 37516 2932 37522 2984
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2904 3387 2907
rect 11146 2904 11152 2916
rect 3375 2876 11152 2904
rect 3375 2873 3387 2876
rect 3329 2867 3387 2873
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 716 2808 1777 2836
rect 716 2796 722 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 16850 2836 16856 2848
rect 16811 2808 16856 2836
rect 1765 2799 1823 2805
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 18693 2839 18751 2845
rect 18693 2805 18705 2839
rect 18739 2836 18751 2839
rect 20622 2836 20628 2848
rect 18739 2808 20628 2836
rect 18739 2805 18751 2808
rect 18693 2799 18751 2805
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 25222 2796 25228 2848
rect 25280 2836 25286 2848
rect 25593 2839 25651 2845
rect 25593 2836 25605 2839
rect 25280 2808 25605 2836
rect 25280 2796 25286 2808
rect 25593 2805 25605 2808
rect 25639 2805 25651 2839
rect 25593 2799 25651 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7193 2635 7251 2641
rect 7193 2632 7205 2635
rect 7156 2604 7205 2632
rect 7156 2592 7162 2604
rect 7193 2601 7205 2604
rect 7239 2601 7251 2635
rect 7193 2595 7251 2601
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 10226 2632 10232 2644
rect 9815 2604 10232 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 14734 2632 14740 2644
rect 14323 2604 14740 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 18230 2632 18236 2644
rect 18191 2604 18236 2632
rect 18230 2592 18236 2604
rect 18288 2592 18294 2644
rect 22002 2632 22008 2644
rect 21963 2604 22008 2632
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 24581 2635 24639 2641
rect 24581 2601 24593 2635
rect 24627 2632 24639 2635
rect 24670 2632 24676 2644
rect 24627 2604 24676 2632
rect 24627 2601 24639 2604
rect 24581 2595 24639 2601
rect 24670 2592 24676 2604
rect 24728 2592 24734 2644
rect 26326 2592 26332 2644
rect 26384 2632 26390 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 26384 2604 27169 2632
rect 26384 2592 26390 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27157 2595 27215 2601
rect 27430 2592 27436 2644
rect 27488 2632 27494 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 27488 2604 28641 2632
rect 27488 2592 27494 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 28629 2595 28687 2601
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 3237 2567 3295 2573
rect 3237 2564 3249 2567
rect 72 2536 3249 2564
rect 72 2524 78 2536
rect 3237 2533 3249 2536
rect 3283 2533 3295 2567
rect 22278 2564 22284 2576
rect 3237 2527 3295 2533
rect 6886 2536 22284 2564
rect 4706 2496 4712 2508
rect 3068 2468 4712 2496
rect 3068 2437 3096 2468
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 6886 2496 6914 2536
rect 22278 2524 22284 2536
rect 22336 2524 22342 2576
rect 31570 2524 31576 2576
rect 31628 2564 31634 2576
rect 31628 2536 34928 2564
rect 31628 2524 31634 2536
rect 5276 2468 6914 2496
rect 5276 2437 5304 2468
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 13170 2496 13176 2508
rect 8536 2468 13032 2496
rect 13131 2468 13176 2496
rect 8536 2456 8542 2468
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 5031 2400 5273 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 1670 2360 1676 2372
rect 1631 2332 1676 2360
rect 1670 2320 1676 2332
rect 1728 2320 1734 2372
rect 2332 2360 2360 2391
rect 3418 2360 3424 2372
rect 2332 2332 3424 2360
rect 3418 2320 3424 2332
rect 3476 2320 3482 2372
rect 3988 2360 4016 2391
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6512 2400 6745 2428
rect 6512 2388 6518 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7156 2400 7389 2428
rect 7156 2388 7162 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 8444 2400 9321 2428
rect 8444 2388 8450 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9732 2400 9965 2428
rect 9732 2388 9738 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 11698 2428 11704 2440
rect 11659 2400 11704 2428
rect 9953 2391 10011 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 12894 2428 12900 2440
rect 12855 2400 12900 2428
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13004 2428 13032 2468
rect 13170 2456 13176 2468
rect 13228 2456 13234 2508
rect 19705 2499 19763 2505
rect 19705 2496 19717 2499
rect 13280 2468 19717 2496
rect 13280 2428 13308 2468
rect 19705 2465 19717 2468
rect 19751 2465 19763 2499
rect 19705 2459 19763 2465
rect 20622 2456 20628 2508
rect 20680 2496 20686 2508
rect 20680 2468 22692 2496
rect 20680 2456 20686 2468
rect 13004 2400 13308 2428
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 14240 2400 14473 2428
rect 14240 2388 14246 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2428 16083 2431
rect 16850 2428 16856 2440
rect 16071 2400 16856 2428
rect 16071 2397 16083 2400
rect 16025 2391 16083 2397
rect 6822 2360 6828 2372
rect 3988 2332 6828 2360
rect 6822 2320 6828 2332
rect 6880 2320 6886 2372
rect 11330 2360 11336 2372
rect 9140 2332 11336 2360
rect 1762 2292 1768 2304
rect 1723 2264 1768 2292
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3936 2264 4169 2292
rect 3936 2252 3942 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5224 2264 5457 2292
rect 5224 2252 5230 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 6549 2295 6607 2301
rect 6549 2261 6561 2295
rect 6595 2292 6607 2295
rect 9030 2292 9036 2304
rect 6595 2264 9036 2292
rect 6595 2261 6607 2264
rect 6549 2255 6607 2261
rect 9030 2252 9036 2264
rect 9088 2252 9094 2304
rect 9140 2301 9168 2332
rect 11330 2320 11336 2332
rect 11388 2320 11394 2372
rect 14936 2360 14964 2391
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18417 2431 18475 2437
rect 18417 2428 18429 2431
rect 18104 2400 18429 2428
rect 18104 2388 18110 2400
rect 18417 2397 18429 2400
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19392 2400 19441 2428
rect 19392 2388 19398 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 20036 2400 20729 2428
rect 20036 2388 20042 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22664 2437 22692 2468
rect 24854 2456 24860 2508
rect 24912 2496 24918 2508
rect 24912 2468 33824 2496
rect 24912 2456 24918 2468
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21968 2400 22201 2428
rect 21968 2388 21974 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 23900 2400 24777 2428
rect 23900 2388 23906 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 25222 2428 25228 2440
rect 25183 2400 25228 2428
rect 24765 2391 24823 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 25958 2428 25964 2440
rect 25919 2400 25964 2428
rect 25958 2388 25964 2400
rect 26016 2388 26022 2440
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 29730 2428 29736 2440
rect 29691 2400 29736 2428
rect 27341 2391 27399 2397
rect 29730 2388 29736 2400
rect 29788 2388 29794 2440
rect 30466 2428 30472 2440
rect 30427 2400 30472 2428
rect 30466 2388 30472 2400
rect 30524 2388 30530 2440
rect 31662 2388 31668 2440
rect 31720 2428 31726 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31720 2400 32321 2428
rect 31720 2388 31726 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33045 2431 33103 2437
rect 33045 2397 33057 2431
rect 33091 2428 33103 2431
rect 33318 2428 33324 2440
rect 33091 2400 33324 2428
rect 33091 2397 33103 2400
rect 33045 2391 33103 2397
rect 33318 2388 33324 2400
rect 33376 2388 33382 2440
rect 33796 2437 33824 2468
rect 34900 2437 34928 2536
rect 37274 2456 37280 2508
rect 37332 2496 37338 2508
rect 37737 2499 37795 2505
rect 37737 2496 37749 2499
rect 37332 2468 37749 2496
rect 37332 2456 37338 2468
rect 37737 2465 37749 2468
rect 37783 2465 37795 2499
rect 37737 2459 37795 2465
rect 33781 2431 33839 2437
rect 33781 2397 33793 2431
rect 33827 2397 33839 2431
rect 33781 2391 33839 2397
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35342 2388 35348 2440
rect 35400 2428 35406 2440
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 35400 2400 36185 2428
rect 35400 2388 35406 2400
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 37458 2428 37464 2440
rect 37419 2400 37464 2428
rect 36173 2391 36231 2397
rect 37458 2388 37464 2400
rect 37516 2388 37522 2440
rect 27798 2360 27804 2372
rect 14936 2332 27804 2360
rect 27798 2320 27804 2332
rect 27856 2320 27862 2372
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28537 2363 28595 2369
rect 28537 2360 28549 2363
rect 28408 2332 28549 2360
rect 28408 2320 28414 2332
rect 28537 2329 28549 2332
rect 28583 2329 28595 2363
rect 28537 2323 28595 2329
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11020 2264 11897 2292
rect 11020 2252 11026 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14884 2264 15117 2292
rect 14884 2252 14890 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16209 2295 16267 2301
rect 16209 2292 16221 2295
rect 16172 2264 16221 2292
rect 16172 2252 16178 2264
rect 16209 2261 16221 2264
rect 16255 2261 16267 2295
rect 16209 2255 16267 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20680 2264 20913 2292
rect 20680 2252 20686 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 22833 2255 22891 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26145 2295 26203 2301
rect 26145 2292 26157 2295
rect 25832 2264 26157 2292
rect 25832 2252 25838 2264
rect 26145 2261 26157 2264
rect 26191 2261 26203 2295
rect 26145 2255 26203 2261
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 29696 2264 29929 2292
rect 29696 2252 29702 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 29917 2255 29975 2261
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 30653 2295 30711 2301
rect 30653 2292 30665 2295
rect 30340 2264 30665 2292
rect 30340 2252 30346 2264
rect 30653 2261 30665 2264
rect 30699 2261 30711 2295
rect 30653 2255 30711 2261
rect 31570 2252 31576 2304
rect 31628 2292 31634 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 31628 2264 32505 2292
rect 31628 2252 31634 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 32858 2252 32864 2304
rect 32916 2292 32922 2304
rect 33229 2295 33287 2301
rect 33229 2292 33241 2295
rect 32916 2264 33241 2292
rect 32916 2252 32922 2264
rect 33229 2261 33241 2264
rect 33275 2261 33287 2295
rect 33229 2255 33287 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33965 2295 34023 2301
rect 33965 2292 33977 2295
rect 33560 2264 33977 2292
rect 33560 2252 33566 2264
rect 33965 2261 33977 2264
rect 34011 2261 34023 2295
rect 33965 2255 34023 2261
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34848 2264 35081 2292
rect 34848 2252 34854 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 36078 2252 36084 2304
rect 36136 2292 36142 2304
rect 36357 2295 36415 2301
rect 36357 2292 36369 2295
rect 36136 2264 36369 2292
rect 36136 2252 36142 2264
rect 36357 2261 36369 2264
rect 36403 2261 36415 2295
rect 36357 2255 36415 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 9030 2048 9036 2100
rect 9088 2088 9094 2100
rect 12986 2088 12992 2100
rect 9088 2060 12992 2088
rect 9088 2048 9094 2060
rect 12986 2048 12992 2060
rect 13044 2048 13050 2100
rect 1762 1980 1768 2032
rect 1820 2020 1826 2032
rect 15010 2020 15016 2032
rect 1820 1992 15016 2020
rect 1820 1980 1826 1992
rect 15010 1980 15016 1992
rect 15068 1980 15074 2032
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1768 37451 1820 37460
rect 1768 37417 1777 37451
rect 1777 37417 1811 37451
rect 1811 37417 1820 37451
rect 1768 37408 1820 37417
rect 25044 37408 25096 37460
rect 6092 37340 6144 37392
rect 25412 37340 25464 37392
rect 26240 37340 26292 37392
rect 12256 37272 12308 37324
rect 2320 37204 2372 37256
rect 2780 37204 2832 37256
rect 2964 37204 3016 37256
rect 4620 37204 4672 37256
rect 6460 37204 6512 37256
rect 6552 37247 6604 37256
rect 6552 37213 6561 37247
rect 6561 37213 6595 37247
rect 6595 37213 6604 37247
rect 6552 37204 6604 37213
rect 7748 37204 7800 37256
rect 9680 37204 9732 37256
rect 3240 37068 3292 37120
rect 5724 37068 5776 37120
rect 6000 37068 6052 37120
rect 8024 37111 8076 37120
rect 8024 37077 8033 37111
rect 8033 37077 8067 37111
rect 8067 37077 8076 37111
rect 8024 37068 8076 37077
rect 9496 37111 9548 37120
rect 9496 37077 9505 37111
rect 9505 37077 9539 37111
rect 9539 37077 9548 37111
rect 9496 37068 9548 37077
rect 10876 37068 10928 37120
rect 11060 37111 11112 37120
rect 11060 37077 11069 37111
rect 11069 37077 11103 37111
rect 11103 37077 11112 37111
rect 11060 37068 11112 37077
rect 14004 37204 14056 37256
rect 14188 37204 14240 37256
rect 15568 37247 15620 37256
rect 13544 37136 13596 37188
rect 15568 37213 15577 37247
rect 15577 37213 15611 37247
rect 15611 37213 15620 37247
rect 15568 37204 15620 37213
rect 17776 37204 17828 37256
rect 17868 37204 17920 37256
rect 21272 37272 21324 37324
rect 23204 37272 23256 37324
rect 19432 37204 19484 37256
rect 20996 37247 21048 37256
rect 14096 37068 14148 37120
rect 14280 37111 14332 37120
rect 14280 37077 14289 37111
rect 14289 37077 14323 37111
rect 14323 37077 14332 37111
rect 14280 37068 14332 37077
rect 14924 37111 14976 37120
rect 14924 37077 14933 37111
rect 14933 37077 14967 37111
rect 14967 37077 14976 37111
rect 14924 37068 14976 37077
rect 15016 37068 15068 37120
rect 18604 37136 18656 37188
rect 20720 37136 20772 37188
rect 15476 37068 15528 37120
rect 17224 37068 17276 37120
rect 17408 37068 17460 37120
rect 18788 37111 18840 37120
rect 18788 37077 18797 37111
rect 18797 37077 18831 37111
rect 18831 37077 18840 37111
rect 18788 37068 18840 37077
rect 19984 37068 20036 37120
rect 20996 37213 21005 37247
rect 21005 37213 21039 37247
rect 21039 37213 21048 37247
rect 20996 37204 21048 37213
rect 22560 37204 22612 37256
rect 23112 37204 23164 37256
rect 23388 37204 23440 37256
rect 25044 37204 25096 37256
rect 26608 37204 26660 37256
rect 27804 37247 27856 37256
rect 20904 37136 20956 37188
rect 21916 37136 21968 37188
rect 25228 37179 25280 37188
rect 25228 37145 25237 37179
rect 25237 37145 25271 37179
rect 25271 37145 25280 37179
rect 25228 37136 25280 37145
rect 25320 37179 25372 37188
rect 25320 37145 25329 37179
rect 25329 37145 25363 37179
rect 25363 37145 25372 37179
rect 27804 37213 27813 37247
rect 27813 37213 27847 37247
rect 27847 37213 27856 37247
rect 27804 37204 27856 37213
rect 28540 37247 28592 37256
rect 28540 37213 28549 37247
rect 28549 37213 28583 37247
rect 28583 37213 28592 37247
rect 30380 37272 30432 37324
rect 30932 37272 30984 37324
rect 32588 37247 32640 37256
rect 28540 37204 28592 37213
rect 25320 37136 25372 37145
rect 23388 37111 23440 37120
rect 23388 37077 23397 37111
rect 23397 37077 23431 37111
rect 23431 37077 23440 37111
rect 23388 37068 23440 37077
rect 24492 37068 24544 37120
rect 28908 37136 28960 37188
rect 32588 37213 32597 37247
rect 32597 37213 32631 37247
rect 32631 37213 32640 37247
rect 32588 37204 32640 37213
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 34796 37204 34848 37256
rect 36084 37204 36136 37256
rect 37372 37204 37424 37256
rect 30472 37179 30524 37188
rect 30472 37145 30481 37179
rect 30481 37145 30515 37179
rect 30515 37145 30524 37179
rect 30472 37136 30524 37145
rect 27712 37068 27764 37120
rect 28632 37111 28684 37120
rect 28632 37077 28641 37111
rect 28641 37077 28675 37111
rect 28675 37077 28684 37111
rect 28632 37068 28684 37077
rect 33140 37068 33192 37120
rect 34520 37068 34572 37120
rect 36360 37111 36412 37120
rect 36360 37077 36369 37111
rect 36369 37077 36403 37111
rect 36403 37077 36412 37111
rect 36360 37068 36412 37077
rect 37648 37111 37700 37120
rect 37648 37077 37657 37111
rect 37657 37077 37691 37111
rect 37691 37077 37700 37111
rect 37648 37068 37700 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 6552 36864 6604 36916
rect 10140 36864 10192 36916
rect 10876 36864 10928 36916
rect 6092 36796 6144 36848
rect 11980 36796 12032 36848
rect 1308 36728 1360 36780
rect 4712 36771 4764 36780
rect 4712 36737 4721 36771
rect 4721 36737 4755 36771
rect 4755 36737 4764 36771
rect 4712 36728 4764 36737
rect 5724 36728 5776 36780
rect 7656 36771 7708 36780
rect 7656 36737 7665 36771
rect 7665 36737 7699 36771
rect 7699 36737 7708 36771
rect 7656 36728 7708 36737
rect 9036 36728 9088 36780
rect 8668 36703 8720 36712
rect 8668 36669 8677 36703
rect 8677 36669 8711 36703
rect 8711 36669 8720 36703
rect 8668 36660 8720 36669
rect 10416 36660 10468 36712
rect 3424 36592 3476 36644
rect 11888 36592 11940 36644
rect 12900 36864 12952 36916
rect 13912 36864 13964 36916
rect 14832 36864 14884 36916
rect 14924 36864 14976 36916
rect 20076 36864 20128 36916
rect 20628 36864 20680 36916
rect 20996 36864 21048 36916
rect 21916 36864 21968 36916
rect 22652 36907 22704 36916
rect 22652 36873 22661 36907
rect 22661 36873 22695 36907
rect 22695 36873 22704 36907
rect 22652 36864 22704 36873
rect 12440 36660 12492 36712
rect 12992 36703 13044 36712
rect 12992 36669 13001 36703
rect 13001 36669 13035 36703
rect 13035 36669 13044 36703
rect 12992 36660 13044 36669
rect 16764 36796 16816 36848
rect 17408 36796 17460 36848
rect 18420 36796 18472 36848
rect 24216 36839 24268 36848
rect 18236 36728 18288 36780
rect 19340 36728 19392 36780
rect 20076 36771 20128 36780
rect 20076 36737 20085 36771
rect 20085 36737 20119 36771
rect 20119 36737 20128 36771
rect 20076 36728 20128 36737
rect 20720 36771 20772 36780
rect 20720 36737 20729 36771
rect 20729 36737 20763 36771
rect 20763 36737 20772 36771
rect 20720 36728 20772 36737
rect 22284 36728 22336 36780
rect 22744 36728 22796 36780
rect 23204 36728 23256 36780
rect 24216 36805 24225 36839
rect 24225 36805 24259 36839
rect 24259 36805 24268 36839
rect 24216 36796 24268 36805
rect 25228 36864 25280 36916
rect 26608 36864 26660 36916
rect 27804 36864 27856 36916
rect 27896 36864 27948 36916
rect 25872 36771 25924 36780
rect 25872 36737 25881 36771
rect 25881 36737 25915 36771
rect 25915 36737 25924 36771
rect 25872 36728 25924 36737
rect 26332 36771 26384 36780
rect 26332 36737 26341 36771
rect 26341 36737 26375 36771
rect 26375 36737 26384 36771
rect 26332 36728 26384 36737
rect 1860 36524 1912 36576
rect 2688 36567 2740 36576
rect 2688 36533 2697 36567
rect 2697 36533 2731 36567
rect 2731 36533 2740 36567
rect 2688 36524 2740 36533
rect 6460 36524 6512 36576
rect 7748 36567 7800 36576
rect 7748 36533 7757 36567
rect 7757 36533 7791 36567
rect 7791 36533 7800 36567
rect 7748 36524 7800 36533
rect 9128 36567 9180 36576
rect 9128 36533 9137 36567
rect 9137 36533 9171 36567
rect 9171 36533 9180 36567
rect 9128 36524 9180 36533
rect 10324 36567 10376 36576
rect 10324 36533 10333 36567
rect 10333 36533 10367 36567
rect 10367 36533 10376 36567
rect 10324 36524 10376 36533
rect 16764 36660 16816 36712
rect 16580 36592 16632 36644
rect 16672 36592 16724 36644
rect 17224 36660 17276 36712
rect 19248 36660 19300 36712
rect 20536 36660 20588 36712
rect 23940 36660 23992 36712
rect 24032 36703 24084 36712
rect 24032 36669 24041 36703
rect 24041 36669 24075 36703
rect 24075 36669 24084 36703
rect 26608 36728 26660 36780
rect 27252 36728 27304 36780
rect 27436 36796 27488 36848
rect 30288 36796 30340 36848
rect 32220 36864 32272 36916
rect 38108 36839 38160 36848
rect 38108 36805 38117 36839
rect 38117 36805 38151 36839
rect 38151 36805 38160 36839
rect 38108 36796 38160 36805
rect 33048 36771 33100 36780
rect 24032 36660 24084 36669
rect 18144 36592 18196 36644
rect 22100 36592 22152 36644
rect 22192 36592 22244 36644
rect 25872 36592 25924 36644
rect 27712 36660 27764 36712
rect 27804 36660 27856 36712
rect 28080 36703 28132 36712
rect 28080 36669 28089 36703
rect 28089 36669 28123 36703
rect 28123 36669 28132 36703
rect 28080 36660 28132 36669
rect 29000 36703 29052 36712
rect 29000 36669 29009 36703
rect 29009 36669 29043 36703
rect 29043 36669 29052 36703
rect 29000 36660 29052 36669
rect 29092 36660 29144 36712
rect 30380 36660 30432 36712
rect 15016 36567 15068 36576
rect 15016 36533 15025 36567
rect 15025 36533 15059 36567
rect 15059 36533 15068 36567
rect 15016 36524 15068 36533
rect 16948 36524 17000 36576
rect 17132 36524 17184 36576
rect 17868 36524 17920 36576
rect 20260 36524 20312 36576
rect 21916 36524 21968 36576
rect 22008 36524 22060 36576
rect 26700 36592 26752 36644
rect 33048 36737 33057 36771
rect 33057 36737 33091 36771
rect 33091 36737 33100 36771
rect 33048 36728 33100 36737
rect 35440 36728 35492 36780
rect 39304 36728 39356 36780
rect 32680 36592 32732 36644
rect 26424 36567 26476 36576
rect 26424 36533 26433 36567
rect 26433 36533 26467 36567
rect 26467 36533 26476 36567
rect 26424 36524 26476 36533
rect 27344 36524 27396 36576
rect 28632 36524 28684 36576
rect 32496 36567 32548 36576
rect 32496 36533 32505 36567
rect 32505 36533 32539 36567
rect 32539 36533 32548 36567
rect 32496 36524 32548 36533
rect 36728 36567 36780 36576
rect 36728 36533 36737 36567
rect 36737 36533 36771 36567
rect 36771 36533 36780 36567
rect 36728 36524 36780 36533
rect 37280 36524 37332 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4712 36320 4764 36372
rect 8668 36320 8720 36372
rect 7656 36252 7708 36304
rect 8116 36252 8168 36304
rect 14004 36320 14056 36372
rect 18420 36320 18472 36372
rect 18788 36320 18840 36372
rect 20536 36320 20588 36372
rect 20812 36320 20864 36372
rect 21640 36320 21692 36372
rect 22652 36320 22704 36372
rect 33048 36320 33100 36372
rect 37188 36320 37240 36372
rect 9128 36252 9180 36304
rect 6460 36227 6512 36236
rect 6460 36193 6469 36227
rect 6469 36193 6503 36227
rect 6503 36193 6512 36227
rect 6460 36184 6512 36193
rect 20 36116 72 36168
rect 2872 36116 2924 36168
rect 9588 36184 9640 36236
rect 10232 36184 10284 36236
rect 10416 36227 10468 36236
rect 10416 36193 10425 36227
rect 10425 36193 10459 36227
rect 10459 36193 10468 36227
rect 10416 36184 10468 36193
rect 6552 36091 6604 36100
rect 6552 36057 6561 36091
rect 6561 36057 6595 36091
rect 6595 36057 6604 36091
rect 6552 36048 6604 36057
rect 6828 36048 6880 36100
rect 10876 36116 10928 36168
rect 12900 36252 12952 36304
rect 12992 36252 13044 36304
rect 16396 36252 16448 36304
rect 18236 36252 18288 36304
rect 11980 36184 12032 36236
rect 9128 36048 9180 36100
rect 9772 36048 9824 36100
rect 9956 36048 10008 36100
rect 11888 36116 11940 36168
rect 13544 36159 13596 36168
rect 13544 36125 13553 36159
rect 13553 36125 13587 36159
rect 13587 36125 13596 36159
rect 13544 36116 13596 36125
rect 15568 36184 15620 36236
rect 20260 36184 20312 36236
rect 21088 36184 21140 36236
rect 16764 36159 16816 36168
rect 16764 36125 16773 36159
rect 16773 36125 16807 36159
rect 16807 36125 16816 36159
rect 16764 36116 16816 36125
rect 18144 36116 18196 36168
rect 18328 36116 18380 36168
rect 14648 36091 14700 36100
rect 14648 36057 14657 36091
rect 14657 36057 14691 36091
rect 14691 36057 14700 36091
rect 14648 36048 14700 36057
rect 15568 36048 15620 36100
rect 11060 35980 11112 36032
rect 11520 36023 11572 36032
rect 11520 35989 11529 36023
rect 11529 35989 11563 36023
rect 11563 35989 11572 36023
rect 11520 35980 11572 35989
rect 11612 35980 11664 36032
rect 14280 35980 14332 36032
rect 19432 36048 19484 36100
rect 19708 36159 19760 36168
rect 19708 36125 19717 36159
rect 19717 36125 19751 36159
rect 19751 36125 19760 36159
rect 19708 36116 19760 36125
rect 20076 36116 20128 36168
rect 20168 36048 20220 36100
rect 20536 36091 20588 36100
rect 20536 36057 20545 36091
rect 20545 36057 20579 36091
rect 20579 36057 20588 36091
rect 20536 36048 20588 36057
rect 20904 36048 20956 36100
rect 26700 36252 26752 36304
rect 27436 36252 27488 36304
rect 18512 36023 18564 36032
rect 18512 35989 18521 36023
rect 18521 35989 18555 36023
rect 18555 35989 18564 36023
rect 18512 35980 18564 35989
rect 18696 35980 18748 36032
rect 19708 35980 19760 36032
rect 22100 35980 22152 36032
rect 23388 36116 23440 36168
rect 23480 36116 23532 36168
rect 25136 36184 25188 36236
rect 27252 36184 27304 36236
rect 24032 36048 24084 36100
rect 31852 36159 31904 36168
rect 31852 36125 31861 36159
rect 31861 36125 31895 36159
rect 31895 36125 31904 36159
rect 31852 36116 31904 36125
rect 32312 36159 32364 36168
rect 32312 36125 32321 36159
rect 32321 36125 32355 36159
rect 32355 36125 32364 36159
rect 32312 36116 32364 36125
rect 38660 36184 38712 36236
rect 24676 36091 24728 36100
rect 24676 36057 24685 36091
rect 24685 36057 24719 36091
rect 24719 36057 24728 36091
rect 24676 36048 24728 36057
rect 24768 36091 24820 36100
rect 24768 36057 24777 36091
rect 24777 36057 24811 36091
rect 24811 36057 24820 36091
rect 24768 36048 24820 36057
rect 25504 36048 25556 36100
rect 25964 36091 26016 36100
rect 25964 36057 25973 36091
rect 25973 36057 26007 36091
rect 26007 36057 26016 36091
rect 25964 36048 26016 36057
rect 26240 36048 26292 36100
rect 27068 36048 27120 36100
rect 28080 36091 28132 36100
rect 28080 36057 28089 36091
rect 28089 36057 28123 36091
rect 28123 36057 28132 36091
rect 28080 36048 28132 36057
rect 29000 36048 29052 36100
rect 30840 36048 30892 36100
rect 31024 36048 31076 36100
rect 37372 36116 37424 36168
rect 38384 36048 38436 36100
rect 30380 35980 30432 36032
rect 34520 35980 34572 36032
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 10876 35819 10928 35828
rect 10876 35785 10885 35819
rect 10885 35785 10919 35819
rect 10919 35785 10928 35819
rect 10876 35776 10928 35785
rect 9312 35751 9364 35760
rect 9312 35717 9321 35751
rect 9321 35717 9355 35751
rect 9355 35717 9364 35751
rect 9312 35708 9364 35717
rect 16948 35776 17000 35828
rect 20720 35776 20772 35828
rect 20904 35776 20956 35828
rect 21180 35776 21232 35828
rect 22100 35776 22152 35828
rect 24676 35776 24728 35828
rect 25964 35776 26016 35828
rect 27620 35776 27672 35828
rect 1676 35683 1728 35692
rect 1676 35649 1685 35683
rect 1685 35649 1719 35683
rect 1719 35649 1728 35683
rect 1676 35640 1728 35649
rect 3424 35683 3476 35692
rect 3424 35649 3433 35683
rect 3433 35649 3467 35683
rect 3467 35649 3476 35683
rect 3424 35640 3476 35649
rect 3608 35640 3660 35692
rect 4068 35572 4120 35624
rect 21548 35708 21600 35760
rect 11520 35640 11572 35692
rect 12440 35615 12492 35624
rect 12440 35581 12449 35615
rect 12449 35581 12483 35615
rect 12483 35581 12492 35615
rect 12440 35572 12492 35581
rect 12808 35572 12860 35624
rect 14648 35572 14700 35624
rect 17224 35572 17276 35624
rect 17868 35572 17920 35624
rect 19984 35640 20036 35692
rect 20352 35640 20404 35692
rect 20720 35683 20772 35692
rect 20720 35649 20729 35683
rect 20729 35649 20763 35683
rect 20763 35649 20772 35683
rect 20720 35640 20772 35649
rect 22284 35708 22336 35760
rect 22468 35708 22520 35760
rect 20168 35572 20220 35624
rect 22192 35683 22244 35692
rect 22192 35649 22201 35683
rect 22201 35649 22235 35683
rect 22235 35649 22244 35683
rect 22192 35640 22244 35649
rect 22376 35640 22428 35692
rect 23480 35640 23532 35692
rect 21272 35572 21324 35624
rect 22100 35572 22152 35624
rect 26424 35708 26476 35760
rect 24584 35683 24636 35692
rect 24584 35649 24593 35683
rect 24593 35649 24627 35683
rect 24627 35649 24636 35683
rect 24584 35640 24636 35649
rect 25412 35640 25464 35692
rect 25688 35640 25740 35692
rect 27712 35708 27764 35760
rect 27988 35751 28040 35760
rect 27988 35717 27997 35751
rect 27997 35717 28031 35751
rect 28031 35717 28040 35751
rect 27988 35708 28040 35717
rect 29828 35708 29880 35760
rect 27160 35683 27212 35692
rect 27160 35649 27169 35683
rect 27169 35649 27203 35683
rect 27203 35649 27212 35683
rect 30840 35776 30892 35828
rect 27160 35640 27212 35649
rect 30564 35640 30616 35692
rect 26884 35572 26936 35624
rect 1492 35436 1544 35488
rect 2596 35436 2648 35488
rect 3976 35436 4028 35488
rect 7840 35436 7892 35488
rect 12256 35436 12308 35488
rect 12532 35436 12584 35488
rect 14188 35479 14240 35488
rect 14188 35445 14197 35479
rect 14197 35445 14231 35479
rect 14231 35445 14240 35479
rect 18420 35504 18472 35556
rect 14188 35436 14240 35445
rect 18512 35436 18564 35488
rect 20536 35504 20588 35556
rect 20996 35436 21048 35488
rect 21180 35436 21232 35488
rect 22468 35504 22520 35556
rect 28172 35615 28224 35624
rect 28172 35581 28181 35615
rect 28181 35581 28215 35615
rect 28215 35581 28224 35615
rect 28172 35572 28224 35581
rect 28264 35572 28316 35624
rect 37464 35615 37516 35624
rect 27436 35504 27488 35556
rect 22284 35436 22336 35488
rect 27160 35436 27212 35488
rect 27896 35436 27948 35488
rect 30012 35504 30064 35556
rect 31852 35504 31904 35556
rect 29092 35436 29144 35488
rect 29736 35436 29788 35488
rect 37464 35581 37473 35615
rect 37473 35581 37507 35615
rect 37507 35581 37516 35615
rect 37464 35572 37516 35581
rect 37740 35615 37792 35624
rect 37740 35581 37749 35615
rect 37749 35581 37783 35615
rect 37783 35581 37792 35615
rect 37740 35572 37792 35581
rect 32036 35436 32088 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3148 35232 3200 35284
rect 3608 35232 3660 35284
rect 4068 35275 4120 35284
rect 4068 35241 4077 35275
rect 4077 35241 4111 35275
rect 4111 35241 4120 35275
rect 4068 35232 4120 35241
rect 4896 35232 4948 35284
rect 9588 35232 9640 35284
rect 9772 35232 9824 35284
rect 12532 35232 12584 35284
rect 12256 35164 12308 35216
rect 16396 35207 16448 35216
rect 16396 35173 16405 35207
rect 16405 35173 16439 35207
rect 16439 35173 16448 35207
rect 16396 35164 16448 35173
rect 5356 35096 5408 35148
rect 8208 35096 8260 35148
rect 12440 35096 12492 35148
rect 13176 35096 13228 35148
rect 13360 35139 13412 35148
rect 13360 35105 13369 35139
rect 13369 35105 13403 35139
rect 13403 35105 13412 35139
rect 13360 35096 13412 35105
rect 14648 35139 14700 35148
rect 14648 35105 14657 35139
rect 14657 35105 14691 35139
rect 14691 35105 14700 35139
rect 14648 35096 14700 35105
rect 16488 35096 16540 35148
rect 17132 35139 17184 35148
rect 17132 35105 17141 35139
rect 17141 35105 17175 35139
rect 17175 35105 17184 35139
rect 17132 35096 17184 35105
rect 17500 35096 17552 35148
rect 19340 35164 19392 35216
rect 19984 35164 20036 35216
rect 21824 35164 21876 35216
rect 24768 35232 24820 35284
rect 26516 35232 26568 35284
rect 29920 35232 29972 35284
rect 30472 35275 30524 35284
rect 30472 35241 30481 35275
rect 30481 35241 30515 35275
rect 30515 35241 30524 35275
rect 30472 35232 30524 35241
rect 32312 35232 32364 35284
rect 28080 35164 28132 35216
rect 28356 35164 28408 35216
rect 30012 35164 30064 35216
rect 3332 35028 3384 35080
rect 10508 35071 10560 35080
rect 2596 34960 2648 35012
rect 10508 35037 10517 35071
rect 10517 35037 10551 35071
rect 10551 35037 10560 35071
rect 10508 35028 10560 35037
rect 13268 35071 13320 35080
rect 13268 35037 13277 35071
rect 13277 35037 13311 35071
rect 13311 35037 13320 35071
rect 13268 35028 13320 35037
rect 16856 35071 16908 35080
rect 16856 35037 16865 35071
rect 16865 35037 16899 35071
rect 16899 35037 16908 35071
rect 16856 35028 16908 35037
rect 26240 35139 26292 35148
rect 26240 35105 26249 35139
rect 26249 35105 26283 35139
rect 26283 35105 26292 35139
rect 26240 35096 26292 35105
rect 27436 35096 27488 35148
rect 19432 35071 19484 35080
rect 19432 35037 19441 35071
rect 19441 35037 19475 35071
rect 19475 35037 19484 35071
rect 19432 35028 19484 35037
rect 20168 35071 20220 35080
rect 20168 35037 20177 35071
rect 20177 35037 20211 35071
rect 20211 35037 20220 35071
rect 20168 35028 20220 35037
rect 20260 35028 20312 35080
rect 20720 35028 20772 35080
rect 21456 35071 21508 35080
rect 21456 35037 21465 35071
rect 21465 35037 21499 35071
rect 21499 35037 21508 35071
rect 21456 35028 21508 35037
rect 22376 35028 22428 35080
rect 2688 34892 2740 34944
rect 4620 34892 4672 34944
rect 14832 34960 14884 35012
rect 7748 34935 7800 34944
rect 7748 34901 7757 34935
rect 7757 34901 7791 34935
rect 7791 34901 7800 34935
rect 7748 34892 7800 34901
rect 12624 34892 12676 34944
rect 12716 34892 12768 34944
rect 16948 34892 17000 34944
rect 18604 34935 18656 34944
rect 18604 34901 18613 34935
rect 18613 34901 18647 34935
rect 18647 34901 18656 34935
rect 18604 34892 18656 34901
rect 20168 34892 20220 34944
rect 20444 34892 20496 34944
rect 20720 34892 20772 34944
rect 20996 34892 21048 34944
rect 21824 34960 21876 35012
rect 23480 35028 23532 35080
rect 23664 35071 23716 35080
rect 23664 35037 23673 35071
rect 23673 35037 23707 35071
rect 23707 35037 23716 35071
rect 23664 35028 23716 35037
rect 25596 35028 25648 35080
rect 28172 35139 28224 35148
rect 28172 35105 28181 35139
rect 28181 35105 28215 35139
rect 28215 35105 28224 35139
rect 28172 35096 28224 35105
rect 28908 35071 28960 35080
rect 22836 34935 22888 34944
rect 22836 34901 22845 34935
rect 22845 34901 22879 34935
rect 22879 34901 22888 34935
rect 22836 34892 22888 34901
rect 22928 34892 22980 34944
rect 26884 34960 26936 35012
rect 28908 35037 28917 35071
rect 28917 35037 28951 35071
rect 28951 35037 28960 35071
rect 28908 35028 28960 35037
rect 29920 35071 29972 35080
rect 29920 35037 29929 35071
rect 29929 35037 29963 35071
rect 29963 35037 29972 35071
rect 29920 35028 29972 35037
rect 30012 35028 30064 35080
rect 27160 34960 27212 35012
rect 27528 34960 27580 35012
rect 27896 35003 27948 35012
rect 27896 34969 27905 35003
rect 27905 34969 27939 35003
rect 27939 34969 27948 35003
rect 27896 34960 27948 34969
rect 27988 34960 28040 35012
rect 31024 34960 31076 35012
rect 28540 34892 28592 34944
rect 29000 34935 29052 34944
rect 29000 34901 29009 34935
rect 29009 34901 29043 34935
rect 29043 34901 29052 34935
rect 29000 34892 29052 34901
rect 29276 34892 29328 34944
rect 38016 34935 38068 34944
rect 38016 34901 38025 34935
rect 38025 34901 38059 34935
rect 38059 34901 38068 34935
rect 38016 34892 38068 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 3332 34688 3384 34740
rect 5356 34731 5408 34740
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 3976 34620 4028 34672
rect 2872 34552 2924 34604
rect 5356 34697 5365 34731
rect 5365 34697 5399 34731
rect 5399 34697 5408 34731
rect 5356 34688 5408 34697
rect 6552 34688 6604 34740
rect 10508 34688 10560 34740
rect 15568 34731 15620 34740
rect 5724 34552 5776 34604
rect 6276 34552 6328 34604
rect 2688 34484 2740 34536
rect 7748 34552 7800 34604
rect 9588 34552 9640 34604
rect 13268 34620 13320 34672
rect 14372 34620 14424 34672
rect 15568 34697 15577 34731
rect 15577 34697 15611 34731
rect 15611 34697 15620 34731
rect 15568 34688 15620 34697
rect 16672 34688 16724 34740
rect 17868 34688 17920 34740
rect 17960 34688 18012 34740
rect 19984 34688 20036 34740
rect 17408 34620 17460 34672
rect 22100 34688 22152 34740
rect 23940 34688 23992 34740
rect 25044 34688 25096 34740
rect 28540 34731 28592 34740
rect 20536 34620 20588 34672
rect 22468 34663 22520 34672
rect 22468 34629 22477 34663
rect 22477 34629 22511 34663
rect 22511 34629 22520 34663
rect 22468 34620 22520 34629
rect 12440 34552 12492 34604
rect 12624 34595 12676 34604
rect 12624 34561 12633 34595
rect 12633 34561 12667 34595
rect 12667 34561 12676 34595
rect 12624 34552 12676 34561
rect 12716 34595 12768 34604
rect 12716 34561 12725 34595
rect 12725 34561 12759 34595
rect 12759 34561 12768 34595
rect 22376 34595 22428 34604
rect 12716 34552 12768 34561
rect 22376 34561 22385 34595
rect 22385 34561 22419 34595
rect 22419 34561 22428 34595
rect 22376 34552 22428 34561
rect 6276 34416 6328 34468
rect 16856 34527 16908 34536
rect 13176 34348 13228 34400
rect 16856 34493 16865 34527
rect 16865 34493 16899 34527
rect 16899 34493 16908 34527
rect 16856 34484 16908 34493
rect 17224 34484 17276 34536
rect 16304 34416 16356 34468
rect 16488 34416 16540 34468
rect 18144 34416 18196 34468
rect 20812 34527 20864 34536
rect 20812 34493 20821 34527
rect 20821 34493 20855 34527
rect 20855 34493 20864 34527
rect 21180 34527 21232 34536
rect 20812 34484 20864 34493
rect 21180 34493 21189 34527
rect 21189 34493 21223 34527
rect 21223 34493 21232 34527
rect 21180 34484 21232 34493
rect 21548 34484 21600 34536
rect 23020 34595 23072 34604
rect 23020 34561 23029 34595
rect 23029 34561 23063 34595
rect 23063 34561 23072 34595
rect 23020 34552 23072 34561
rect 23388 34552 23440 34604
rect 23848 34552 23900 34604
rect 25596 34595 25648 34604
rect 23112 34527 23164 34536
rect 23112 34493 23121 34527
rect 23121 34493 23155 34527
rect 23155 34493 23164 34527
rect 23112 34484 23164 34493
rect 23480 34484 23532 34536
rect 23756 34527 23808 34536
rect 23756 34493 23765 34527
rect 23765 34493 23799 34527
rect 23799 34493 23808 34527
rect 23756 34484 23808 34493
rect 25596 34561 25605 34595
rect 25605 34561 25639 34595
rect 25639 34561 25648 34595
rect 25596 34552 25648 34561
rect 26424 34552 26476 34604
rect 14648 34348 14700 34400
rect 15844 34348 15896 34400
rect 16672 34348 16724 34400
rect 16948 34348 17000 34400
rect 18512 34348 18564 34400
rect 22284 34416 22336 34468
rect 23204 34416 23256 34468
rect 23572 34416 23624 34468
rect 25228 34484 25280 34536
rect 25320 34484 25372 34536
rect 26884 34484 26936 34536
rect 27804 34595 27856 34604
rect 27804 34561 27813 34595
rect 27813 34561 27847 34595
rect 27847 34561 27856 34595
rect 27804 34552 27856 34561
rect 28540 34697 28549 34731
rect 28549 34697 28583 34731
rect 28583 34697 28592 34731
rect 28540 34688 28592 34697
rect 29828 34731 29880 34740
rect 29828 34697 29837 34731
rect 29837 34697 29871 34731
rect 29871 34697 29880 34731
rect 29828 34688 29880 34697
rect 30380 34688 30432 34740
rect 28080 34620 28132 34672
rect 28448 34595 28500 34604
rect 28448 34561 28457 34595
rect 28457 34561 28491 34595
rect 28491 34561 28500 34595
rect 28448 34552 28500 34561
rect 27436 34484 27488 34536
rect 36728 34552 36780 34604
rect 37832 34552 37884 34604
rect 22560 34348 22612 34400
rect 24400 34391 24452 34400
rect 24400 34357 24409 34391
rect 24409 34357 24443 34391
rect 24443 34357 24452 34391
rect 24400 34348 24452 34357
rect 26700 34348 26752 34400
rect 27528 34348 27580 34400
rect 30012 34484 30064 34536
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 4620 34144 4672 34196
rect 8208 34144 8260 34196
rect 13728 34144 13780 34196
rect 8944 34008 8996 34060
rect 11060 34051 11112 34060
rect 11060 34017 11069 34051
rect 11069 34017 11103 34051
rect 11103 34017 11112 34051
rect 11060 34008 11112 34017
rect 13268 34008 13320 34060
rect 15844 34076 15896 34128
rect 14648 34008 14700 34060
rect 16856 34008 16908 34060
rect 16948 34008 17000 34060
rect 18512 34076 18564 34128
rect 18604 34076 18656 34128
rect 27252 34144 27304 34196
rect 23572 34119 23624 34128
rect 23572 34085 23581 34119
rect 23581 34085 23615 34119
rect 23615 34085 23624 34119
rect 23572 34076 23624 34085
rect 17408 34008 17460 34060
rect 18420 34008 18472 34060
rect 23940 34008 23992 34060
rect 25504 34076 25556 34128
rect 24952 34051 25004 34060
rect 24952 34017 24961 34051
rect 24961 34017 24995 34051
rect 24995 34017 25004 34051
rect 24952 34008 25004 34017
rect 25412 34008 25464 34060
rect 27436 34008 27488 34060
rect 3424 33940 3476 33992
rect 8116 33940 8168 33992
rect 15384 33940 15436 33992
rect 19156 33940 19208 33992
rect 20260 33940 20312 33992
rect 22376 33940 22428 33992
rect 24492 33940 24544 33992
rect 25596 33940 25648 33992
rect 28172 34076 28224 34128
rect 29092 34144 29144 34196
rect 37832 34187 37884 34196
rect 37832 34153 37841 34187
rect 37841 34153 37875 34187
rect 37875 34153 37884 34187
rect 37832 34144 37884 34153
rect 29184 34076 29236 34128
rect 29000 34008 29052 34060
rect 28540 33940 28592 33992
rect 33048 33940 33100 33992
rect 38016 33983 38068 33992
rect 38016 33949 38025 33983
rect 38025 33949 38059 33983
rect 38059 33949 38068 33983
rect 38016 33940 38068 33949
rect 10324 33872 10376 33924
rect 10600 33915 10652 33924
rect 10600 33881 10609 33915
rect 10609 33881 10643 33915
rect 10643 33881 10652 33915
rect 10600 33872 10652 33881
rect 12532 33872 12584 33924
rect 11428 33804 11480 33856
rect 11704 33804 11756 33856
rect 16028 33804 16080 33856
rect 16212 33915 16264 33924
rect 16212 33881 16221 33915
rect 16221 33881 16255 33915
rect 16255 33881 16264 33915
rect 16212 33872 16264 33881
rect 22836 33872 22888 33924
rect 17684 33847 17736 33856
rect 17684 33813 17693 33847
rect 17693 33813 17727 33847
rect 17727 33813 17736 33847
rect 17684 33804 17736 33813
rect 17868 33804 17920 33856
rect 21180 33804 21232 33856
rect 25412 33804 25464 33856
rect 25872 33847 25924 33856
rect 25872 33813 25881 33847
rect 25881 33813 25915 33847
rect 25915 33813 25924 33847
rect 25872 33804 25924 33813
rect 26700 33915 26752 33924
rect 26700 33881 26709 33915
rect 26709 33881 26743 33915
rect 26743 33881 26752 33915
rect 26700 33872 26752 33881
rect 27804 33872 27856 33924
rect 27988 33804 28040 33856
rect 29736 33847 29788 33856
rect 29736 33813 29745 33847
rect 29745 33813 29779 33847
rect 29779 33813 29788 33847
rect 29736 33804 29788 33813
rect 29828 33804 29880 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4804 33600 4856 33652
rect 10600 33600 10652 33652
rect 15844 33600 15896 33652
rect 16212 33600 16264 33652
rect 17408 33600 17460 33652
rect 17500 33600 17552 33652
rect 20904 33600 20956 33652
rect 21088 33643 21140 33652
rect 21088 33609 21097 33643
rect 21097 33609 21131 33643
rect 21131 33609 21140 33643
rect 21088 33600 21140 33609
rect 21180 33600 21232 33652
rect 24492 33600 24544 33652
rect 2688 33532 2740 33584
rect 2780 33532 2832 33584
rect 7840 33532 7892 33584
rect 13728 33532 13780 33584
rect 17132 33532 17184 33584
rect 6184 33464 6236 33516
rect 11704 33507 11756 33516
rect 3148 33396 3200 33448
rect 5540 33396 5592 33448
rect 7472 33439 7524 33448
rect 7472 33405 7481 33439
rect 7481 33405 7515 33439
rect 7515 33405 7524 33439
rect 7472 33396 7524 33405
rect 8208 33396 8260 33448
rect 11704 33473 11713 33507
rect 11713 33473 11747 33507
rect 11747 33473 11756 33507
rect 11704 33464 11756 33473
rect 13176 33507 13228 33516
rect 13176 33473 13185 33507
rect 13185 33473 13219 33507
rect 13219 33473 13228 33507
rect 13176 33464 13228 33473
rect 20996 33507 21048 33516
rect 9404 33396 9456 33448
rect 14004 33396 14056 33448
rect 16856 33396 16908 33448
rect 1768 33371 1820 33380
rect 1768 33337 1777 33371
rect 1777 33337 1811 33371
rect 1811 33337 1820 33371
rect 1768 33328 1820 33337
rect 15108 33328 15160 33380
rect 17868 33396 17920 33448
rect 20996 33473 21005 33507
rect 21005 33473 21039 33507
rect 21039 33473 21048 33507
rect 20996 33464 21048 33473
rect 23940 33532 23992 33584
rect 24308 33532 24360 33584
rect 24400 33532 24452 33584
rect 29736 33600 29788 33652
rect 29000 33575 29052 33584
rect 29000 33541 29009 33575
rect 29009 33541 29043 33575
rect 29043 33541 29052 33575
rect 29000 33532 29052 33541
rect 22744 33464 22796 33516
rect 23112 33464 23164 33516
rect 23480 33464 23532 33516
rect 24032 33507 24084 33516
rect 24032 33473 24041 33507
rect 24041 33473 24075 33507
rect 24075 33473 24084 33507
rect 24032 33464 24084 33473
rect 22928 33396 22980 33448
rect 25044 33396 25096 33448
rect 25964 33439 26016 33448
rect 25964 33405 25973 33439
rect 25973 33405 26007 33439
rect 26007 33405 26016 33439
rect 25964 33396 26016 33405
rect 26792 33464 26844 33516
rect 27252 33464 27304 33516
rect 27896 33396 27948 33448
rect 29184 33439 29236 33448
rect 29184 33405 29193 33439
rect 29193 33405 29227 33439
rect 29227 33405 29236 33439
rect 29184 33396 29236 33405
rect 4620 33260 4672 33312
rect 4712 33260 4764 33312
rect 15660 33260 15712 33312
rect 28080 33328 28132 33380
rect 18512 33260 18564 33312
rect 22560 33260 22612 33312
rect 22652 33260 22704 33312
rect 24860 33260 24912 33312
rect 27620 33260 27672 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4804 33056 4856 33108
rect 14372 33099 14424 33108
rect 14372 33065 14381 33099
rect 14381 33065 14415 33099
rect 14415 33065 14424 33099
rect 14372 33056 14424 33065
rect 6828 32988 6880 33040
rect 14004 32988 14056 33040
rect 18972 33056 19024 33108
rect 19156 33056 19208 33108
rect 23940 33099 23992 33108
rect 23940 33065 23949 33099
rect 23949 33065 23983 33099
rect 23983 33065 23992 33099
rect 23940 33056 23992 33065
rect 2596 32920 2648 32972
rect 5540 32963 5592 32972
rect 5540 32929 5549 32963
rect 5549 32929 5583 32963
rect 5583 32929 5592 32963
rect 5540 32920 5592 32929
rect 14188 32920 14240 32972
rect 4712 32895 4764 32904
rect 4712 32861 4721 32895
rect 4721 32861 4755 32895
rect 4755 32861 4764 32895
rect 4712 32852 4764 32861
rect 6184 32895 6236 32904
rect 6184 32861 6193 32895
rect 6193 32861 6227 32895
rect 6227 32861 6236 32895
rect 6828 32895 6880 32904
rect 6184 32852 6236 32861
rect 6828 32861 6837 32895
rect 6837 32861 6871 32895
rect 6871 32861 6880 32895
rect 6828 32852 6880 32861
rect 2872 32784 2924 32836
rect 8944 32852 8996 32904
rect 11428 32852 11480 32904
rect 4896 32716 4948 32768
rect 10232 32784 10284 32836
rect 11612 32784 11664 32836
rect 16764 32920 16816 32972
rect 18880 32988 18932 33040
rect 19432 32988 19484 33040
rect 20628 32988 20680 33040
rect 21548 32988 21600 33040
rect 23204 32988 23256 33040
rect 27436 33056 27488 33108
rect 16856 32895 16908 32904
rect 16856 32861 16865 32895
rect 16865 32861 16899 32895
rect 16899 32861 16908 32895
rect 16856 32852 16908 32861
rect 18696 32852 18748 32904
rect 6920 32716 6972 32768
rect 7564 32716 7616 32768
rect 15384 32784 15436 32836
rect 15936 32827 15988 32836
rect 15936 32793 15945 32827
rect 15945 32793 15979 32827
rect 15979 32793 15988 32827
rect 15936 32784 15988 32793
rect 16580 32784 16632 32836
rect 17040 32784 17092 32836
rect 19616 32920 19668 32972
rect 18880 32895 18932 32904
rect 18880 32861 18889 32895
rect 18889 32861 18923 32895
rect 18923 32861 18932 32895
rect 18880 32852 18932 32861
rect 19432 32852 19484 32904
rect 20536 32852 20588 32904
rect 22376 32852 22428 32904
rect 22928 32852 22980 32904
rect 23112 32852 23164 32904
rect 24124 32988 24176 33040
rect 24308 32920 24360 32972
rect 25136 32963 25188 32972
rect 25136 32929 25145 32963
rect 25145 32929 25179 32963
rect 25179 32929 25188 32963
rect 25136 32920 25188 32929
rect 26976 32920 27028 32972
rect 13084 32716 13136 32768
rect 15108 32716 15160 32768
rect 15292 32716 15344 32768
rect 20260 32784 20312 32836
rect 21088 32827 21140 32836
rect 21088 32793 21097 32827
rect 21097 32793 21131 32827
rect 21131 32793 21140 32827
rect 21088 32784 21140 32793
rect 21180 32827 21232 32836
rect 21180 32793 21189 32827
rect 21189 32793 21223 32827
rect 21223 32793 21232 32827
rect 22100 32827 22152 32836
rect 21180 32784 21232 32793
rect 22100 32793 22109 32827
rect 22109 32793 22143 32827
rect 22143 32793 22152 32827
rect 22100 32784 22152 32793
rect 22008 32716 22060 32768
rect 22192 32716 22244 32768
rect 23664 32716 23716 32768
rect 24492 32716 24544 32768
rect 25412 32784 25464 32836
rect 28356 32827 28408 32836
rect 24952 32716 25004 32768
rect 25504 32716 25556 32768
rect 27620 32716 27672 32768
rect 28356 32793 28365 32827
rect 28365 32793 28399 32827
rect 28399 32793 28408 32827
rect 28356 32784 28408 32793
rect 29828 32784 29880 32836
rect 38108 32827 38160 32836
rect 38108 32793 38117 32827
rect 38117 32793 38151 32827
rect 38151 32793 38160 32827
rect 38108 32784 38160 32793
rect 37832 32716 37884 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 7564 32512 7616 32564
rect 7472 32487 7524 32496
rect 7472 32453 7481 32487
rect 7481 32453 7515 32487
rect 7515 32453 7524 32487
rect 7472 32444 7524 32453
rect 13084 32444 13136 32496
rect 2044 32376 2096 32428
rect 6552 32308 6604 32360
rect 1768 32215 1820 32224
rect 1768 32181 1777 32215
rect 1777 32181 1811 32215
rect 1811 32181 1820 32215
rect 1768 32172 1820 32181
rect 5632 32172 5684 32224
rect 8300 32376 8352 32428
rect 8944 32419 8996 32428
rect 8944 32385 8953 32419
rect 8953 32385 8987 32419
rect 8987 32385 8996 32419
rect 8944 32376 8996 32385
rect 15936 32512 15988 32564
rect 13544 32487 13596 32496
rect 13544 32453 13553 32487
rect 13553 32453 13587 32487
rect 13587 32453 13596 32487
rect 13544 32444 13596 32453
rect 15292 32487 15344 32496
rect 15292 32453 15301 32487
rect 15301 32453 15335 32487
rect 15335 32453 15344 32487
rect 15292 32444 15344 32453
rect 15660 32376 15712 32428
rect 18880 32512 18932 32564
rect 18972 32512 19024 32564
rect 26332 32555 26384 32564
rect 19248 32444 19300 32496
rect 19984 32444 20036 32496
rect 26332 32521 26341 32555
rect 26341 32521 26375 32555
rect 26375 32521 26384 32555
rect 26332 32512 26384 32521
rect 27804 32512 27856 32564
rect 29000 32512 29052 32564
rect 33048 32512 33100 32564
rect 22744 32444 22796 32496
rect 23296 32487 23348 32496
rect 23296 32453 23305 32487
rect 23305 32453 23339 32487
rect 23339 32453 23348 32487
rect 23296 32444 23348 32453
rect 24860 32487 24912 32496
rect 24860 32453 24862 32487
rect 24862 32453 24896 32487
rect 24896 32453 24912 32487
rect 24860 32444 24912 32453
rect 16764 32376 16816 32428
rect 18512 32376 18564 32428
rect 18696 32240 18748 32292
rect 18972 32308 19024 32360
rect 20260 32376 20312 32428
rect 20536 32376 20588 32428
rect 21456 32376 21508 32428
rect 21732 32376 21784 32428
rect 21916 32376 21968 32428
rect 22468 32376 22520 32428
rect 22928 32376 22980 32428
rect 22560 32308 22612 32360
rect 23204 32351 23256 32360
rect 23204 32317 23213 32351
rect 23213 32317 23247 32351
rect 23247 32317 23256 32351
rect 23204 32308 23256 32317
rect 24124 32240 24176 32292
rect 24952 32308 25004 32360
rect 26976 32376 27028 32428
rect 27620 32376 27672 32428
rect 38292 32419 38344 32428
rect 38292 32385 38301 32419
rect 38301 32385 38335 32419
rect 38335 32385 38344 32419
rect 38292 32376 38344 32385
rect 24860 32240 24912 32292
rect 10232 32172 10284 32224
rect 10692 32215 10744 32224
rect 10692 32181 10701 32215
rect 10701 32181 10735 32215
rect 10735 32181 10744 32215
rect 10692 32172 10744 32181
rect 18972 32172 19024 32224
rect 19340 32172 19392 32224
rect 21088 32215 21140 32224
rect 21088 32181 21097 32215
rect 21097 32181 21131 32215
rect 21131 32181 21140 32215
rect 21088 32172 21140 32181
rect 22100 32215 22152 32224
rect 22100 32181 22109 32215
rect 22109 32181 22143 32215
rect 22143 32181 22152 32215
rect 22100 32172 22152 32181
rect 23112 32172 23164 32224
rect 27528 32308 27580 32360
rect 25504 32172 25556 32224
rect 28540 32172 28592 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2964 32011 3016 32020
rect 2964 31977 2973 32011
rect 2973 31977 3007 32011
rect 3007 31977 3016 32011
rect 2964 31968 3016 31977
rect 6828 31968 6880 32020
rect 12716 31968 12768 32020
rect 15936 31968 15988 32020
rect 22100 31968 22152 32020
rect 23296 31968 23348 32020
rect 10324 31900 10376 31952
rect 2688 31832 2740 31884
rect 4160 31832 4212 31884
rect 7472 31832 7524 31884
rect 10232 31832 10284 31884
rect 15384 31900 15436 31952
rect 16764 31875 16816 31884
rect 1860 31807 1912 31816
rect 1860 31773 1869 31807
rect 1869 31773 1903 31807
rect 1903 31773 1912 31807
rect 1860 31764 1912 31773
rect 2412 31764 2464 31816
rect 3148 31807 3200 31816
rect 3148 31773 3157 31807
rect 3157 31773 3191 31807
rect 3191 31773 3200 31807
rect 3148 31764 3200 31773
rect 6460 31764 6512 31816
rect 7104 31807 7156 31816
rect 7104 31773 7113 31807
rect 7113 31773 7147 31807
rect 7147 31773 7156 31807
rect 7104 31764 7156 31773
rect 7840 31764 7892 31816
rect 8944 31764 8996 31816
rect 11796 31807 11848 31816
rect 11796 31773 11805 31807
rect 11805 31773 11839 31807
rect 11839 31773 11848 31807
rect 11796 31764 11848 31773
rect 16764 31841 16773 31875
rect 16773 31841 16807 31875
rect 16807 31841 16816 31875
rect 16764 31832 16816 31841
rect 18512 31875 18564 31884
rect 18512 31841 18521 31875
rect 18521 31841 18555 31875
rect 18555 31841 18564 31875
rect 18512 31832 18564 31841
rect 20628 31900 20680 31952
rect 22008 31832 22060 31884
rect 22192 31832 22244 31884
rect 22836 31832 22888 31884
rect 23112 31875 23164 31884
rect 23112 31841 23121 31875
rect 23121 31841 23155 31875
rect 23155 31841 23164 31875
rect 23112 31832 23164 31841
rect 23388 31900 23440 31952
rect 27620 31900 27672 31952
rect 11152 31739 11204 31748
rect 6000 31628 6052 31680
rect 10232 31628 10284 31680
rect 11152 31705 11161 31739
rect 11161 31705 11195 31739
rect 11195 31705 11204 31739
rect 11152 31696 11204 31705
rect 15936 31696 15988 31748
rect 18788 31764 18840 31816
rect 16948 31696 17000 31748
rect 17132 31696 17184 31748
rect 24768 31764 24820 31816
rect 22560 31739 22612 31748
rect 22560 31705 22569 31739
rect 22569 31705 22603 31739
rect 22603 31705 22612 31739
rect 22560 31696 22612 31705
rect 23388 31696 23440 31748
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 25780 31764 25832 31816
rect 26884 31739 26936 31748
rect 26884 31705 26893 31739
rect 26893 31705 26927 31739
rect 26927 31705 26936 31739
rect 26884 31696 26936 31705
rect 26976 31696 27028 31748
rect 27252 31696 27304 31748
rect 28356 31832 28408 31884
rect 28908 31875 28960 31884
rect 28908 31841 28917 31875
rect 28917 31841 28951 31875
rect 28951 31841 28960 31875
rect 28908 31832 28960 31841
rect 32128 31832 32180 31884
rect 30380 31764 30432 31816
rect 28080 31739 28132 31748
rect 28080 31705 28089 31739
rect 28089 31705 28123 31739
rect 28123 31705 28132 31739
rect 28080 31696 28132 31705
rect 10968 31628 11020 31680
rect 11244 31628 11296 31680
rect 22376 31628 22428 31680
rect 22928 31628 22980 31680
rect 23112 31628 23164 31680
rect 25872 31628 25924 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 3148 31424 3200 31476
rect 1768 31331 1820 31340
rect 1768 31297 1777 31331
rect 1777 31297 1811 31331
rect 1811 31297 1820 31331
rect 1768 31288 1820 31297
rect 3424 31288 3476 31340
rect 4068 31424 4120 31476
rect 6552 31424 6604 31476
rect 5356 31288 5408 31340
rect 6920 31331 6972 31340
rect 6920 31297 6929 31331
rect 6929 31297 6963 31331
rect 6963 31297 6972 31331
rect 6920 31288 6972 31297
rect 8300 31356 8352 31408
rect 23112 31424 23164 31476
rect 23572 31424 23624 31476
rect 24400 31424 24452 31476
rect 27896 31424 27948 31476
rect 12348 31399 12400 31408
rect 12348 31365 12357 31399
rect 12357 31365 12391 31399
rect 12391 31365 12400 31399
rect 12348 31356 12400 31365
rect 12440 31356 12492 31408
rect 11796 31288 11848 31340
rect 4896 31220 4948 31272
rect 6000 31263 6052 31272
rect 6000 31229 6009 31263
rect 6009 31229 6043 31263
rect 6043 31229 6052 31263
rect 6000 31220 6052 31229
rect 10692 31220 10744 31272
rect 15384 31331 15436 31340
rect 15384 31297 15393 31331
rect 15393 31297 15427 31331
rect 15427 31297 15436 31331
rect 15384 31288 15436 31297
rect 17408 31356 17460 31408
rect 22928 31356 22980 31408
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 20352 31288 20404 31340
rect 20812 31288 20864 31340
rect 21824 31288 21876 31340
rect 23480 31288 23532 31340
rect 23664 31331 23716 31340
rect 23664 31297 23673 31331
rect 23673 31297 23707 31331
rect 23707 31297 23716 31331
rect 23664 31288 23716 31297
rect 26056 31356 26108 31408
rect 27620 31356 27672 31408
rect 24952 31288 25004 31340
rect 25504 31288 25556 31340
rect 3884 31084 3936 31136
rect 11244 31152 11296 31204
rect 13912 31152 13964 31204
rect 9864 31127 9916 31136
rect 9864 31093 9873 31127
rect 9873 31093 9907 31127
rect 9907 31093 9916 31127
rect 9864 31084 9916 31093
rect 10140 31084 10192 31136
rect 16672 31220 16724 31272
rect 22192 31220 22244 31272
rect 22652 31220 22704 31272
rect 23572 31220 23624 31272
rect 23848 31220 23900 31272
rect 17500 31084 17552 31136
rect 17592 31084 17644 31136
rect 22284 31152 22336 31204
rect 25596 31152 25648 31204
rect 18604 31127 18656 31136
rect 18604 31093 18613 31127
rect 18613 31093 18647 31127
rect 18647 31093 18656 31127
rect 18604 31084 18656 31093
rect 23572 31084 23624 31136
rect 24768 31084 24820 31136
rect 27160 31331 27212 31340
rect 27160 31297 27169 31331
rect 27169 31297 27203 31331
rect 27203 31297 27212 31331
rect 27160 31288 27212 31297
rect 29092 31331 29144 31340
rect 25780 31220 25832 31272
rect 29092 31297 29101 31331
rect 29101 31297 29135 31331
rect 29135 31297 29144 31331
rect 29092 31288 29144 31297
rect 31760 31288 31812 31340
rect 32588 31288 32640 31340
rect 28448 31263 28500 31272
rect 28448 31229 28457 31263
rect 28457 31229 28491 31263
rect 28491 31229 28500 31263
rect 28448 31220 28500 31229
rect 27804 31152 27856 31204
rect 26516 31084 26568 31136
rect 26700 31084 26752 31136
rect 29184 31127 29236 31136
rect 29184 31093 29193 31127
rect 29193 31093 29227 31127
rect 29227 31093 29236 31127
rect 29184 31084 29236 31093
rect 30104 31084 30156 31136
rect 32680 31084 32732 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 17592 30880 17644 30932
rect 15752 30812 15804 30864
rect 24952 30880 25004 30932
rect 25504 30880 25556 30932
rect 17776 30812 17828 30864
rect 24032 30812 24084 30864
rect 11152 30744 11204 30796
rect 18420 30744 18472 30796
rect 20168 30744 20220 30796
rect 20444 30787 20496 30796
rect 20444 30753 20453 30787
rect 20453 30753 20487 30787
rect 20487 30753 20496 30787
rect 20444 30744 20496 30753
rect 16212 30676 16264 30728
rect 19248 30676 19300 30728
rect 19984 30676 20036 30728
rect 20260 30676 20312 30728
rect 21456 30676 21508 30728
rect 19340 30608 19392 30660
rect 20536 30651 20588 30660
rect 20536 30617 20545 30651
rect 20545 30617 20579 30651
rect 20579 30617 20588 30651
rect 21088 30651 21140 30660
rect 20536 30608 20588 30617
rect 21088 30617 21097 30651
rect 21097 30617 21131 30651
rect 21131 30617 21140 30651
rect 21824 30651 21876 30660
rect 21088 30608 21140 30617
rect 21824 30617 21833 30651
rect 21833 30617 21867 30651
rect 21867 30617 21876 30651
rect 21824 30608 21876 30617
rect 23756 30676 23808 30728
rect 27160 30880 27212 30932
rect 30104 30812 30156 30864
rect 30380 30855 30432 30864
rect 30380 30821 30389 30855
rect 30389 30821 30423 30855
rect 30423 30821 30432 30855
rect 30380 30812 30432 30821
rect 37372 30812 37424 30864
rect 29184 30744 29236 30796
rect 37464 30719 37516 30728
rect 23112 30608 23164 30660
rect 25504 30651 25556 30660
rect 25504 30617 25513 30651
rect 25513 30617 25547 30651
rect 25547 30617 25556 30651
rect 25504 30608 25556 30617
rect 25596 30651 25648 30660
rect 25596 30617 25605 30651
rect 25605 30617 25639 30651
rect 25639 30617 25648 30651
rect 37464 30685 37473 30719
rect 37473 30685 37507 30719
rect 37507 30685 37516 30719
rect 37464 30676 37516 30685
rect 29828 30651 29880 30660
rect 25596 30608 25648 30617
rect 9864 30540 9916 30592
rect 17776 30540 17828 30592
rect 18236 30540 18288 30592
rect 20168 30540 20220 30592
rect 25688 30540 25740 30592
rect 26700 30583 26752 30592
rect 26700 30549 26709 30583
rect 26709 30549 26743 30583
rect 26743 30549 26752 30583
rect 26700 30540 26752 30549
rect 27712 30540 27764 30592
rect 27896 30540 27948 30592
rect 28632 30583 28684 30592
rect 28632 30549 28641 30583
rect 28641 30549 28675 30583
rect 28675 30549 28684 30583
rect 28632 30540 28684 30549
rect 29828 30617 29837 30651
rect 29837 30617 29871 30651
rect 29871 30617 29880 30651
rect 29828 30608 29880 30617
rect 29920 30651 29972 30660
rect 29920 30617 29929 30651
rect 29929 30617 29963 30651
rect 29963 30617 29972 30651
rect 29920 30608 29972 30617
rect 32036 30540 32088 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 7104 30336 7156 30388
rect 16212 30336 16264 30388
rect 16396 30336 16448 30388
rect 18880 30336 18932 30388
rect 20536 30336 20588 30388
rect 22652 30336 22704 30388
rect 27528 30336 27580 30388
rect 16672 30268 16724 30320
rect 17316 30268 17368 30320
rect 20168 30268 20220 30320
rect 1860 30200 1912 30252
rect 2044 30243 2096 30252
rect 2044 30209 2053 30243
rect 2053 30209 2087 30243
rect 2087 30209 2096 30243
rect 2044 30200 2096 30209
rect 13452 30200 13504 30252
rect 16764 30200 16816 30252
rect 16856 30200 16908 30252
rect 19340 30200 19392 30252
rect 19708 30243 19760 30252
rect 19708 30209 19717 30243
rect 19717 30209 19751 30243
rect 19751 30209 19760 30243
rect 19708 30200 19760 30209
rect 11612 30132 11664 30184
rect 17960 30132 18012 30184
rect 23664 30268 23716 30320
rect 24124 30268 24176 30320
rect 26056 30311 26108 30320
rect 26056 30277 26065 30311
rect 26065 30277 26099 30311
rect 26099 30277 26108 30311
rect 26056 30268 26108 30277
rect 29920 30268 29972 30320
rect 20812 30243 20864 30252
rect 20812 30209 20821 30243
rect 20821 30209 20855 30243
rect 20855 30209 20864 30243
rect 20812 30200 20864 30209
rect 12992 30064 13044 30116
rect 13452 30107 13504 30116
rect 13452 30073 13461 30107
rect 13461 30073 13495 30107
rect 13495 30073 13504 30107
rect 13452 30064 13504 30073
rect 15016 30064 15068 30116
rect 16948 30064 17000 30116
rect 4712 29996 4764 30048
rect 13912 29996 13964 30048
rect 18328 30064 18380 30116
rect 22376 30175 22428 30184
rect 22376 30141 22385 30175
rect 22385 30141 22419 30175
rect 22419 30141 22428 30175
rect 22376 30132 22428 30141
rect 25044 30132 25096 30184
rect 20536 30064 20588 30116
rect 25596 30200 25648 30252
rect 28448 30200 28500 30252
rect 28724 30243 28776 30252
rect 28724 30209 28733 30243
rect 28733 30209 28767 30243
rect 28767 30209 28776 30243
rect 28724 30200 28776 30209
rect 34520 30200 34572 30252
rect 25504 30132 25556 30184
rect 27804 30175 27856 30184
rect 27804 30141 27813 30175
rect 27813 30141 27847 30175
rect 27847 30141 27856 30175
rect 27804 30132 27856 30141
rect 18696 30039 18748 30048
rect 18696 30005 18705 30039
rect 18705 30005 18739 30039
rect 18739 30005 18748 30039
rect 18696 29996 18748 30005
rect 19064 29996 19116 30048
rect 22100 29996 22152 30048
rect 22376 29996 22428 30048
rect 24032 29996 24084 30048
rect 27988 30039 28040 30048
rect 27988 30005 27997 30039
rect 27997 30005 28031 30039
rect 28031 30005 28040 30039
rect 27988 29996 28040 30005
rect 29092 29996 29144 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2320 29724 2372 29776
rect 14004 29724 14056 29776
rect 17776 29792 17828 29844
rect 18420 29792 18472 29844
rect 18880 29792 18932 29844
rect 21548 29792 21600 29844
rect 16764 29656 16816 29708
rect 17040 29656 17092 29708
rect 21640 29699 21692 29708
rect 1768 29631 1820 29640
rect 1768 29597 1777 29631
rect 1777 29597 1811 29631
rect 1811 29597 1820 29631
rect 1768 29588 1820 29597
rect 11612 29631 11664 29640
rect 11612 29597 11621 29631
rect 11621 29597 11655 29631
rect 11655 29597 11664 29631
rect 11612 29588 11664 29597
rect 18236 29588 18288 29640
rect 21640 29665 21649 29699
rect 21649 29665 21683 29699
rect 21683 29665 21692 29699
rect 21640 29656 21692 29665
rect 28632 29656 28684 29708
rect 18788 29631 18840 29640
rect 18788 29597 18797 29631
rect 18797 29597 18831 29631
rect 18831 29597 18840 29631
rect 18788 29588 18840 29597
rect 20168 29588 20220 29640
rect 20352 29588 20404 29640
rect 20904 29631 20956 29640
rect 20904 29597 20913 29631
rect 20913 29597 20947 29631
rect 20947 29597 20956 29631
rect 20904 29588 20956 29597
rect 23112 29631 23164 29640
rect 11796 29520 11848 29572
rect 13728 29520 13780 29572
rect 16672 29563 16724 29572
rect 16672 29529 16681 29563
rect 16681 29529 16715 29563
rect 16715 29529 16724 29563
rect 16672 29520 16724 29529
rect 1952 29452 2004 29504
rect 14188 29452 14240 29504
rect 18420 29520 18472 29572
rect 19432 29520 19484 29572
rect 23112 29597 23121 29631
rect 23121 29597 23155 29631
rect 23155 29597 23164 29631
rect 23112 29588 23164 29597
rect 23756 29631 23808 29640
rect 23756 29597 23765 29631
rect 23765 29597 23799 29631
rect 23799 29597 23808 29631
rect 23756 29588 23808 29597
rect 27160 29588 27212 29640
rect 36636 29588 36688 29640
rect 23388 29520 23440 29572
rect 20628 29452 20680 29504
rect 22376 29452 22428 29504
rect 22560 29452 22612 29504
rect 23756 29452 23808 29504
rect 23940 29452 23992 29504
rect 24768 29563 24820 29572
rect 24768 29529 24777 29563
rect 24777 29529 24811 29563
rect 24811 29529 24820 29563
rect 24768 29520 24820 29529
rect 24952 29520 25004 29572
rect 25228 29520 25280 29572
rect 27712 29563 27764 29572
rect 27712 29529 27721 29563
rect 27721 29529 27755 29563
rect 27755 29529 27764 29563
rect 27712 29520 27764 29529
rect 27344 29452 27396 29504
rect 27804 29452 27856 29504
rect 38200 29495 38252 29504
rect 38200 29461 38209 29495
rect 38209 29461 38243 29495
rect 38243 29461 38252 29495
rect 38200 29452 38252 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4068 29248 4120 29300
rect 5632 29180 5684 29232
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 3792 29112 3844 29164
rect 13912 29248 13964 29300
rect 11060 29180 11112 29232
rect 14188 29180 14240 29232
rect 16764 29248 16816 29300
rect 19064 29248 19116 29300
rect 19156 29248 19208 29300
rect 17224 29180 17276 29232
rect 20628 29180 20680 29232
rect 20904 29248 20956 29300
rect 22284 29248 22336 29300
rect 23112 29248 23164 29300
rect 23940 29248 23992 29300
rect 27988 29248 28040 29300
rect 24676 29180 24728 29232
rect 25320 29180 25372 29232
rect 26424 29180 26476 29232
rect 1860 29044 1912 29096
rect 4804 29044 4856 29096
rect 6552 29087 6604 29096
rect 6552 29053 6561 29087
rect 6561 29053 6595 29087
rect 6595 29053 6604 29087
rect 6552 29044 6604 29053
rect 21640 29112 21692 29164
rect 22468 29112 22520 29164
rect 26700 29112 26752 29164
rect 27988 29112 28040 29164
rect 3148 28976 3200 29028
rect 11244 29044 11296 29096
rect 11612 29044 11664 29096
rect 16120 29044 16172 29096
rect 16856 29087 16908 29096
rect 16856 29053 16865 29087
rect 16865 29053 16899 29087
rect 16899 29053 16908 29087
rect 16856 29044 16908 29053
rect 11152 28976 11204 29028
rect 16672 28976 16724 29028
rect 17868 29044 17920 29096
rect 18144 29044 18196 29096
rect 20444 29044 20496 29096
rect 23388 29044 23440 29096
rect 26056 29044 26108 29096
rect 24032 28976 24084 29028
rect 29000 29044 29052 29096
rect 1584 28951 1636 28960
rect 1584 28917 1593 28951
rect 1593 28917 1627 28951
rect 1627 28917 1636 28951
rect 1584 28908 1636 28917
rect 9680 28908 9732 28960
rect 14372 28908 14424 28960
rect 15936 28908 15988 28960
rect 16120 28908 16172 28960
rect 27804 28908 27856 28960
rect 28172 28908 28224 28960
rect 31484 28908 31536 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 9680 28704 9732 28756
rect 14004 28704 14056 28756
rect 14096 28704 14148 28756
rect 15936 28704 15988 28756
rect 18604 28704 18656 28756
rect 22100 28704 22152 28756
rect 23204 28704 23256 28756
rect 28172 28747 28224 28756
rect 28172 28713 28181 28747
rect 28181 28713 28215 28747
rect 28215 28713 28224 28747
rect 28172 28704 28224 28713
rect 12532 28636 12584 28688
rect 14556 28636 14608 28688
rect 17224 28636 17276 28688
rect 19340 28636 19392 28688
rect 19432 28636 19484 28688
rect 26424 28679 26476 28688
rect 1860 28543 1912 28552
rect 1860 28509 1869 28543
rect 1869 28509 1903 28543
rect 1903 28509 1912 28543
rect 1860 28500 1912 28509
rect 6000 28568 6052 28620
rect 3976 28500 4028 28552
rect 6552 28500 6604 28552
rect 11244 28543 11296 28552
rect 11244 28509 11253 28543
rect 11253 28509 11287 28543
rect 11287 28509 11296 28543
rect 11244 28500 11296 28509
rect 13820 28500 13872 28552
rect 14464 28543 14516 28552
rect 14464 28509 14473 28543
rect 14473 28509 14507 28543
rect 14507 28509 14516 28543
rect 14464 28500 14516 28509
rect 15200 28543 15252 28552
rect 15200 28509 15232 28543
rect 15232 28509 15252 28543
rect 15200 28500 15252 28509
rect 16580 28500 16632 28552
rect 16856 28500 16908 28552
rect 20076 28500 20128 28552
rect 20352 28500 20404 28552
rect 20628 28543 20680 28552
rect 20628 28509 20637 28543
rect 20637 28509 20671 28543
rect 20671 28509 20680 28543
rect 20628 28500 20680 28509
rect 3332 28432 3384 28484
rect 5632 28432 5684 28484
rect 11612 28432 11664 28484
rect 15752 28432 15804 28484
rect 16764 28432 16816 28484
rect 17500 28475 17552 28484
rect 2872 28407 2924 28416
rect 2872 28373 2881 28407
rect 2881 28373 2915 28407
rect 2915 28373 2924 28407
rect 2872 28364 2924 28373
rect 6000 28364 6052 28416
rect 12532 28364 12584 28416
rect 12992 28407 13044 28416
rect 12992 28373 13001 28407
rect 13001 28373 13035 28407
rect 13035 28373 13044 28407
rect 12992 28364 13044 28373
rect 13636 28407 13688 28416
rect 13636 28373 13645 28407
rect 13645 28373 13679 28407
rect 13679 28373 13688 28407
rect 13636 28364 13688 28373
rect 14004 28364 14056 28416
rect 16948 28407 17000 28416
rect 16948 28373 16957 28407
rect 16957 28373 16991 28407
rect 16991 28373 17000 28407
rect 16948 28364 17000 28373
rect 17500 28441 17509 28475
rect 17509 28441 17543 28475
rect 17543 28441 17552 28475
rect 17500 28432 17552 28441
rect 20904 28475 20956 28484
rect 20904 28441 20913 28475
rect 20913 28441 20947 28475
rect 20947 28441 20956 28475
rect 20904 28432 20956 28441
rect 21824 28500 21876 28552
rect 22284 28500 22336 28552
rect 22008 28432 22060 28484
rect 23940 28432 23992 28484
rect 24124 28432 24176 28484
rect 26424 28645 26433 28679
rect 26433 28645 26467 28679
rect 26467 28645 26476 28679
rect 26424 28636 26476 28645
rect 27804 28636 27856 28688
rect 28356 28636 28408 28688
rect 27620 28568 27672 28620
rect 17868 28364 17920 28416
rect 19432 28364 19484 28416
rect 20076 28407 20128 28416
rect 20076 28373 20085 28407
rect 20085 28373 20119 28407
rect 20119 28373 20128 28407
rect 20076 28364 20128 28373
rect 20168 28364 20220 28416
rect 24492 28364 24544 28416
rect 25596 28432 25648 28484
rect 27252 28432 27304 28484
rect 28540 28500 28592 28552
rect 29644 28500 29696 28552
rect 37280 28568 37332 28620
rect 31484 28543 31536 28552
rect 31484 28509 31493 28543
rect 31493 28509 31527 28543
rect 31527 28509 31536 28543
rect 31484 28500 31536 28509
rect 27896 28364 27948 28416
rect 33048 28364 33100 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 6000 28135 6052 28144
rect 6000 28101 6009 28135
rect 6009 28101 6043 28135
rect 6043 28101 6052 28135
rect 6000 28092 6052 28101
rect 22560 28160 22612 28212
rect 13636 28092 13688 28144
rect 15016 28092 15068 28144
rect 17224 28092 17276 28144
rect 20076 28092 20128 28144
rect 22284 28092 22336 28144
rect 23756 28135 23808 28144
rect 1768 28067 1820 28076
rect 1768 28033 1777 28067
rect 1777 28033 1811 28067
rect 1811 28033 1820 28067
rect 1768 28024 1820 28033
rect 6552 28024 6604 28076
rect 12808 28067 12860 28076
rect 12808 28033 12817 28067
rect 12817 28033 12851 28067
rect 12851 28033 12860 28067
rect 12808 28024 12860 28033
rect 14556 28024 14608 28076
rect 16764 28024 16816 28076
rect 19064 28067 19116 28076
rect 19064 28033 19073 28067
rect 19073 28033 19107 28067
rect 19107 28033 19116 28067
rect 19064 28024 19116 28033
rect 19156 28067 19208 28076
rect 19156 28033 19165 28067
rect 19165 28033 19199 28067
rect 19199 28033 19208 28067
rect 19156 28024 19208 28033
rect 20812 28024 20864 28076
rect 3976 27999 4028 28008
rect 3976 27965 3985 27999
rect 3985 27965 4019 27999
rect 4019 27965 4028 27999
rect 3976 27956 4028 27965
rect 4988 27956 5040 28008
rect 5448 27956 5500 28008
rect 2228 27820 2280 27872
rect 9956 27863 10008 27872
rect 9956 27829 9965 27863
rect 9965 27829 9999 27863
rect 9999 27829 10008 27863
rect 9956 27820 10008 27829
rect 15200 27956 15252 28008
rect 16856 27999 16908 28008
rect 16856 27965 16865 27999
rect 16865 27965 16899 27999
rect 16899 27965 16908 27999
rect 16856 27956 16908 27965
rect 17684 27956 17736 28008
rect 17868 27956 17920 28008
rect 14556 27863 14608 27872
rect 14556 27829 14565 27863
rect 14565 27829 14599 27863
rect 14599 27829 14608 27863
rect 14556 27820 14608 27829
rect 16304 27888 16356 27940
rect 18236 27888 18288 27940
rect 21916 27888 21968 27940
rect 23204 27956 23256 28008
rect 23756 28101 23765 28135
rect 23765 28101 23799 28135
rect 23799 28101 23808 28135
rect 23756 28092 23808 28101
rect 26424 28160 26476 28212
rect 29000 28203 29052 28212
rect 29000 28169 29009 28203
rect 29009 28169 29043 28203
rect 29043 28169 29052 28203
rect 29000 28160 29052 28169
rect 25688 28135 25740 28144
rect 25688 28101 25697 28135
rect 25697 28101 25731 28135
rect 25731 28101 25740 28135
rect 25688 28092 25740 28101
rect 26516 28092 26568 28144
rect 27344 28135 27396 28144
rect 27344 28101 27353 28135
rect 27353 28101 27387 28135
rect 27387 28101 27396 28135
rect 27344 28092 27396 28101
rect 28264 28092 28316 28144
rect 23296 27888 23348 27940
rect 24032 27956 24084 28008
rect 25044 28024 25096 28076
rect 29276 28092 29328 28144
rect 29184 28067 29236 28076
rect 29184 28033 29193 28067
rect 29193 28033 29227 28067
rect 29227 28033 29236 28067
rect 29184 28024 29236 28033
rect 38016 28067 38068 28076
rect 38016 28033 38025 28067
rect 38025 28033 38059 28067
rect 38059 28033 38068 28067
rect 38016 28024 38068 28033
rect 25596 27999 25648 28008
rect 25596 27965 25605 27999
rect 25605 27965 25639 27999
rect 25639 27965 25648 27999
rect 25596 27956 25648 27965
rect 27252 27999 27304 28008
rect 27252 27965 27261 27999
rect 27261 27965 27295 27999
rect 27295 27965 27304 27999
rect 27252 27956 27304 27965
rect 24860 27931 24912 27940
rect 24860 27897 24869 27931
rect 24869 27897 24903 27931
rect 24903 27897 24912 27931
rect 38200 27931 38252 27940
rect 24860 27888 24912 27897
rect 38200 27897 38209 27931
rect 38209 27897 38243 27931
rect 38243 27897 38252 27931
rect 38200 27888 38252 27897
rect 17868 27820 17920 27872
rect 18144 27820 18196 27872
rect 19432 27820 19484 27872
rect 25228 27820 25280 27872
rect 28080 27820 28132 27872
rect 28448 27863 28500 27872
rect 28448 27829 28457 27863
rect 28457 27829 28491 27863
rect 28491 27829 28500 27863
rect 28448 27820 28500 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1584 27616 1636 27668
rect 12992 27616 13044 27668
rect 17960 27616 18012 27668
rect 18052 27616 18104 27668
rect 18696 27616 18748 27668
rect 18788 27616 18840 27668
rect 20260 27616 20312 27668
rect 21548 27616 21600 27668
rect 4896 27548 4948 27600
rect 17132 27548 17184 27600
rect 19248 27548 19300 27600
rect 21824 27548 21876 27600
rect 24676 27591 24728 27600
rect 24676 27557 24685 27591
rect 24685 27557 24719 27591
rect 24719 27557 24728 27591
rect 24676 27548 24728 27557
rect 24768 27548 24820 27600
rect 3976 27480 4028 27532
rect 12808 27480 12860 27532
rect 15200 27480 15252 27532
rect 16212 27480 16264 27532
rect 16488 27480 16540 27532
rect 21364 27480 21416 27532
rect 4804 27412 4856 27464
rect 5264 27412 5316 27464
rect 18236 27412 18288 27464
rect 18604 27412 18656 27464
rect 19432 27412 19484 27464
rect 23388 27455 23440 27464
rect 23388 27421 23397 27455
rect 23397 27421 23431 27455
rect 23431 27421 23440 27455
rect 23388 27412 23440 27421
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 24860 27412 24912 27464
rect 25320 27455 25372 27464
rect 25320 27421 25329 27455
rect 25329 27421 25363 27455
rect 25363 27421 25372 27455
rect 27344 27548 27396 27600
rect 29184 27548 29236 27600
rect 36636 27548 36688 27600
rect 25320 27412 25372 27421
rect 3148 27344 3200 27396
rect 3516 27344 3568 27396
rect 10508 27344 10560 27396
rect 16396 27344 16448 27396
rect 17408 27344 17460 27396
rect 21364 27387 21416 27396
rect 21364 27353 21373 27387
rect 21373 27353 21407 27387
rect 21407 27353 21416 27387
rect 21364 27344 21416 27353
rect 22008 27387 22060 27396
rect 22008 27353 22017 27387
rect 22017 27353 22051 27387
rect 22051 27353 22060 27387
rect 22928 27387 22980 27396
rect 22008 27344 22060 27353
rect 22928 27353 22937 27387
rect 22937 27353 22971 27387
rect 22971 27353 22980 27387
rect 22928 27344 22980 27353
rect 27436 27412 27488 27464
rect 28356 27480 28408 27532
rect 28540 27412 28592 27464
rect 30380 27455 30432 27464
rect 28356 27344 28408 27396
rect 30380 27421 30389 27455
rect 30389 27421 30423 27455
rect 30423 27421 30432 27455
rect 30380 27412 30432 27421
rect 31576 27412 31628 27464
rect 33048 27412 33100 27464
rect 37464 27344 37516 27396
rect 37924 27344 37976 27396
rect 7012 27276 7064 27328
rect 11520 27319 11572 27328
rect 11520 27285 11529 27319
rect 11529 27285 11563 27319
rect 11563 27285 11572 27319
rect 11520 27276 11572 27285
rect 12992 27276 13044 27328
rect 21824 27276 21876 27328
rect 23480 27319 23532 27328
rect 23480 27285 23489 27319
rect 23489 27285 23523 27319
rect 23523 27285 23532 27319
rect 23480 27276 23532 27285
rect 24216 27276 24268 27328
rect 24768 27276 24820 27328
rect 26424 27276 26476 27328
rect 27344 27276 27396 27328
rect 27988 27276 28040 27328
rect 30472 27319 30524 27328
rect 30472 27285 30481 27319
rect 30481 27285 30515 27319
rect 30515 27285 30524 27319
rect 30472 27276 30524 27285
rect 38200 27319 38252 27328
rect 38200 27285 38209 27319
rect 38209 27285 38243 27319
rect 38243 27285 38252 27319
rect 38200 27276 38252 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 22008 27072 22060 27124
rect 22100 27072 22152 27124
rect 31576 27115 31628 27124
rect 3976 27004 4028 27056
rect 4712 27004 4764 27056
rect 13728 27047 13780 27056
rect 13728 27013 13737 27047
rect 13737 27013 13771 27047
rect 13771 27013 13780 27047
rect 13728 27004 13780 27013
rect 17132 27047 17184 27056
rect 17132 27013 17141 27047
rect 17141 27013 17175 27047
rect 17175 27013 17184 27047
rect 17132 27004 17184 27013
rect 19156 27004 19208 27056
rect 19340 27004 19392 27056
rect 22468 27004 22520 27056
rect 24216 27004 24268 27056
rect 24492 27047 24544 27056
rect 24492 27013 24501 27047
rect 24501 27013 24535 27047
rect 24535 27013 24544 27047
rect 24492 27004 24544 27013
rect 1676 26979 1728 26988
rect 1676 26945 1685 26979
rect 1685 26945 1719 26979
rect 1719 26945 1728 26979
rect 1676 26936 1728 26945
rect 11244 26936 11296 26988
rect 13084 26936 13136 26988
rect 16856 26979 16908 26988
rect 1860 26843 1912 26852
rect 1860 26809 1869 26843
rect 1869 26809 1903 26843
rect 1903 26809 1912 26843
rect 1860 26800 1912 26809
rect 9220 26868 9272 26920
rect 16856 26945 16865 26979
rect 16865 26945 16899 26979
rect 16899 26945 16908 26979
rect 16856 26936 16908 26945
rect 18512 26936 18564 26988
rect 18972 26936 19024 26988
rect 19248 26936 19300 26988
rect 31576 27081 31585 27115
rect 31585 27081 31619 27115
rect 31619 27081 31628 27115
rect 31576 27072 31628 27081
rect 38384 27072 38436 27124
rect 27344 27047 27396 27056
rect 27344 27013 27353 27047
rect 27353 27013 27387 27047
rect 27387 27013 27396 27047
rect 27344 27004 27396 27013
rect 29184 26936 29236 26988
rect 37924 26936 37976 26988
rect 4068 26732 4120 26784
rect 5356 26732 5408 26784
rect 11060 26732 11112 26784
rect 19892 26868 19944 26920
rect 18972 26800 19024 26852
rect 21640 26868 21692 26920
rect 23204 26868 23256 26920
rect 23848 26911 23900 26920
rect 23848 26877 23857 26911
rect 23857 26877 23891 26911
rect 23891 26877 23900 26911
rect 23848 26868 23900 26877
rect 21364 26800 21416 26852
rect 24216 26800 24268 26852
rect 24952 26868 25004 26920
rect 26516 26868 26568 26920
rect 27896 26868 27948 26920
rect 28172 26911 28224 26920
rect 28172 26877 28181 26911
rect 28181 26877 28215 26911
rect 28215 26877 28224 26911
rect 28172 26868 28224 26877
rect 30472 26800 30524 26852
rect 18788 26732 18840 26784
rect 21640 26732 21692 26784
rect 24584 26732 24636 26784
rect 27528 26732 27580 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5448 26528 5500 26580
rect 12992 26528 13044 26580
rect 13084 26528 13136 26580
rect 23940 26528 23992 26580
rect 29184 26571 29236 26580
rect 29184 26537 29193 26571
rect 29193 26537 29227 26571
rect 29227 26537 29236 26571
rect 29184 26528 29236 26537
rect 30380 26528 30432 26580
rect 15752 26460 15804 26512
rect 2412 26435 2464 26444
rect 2412 26401 2421 26435
rect 2421 26401 2455 26435
rect 2455 26401 2464 26435
rect 2412 26392 2464 26401
rect 7932 26392 7984 26444
rect 6092 26324 6144 26376
rect 2872 26256 2924 26308
rect 3424 26299 3476 26308
rect 3424 26265 3433 26299
rect 3433 26265 3467 26299
rect 3467 26265 3476 26299
rect 3424 26256 3476 26265
rect 6644 26256 6696 26308
rect 7012 26256 7064 26308
rect 12256 26392 12308 26444
rect 16856 26392 16908 26444
rect 17316 26392 17368 26444
rect 19248 26460 19300 26512
rect 19984 26460 20036 26512
rect 20168 26392 20220 26444
rect 22744 26392 22796 26444
rect 26424 26435 26476 26444
rect 18788 26324 18840 26376
rect 10508 26299 10560 26308
rect 10508 26265 10517 26299
rect 10517 26265 10551 26299
rect 10551 26265 10560 26299
rect 10508 26256 10560 26265
rect 11152 26256 11204 26308
rect 16580 26256 16632 26308
rect 16948 26256 17000 26308
rect 19248 26256 19300 26308
rect 20076 26324 20128 26376
rect 20352 26367 20404 26376
rect 20352 26333 20361 26367
rect 20361 26333 20395 26367
rect 20395 26333 20404 26367
rect 20352 26324 20404 26333
rect 22468 26324 22520 26376
rect 22652 26367 22704 26376
rect 22652 26333 22661 26367
rect 22661 26333 22695 26367
rect 22695 26333 22704 26367
rect 22652 26324 22704 26333
rect 22836 26324 22888 26376
rect 26424 26401 26433 26435
rect 26433 26401 26467 26435
rect 26467 26401 26476 26435
rect 26424 26392 26476 26401
rect 38016 26460 38068 26512
rect 36360 26392 36412 26444
rect 23388 26367 23440 26376
rect 23388 26333 23397 26367
rect 23397 26333 23431 26367
rect 23431 26333 23440 26367
rect 23388 26324 23440 26333
rect 24492 26324 24544 26376
rect 25044 26324 25096 26376
rect 26516 26324 26568 26376
rect 28540 26367 28592 26376
rect 28540 26333 28549 26367
rect 28549 26333 28583 26367
rect 28583 26333 28592 26367
rect 28540 26324 28592 26333
rect 28724 26367 28776 26376
rect 28724 26333 28733 26367
rect 28733 26333 28767 26367
rect 28767 26333 28776 26367
rect 28724 26324 28776 26333
rect 29092 26324 29144 26376
rect 38292 26367 38344 26376
rect 38292 26333 38301 26367
rect 38301 26333 38335 26367
rect 38335 26333 38344 26367
rect 38292 26324 38344 26333
rect 20444 26299 20496 26308
rect 20444 26265 20453 26299
rect 20453 26265 20487 26299
rect 20487 26265 20496 26299
rect 20444 26256 20496 26265
rect 17224 26188 17276 26240
rect 24768 26256 24820 26308
rect 22284 26188 22336 26240
rect 24952 26188 25004 26240
rect 25320 26231 25372 26240
rect 25320 26197 25329 26231
rect 25329 26197 25363 26231
rect 25363 26197 25372 26231
rect 25320 26188 25372 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 10784 26027 10836 26036
rect 10784 25993 10793 26027
rect 10793 25993 10827 26027
rect 10827 25993 10836 26027
rect 10784 25984 10836 25993
rect 3884 25916 3936 25968
rect 18420 25984 18472 26036
rect 19156 26027 19208 26036
rect 19156 25993 19165 26027
rect 19165 25993 19199 26027
rect 19199 25993 19208 26027
rect 19156 25984 19208 25993
rect 17224 25916 17276 25968
rect 20444 25916 20496 25968
rect 20536 25916 20588 25968
rect 24492 25984 24544 26036
rect 28540 25984 28592 26036
rect 23480 25916 23532 25968
rect 26608 25916 26660 25968
rect 27528 25916 27580 25968
rect 3792 25848 3844 25900
rect 12256 25891 12308 25900
rect 12256 25857 12265 25891
rect 12265 25857 12299 25891
rect 12299 25857 12308 25891
rect 12256 25848 12308 25857
rect 18788 25848 18840 25900
rect 19156 25848 19208 25900
rect 22284 25891 22336 25900
rect 22284 25857 22293 25891
rect 22293 25857 22327 25891
rect 22327 25857 22336 25891
rect 22284 25848 22336 25857
rect 4068 25780 4120 25832
rect 4528 25780 4580 25832
rect 6092 25780 6144 25832
rect 7472 25780 7524 25832
rect 9956 25780 10008 25832
rect 3700 25644 3752 25696
rect 6644 25644 6696 25696
rect 12624 25780 12676 25832
rect 12900 25780 12952 25832
rect 16028 25780 16080 25832
rect 16856 25823 16908 25832
rect 16856 25789 16865 25823
rect 16865 25789 16899 25823
rect 16899 25789 16908 25823
rect 16856 25780 16908 25789
rect 18144 25780 18196 25832
rect 18420 25780 18472 25832
rect 22468 25823 22520 25832
rect 18328 25712 18380 25764
rect 22468 25789 22477 25823
rect 22477 25789 22511 25823
rect 22511 25789 22520 25823
rect 22468 25780 22520 25789
rect 24216 25780 24268 25832
rect 24308 25780 24360 25832
rect 18236 25644 18288 25696
rect 18604 25687 18656 25696
rect 18604 25653 18613 25687
rect 18613 25653 18647 25687
rect 18647 25653 18656 25687
rect 18604 25644 18656 25653
rect 18696 25644 18748 25696
rect 25320 25712 25372 25764
rect 29920 25780 29972 25832
rect 30840 25823 30892 25832
rect 30840 25789 30849 25823
rect 30849 25789 30883 25823
rect 30883 25789 30892 25823
rect 30840 25780 30892 25789
rect 30288 25644 30340 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 18604 25440 18656 25492
rect 16028 25372 16080 25424
rect 19064 25372 19116 25424
rect 19156 25372 19208 25424
rect 19892 25372 19944 25424
rect 6092 25347 6144 25356
rect 6092 25313 6101 25347
rect 6101 25313 6135 25347
rect 6135 25313 6144 25347
rect 6092 25304 6144 25313
rect 8024 25304 8076 25356
rect 20168 25347 20220 25356
rect 20168 25313 20178 25347
rect 20178 25313 20212 25347
rect 20212 25313 20220 25347
rect 23664 25440 23716 25492
rect 25320 25440 25372 25492
rect 27804 25440 27856 25492
rect 28264 25440 28316 25492
rect 28724 25440 28776 25492
rect 23296 25372 23348 25424
rect 26792 25372 26844 25424
rect 20168 25304 20220 25313
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 3608 25236 3660 25288
rect 4068 25236 4120 25288
rect 14280 25236 14332 25288
rect 18052 25279 18104 25288
rect 18052 25245 18061 25279
rect 18061 25245 18095 25279
rect 18095 25245 18104 25279
rect 18052 25236 18104 25245
rect 18236 25236 18288 25288
rect 21640 25279 21692 25288
rect 21640 25245 21649 25279
rect 21649 25245 21683 25279
rect 21683 25245 21692 25279
rect 21640 25236 21692 25245
rect 22284 25279 22336 25288
rect 22284 25245 22293 25279
rect 22293 25245 22327 25279
rect 22327 25245 22336 25279
rect 22284 25236 22336 25245
rect 23112 25236 23164 25288
rect 23480 25236 23532 25288
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 25504 25236 25556 25288
rect 29092 25304 29144 25356
rect 29920 25347 29972 25356
rect 29920 25313 29929 25347
rect 29929 25313 29963 25347
rect 29963 25313 29972 25347
rect 29920 25304 29972 25313
rect 27068 25279 27120 25288
rect 27068 25245 27077 25279
rect 27077 25245 27111 25279
rect 27111 25245 27120 25279
rect 27068 25236 27120 25245
rect 28356 25279 28408 25288
rect 28356 25245 28365 25279
rect 28365 25245 28399 25279
rect 28399 25245 28408 25279
rect 28356 25236 28408 25245
rect 5632 25168 5684 25220
rect 6368 25211 6420 25220
rect 6368 25177 6377 25211
rect 6377 25177 6411 25211
rect 6411 25177 6420 25211
rect 6368 25168 6420 25177
rect 11060 25168 11112 25220
rect 1768 25143 1820 25152
rect 1768 25109 1777 25143
rect 1777 25109 1811 25143
rect 1811 25109 1820 25143
rect 1768 25100 1820 25109
rect 7104 25100 7156 25152
rect 16488 25143 16540 25152
rect 16488 25109 16497 25143
rect 16497 25109 16531 25143
rect 16531 25109 16540 25143
rect 16488 25100 16540 25109
rect 19800 25168 19852 25220
rect 20444 25168 20496 25220
rect 21180 25211 21232 25220
rect 21180 25177 21189 25211
rect 21189 25177 21223 25211
rect 21223 25177 21232 25211
rect 21180 25168 21232 25177
rect 21364 25168 21416 25220
rect 23848 25168 23900 25220
rect 24492 25168 24544 25220
rect 24768 25211 24820 25220
rect 24768 25177 24777 25211
rect 24777 25177 24811 25211
rect 24811 25177 24820 25211
rect 31760 25236 31812 25288
rect 24768 25168 24820 25177
rect 19248 25100 19300 25152
rect 19984 25100 20036 25152
rect 21916 25100 21968 25152
rect 23572 25100 23624 25152
rect 24860 25100 24912 25152
rect 27160 25143 27212 25152
rect 27160 25109 27169 25143
rect 27169 25109 27203 25143
rect 27203 25109 27212 25143
rect 27160 25100 27212 25109
rect 31576 25143 31628 25152
rect 31576 25109 31585 25143
rect 31585 25109 31619 25143
rect 31619 25109 31628 25143
rect 31576 25100 31628 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4620 24828 4672 24880
rect 1400 24760 1452 24812
rect 16304 24896 16356 24948
rect 18052 24896 18104 24948
rect 18144 24896 18196 24948
rect 23112 24896 23164 24948
rect 24216 24896 24268 24948
rect 27896 24896 27948 24948
rect 16488 24828 16540 24880
rect 7748 24760 7800 24812
rect 3608 24735 3660 24744
rect 3608 24701 3617 24735
rect 3617 24701 3651 24735
rect 3651 24701 3660 24735
rect 3608 24692 3660 24701
rect 13268 24735 13320 24744
rect 13268 24701 13277 24735
rect 13277 24701 13311 24735
rect 13311 24701 13320 24735
rect 13268 24692 13320 24701
rect 14188 24692 14240 24744
rect 15200 24760 15252 24812
rect 17500 24760 17552 24812
rect 18328 24803 18380 24812
rect 18328 24769 18337 24803
rect 18337 24769 18371 24803
rect 18371 24769 18380 24803
rect 18328 24760 18380 24769
rect 20076 24828 20128 24880
rect 23572 24828 23624 24880
rect 24952 24871 25004 24880
rect 24952 24837 24961 24871
rect 24961 24837 24995 24871
rect 24995 24837 25004 24871
rect 24952 24828 25004 24837
rect 15016 24735 15068 24744
rect 15016 24701 15025 24735
rect 15025 24701 15059 24735
rect 15059 24701 15068 24735
rect 15016 24692 15068 24701
rect 16948 24692 17000 24744
rect 17684 24692 17736 24744
rect 19340 24692 19392 24744
rect 20444 24692 20496 24744
rect 21180 24735 21232 24744
rect 21180 24701 21189 24735
rect 21189 24701 21223 24735
rect 21223 24701 21232 24735
rect 21640 24760 21692 24812
rect 22192 24803 22244 24812
rect 22192 24769 22201 24803
rect 22201 24769 22235 24803
rect 22235 24769 22244 24803
rect 22192 24760 22244 24769
rect 22560 24760 22612 24812
rect 23480 24760 23532 24812
rect 25596 24760 25648 24812
rect 27160 24760 27212 24812
rect 21180 24692 21232 24701
rect 2688 24556 2740 24608
rect 6828 24556 6880 24608
rect 17500 24556 17552 24608
rect 18420 24599 18472 24608
rect 18420 24565 18429 24599
rect 18429 24565 18463 24599
rect 18463 24565 18472 24599
rect 18420 24556 18472 24565
rect 22468 24692 22520 24744
rect 23388 24692 23440 24744
rect 22836 24624 22888 24676
rect 37832 24760 37884 24812
rect 38016 24803 38068 24812
rect 38016 24769 38025 24803
rect 38025 24769 38059 24803
rect 38059 24769 38068 24803
rect 38016 24760 38068 24769
rect 29276 24692 29328 24744
rect 22100 24556 22152 24608
rect 25504 24556 25556 24608
rect 27160 24599 27212 24608
rect 27160 24565 27169 24599
rect 27169 24565 27203 24599
rect 27203 24565 27212 24599
rect 27160 24556 27212 24565
rect 28356 24556 28408 24608
rect 29092 24599 29144 24608
rect 29092 24565 29101 24599
rect 29101 24565 29135 24599
rect 29135 24565 29144 24599
rect 29092 24556 29144 24565
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 6828 24395 6880 24404
rect 6828 24361 6837 24395
rect 6837 24361 6871 24395
rect 6871 24361 6880 24395
rect 6828 24352 6880 24361
rect 6920 24352 6972 24404
rect 9404 24352 9456 24404
rect 22192 24352 22244 24404
rect 3608 24216 3660 24268
rect 5356 24259 5408 24268
rect 5356 24225 5365 24259
rect 5365 24225 5399 24259
rect 5399 24225 5408 24259
rect 5356 24216 5408 24225
rect 7472 24216 7524 24268
rect 12256 24216 12308 24268
rect 4712 24148 4764 24200
rect 3332 24080 3384 24132
rect 6736 24080 6788 24132
rect 11520 24080 11572 24132
rect 11888 24080 11940 24132
rect 14280 24216 14332 24268
rect 16856 24216 16908 24268
rect 18696 24284 18748 24336
rect 19248 24284 19300 24336
rect 22836 24284 22888 24336
rect 23112 24284 23164 24336
rect 25596 24352 25648 24404
rect 32496 24352 32548 24404
rect 37832 24352 37884 24404
rect 13268 24080 13320 24132
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 8116 24012 8168 24064
rect 15200 24012 15252 24064
rect 16764 24123 16816 24132
rect 16764 24089 16773 24123
rect 16773 24089 16807 24123
rect 16807 24089 16816 24123
rect 16764 24080 16816 24089
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 19248 24148 19300 24200
rect 20352 24148 20404 24200
rect 21456 24148 21508 24200
rect 21824 24191 21876 24200
rect 21824 24157 21833 24191
rect 21833 24157 21867 24191
rect 21867 24157 21876 24191
rect 21824 24148 21876 24157
rect 21916 24148 21968 24200
rect 22560 24148 22612 24200
rect 23112 24191 23164 24200
rect 18144 24012 18196 24064
rect 19156 24080 19208 24132
rect 20720 24123 20772 24132
rect 20720 24089 20729 24123
rect 20729 24089 20763 24123
rect 20763 24089 20772 24123
rect 20720 24080 20772 24089
rect 18788 24055 18840 24064
rect 18788 24021 18797 24055
rect 18797 24021 18831 24055
rect 18831 24021 18840 24055
rect 18788 24012 18840 24021
rect 18880 24012 18932 24064
rect 20628 24012 20680 24064
rect 22192 24080 22244 24132
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 27160 24284 27212 24336
rect 38016 24284 38068 24336
rect 24952 24216 25004 24268
rect 26884 24216 26936 24268
rect 26148 24191 26200 24200
rect 26148 24157 26157 24191
rect 26157 24157 26191 24191
rect 26191 24157 26200 24191
rect 26148 24148 26200 24157
rect 22744 24012 22796 24064
rect 23296 24012 23348 24064
rect 24860 24080 24912 24132
rect 25688 24123 25740 24132
rect 25688 24089 25697 24123
rect 25697 24089 25731 24123
rect 25731 24089 25740 24123
rect 25688 24080 25740 24089
rect 25504 24012 25556 24064
rect 25596 24012 25648 24064
rect 38292 24191 38344 24200
rect 38292 24157 38301 24191
rect 38301 24157 38335 24191
rect 38335 24157 38344 24191
rect 38292 24148 38344 24157
rect 26884 24055 26936 24064
rect 26884 24021 26893 24055
rect 26893 24021 26927 24055
rect 26927 24021 26936 24055
rect 26884 24012 26936 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4620 23808 4672 23860
rect 4712 23808 4764 23860
rect 5540 23808 5592 23860
rect 5724 23808 5776 23860
rect 9220 23851 9272 23860
rect 9220 23817 9229 23851
rect 9229 23817 9263 23851
rect 9263 23817 9272 23851
rect 9220 23808 9272 23817
rect 2780 23740 2832 23792
rect 3700 23740 3752 23792
rect 5264 23715 5316 23724
rect 5264 23681 5273 23715
rect 5273 23681 5307 23715
rect 5307 23681 5316 23715
rect 5264 23672 5316 23681
rect 5724 23672 5776 23724
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 7472 23715 7524 23724
rect 7472 23681 7481 23715
rect 7481 23681 7515 23715
rect 7515 23681 7524 23715
rect 7472 23672 7524 23681
rect 12072 23672 12124 23724
rect 13912 23808 13964 23860
rect 14372 23808 14424 23860
rect 15016 23851 15068 23860
rect 15016 23817 15025 23851
rect 15025 23817 15059 23851
rect 15059 23817 15068 23851
rect 15016 23808 15068 23817
rect 16764 23808 16816 23860
rect 21824 23808 21876 23860
rect 25504 23851 25556 23860
rect 25504 23817 25513 23851
rect 25513 23817 25547 23851
rect 25547 23817 25556 23851
rect 25504 23808 25556 23817
rect 26148 23808 26200 23860
rect 29000 23808 29052 23860
rect 2412 23647 2464 23656
rect 2412 23613 2421 23647
rect 2421 23613 2455 23647
rect 2455 23613 2464 23647
rect 2412 23604 2464 23613
rect 4896 23604 4948 23656
rect 5080 23604 5132 23656
rect 7288 23604 7340 23656
rect 7748 23647 7800 23656
rect 7748 23613 7757 23647
rect 7757 23613 7791 23647
rect 7791 23613 7800 23647
rect 7748 23604 7800 23613
rect 11244 23604 11296 23656
rect 18420 23740 18472 23792
rect 19984 23740 20036 23792
rect 22560 23783 22612 23792
rect 22560 23749 22569 23783
rect 22569 23749 22603 23783
rect 22603 23749 22612 23783
rect 22560 23740 22612 23749
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 24676 23672 24728 23724
rect 26884 23740 26936 23792
rect 25780 23672 25832 23724
rect 13268 23647 13320 23656
rect 13268 23613 13277 23647
rect 13277 23613 13311 23647
rect 13311 23613 13320 23647
rect 13268 23604 13320 23613
rect 13544 23647 13596 23656
rect 13544 23613 13553 23647
rect 13553 23613 13587 23647
rect 13587 23613 13596 23647
rect 13544 23604 13596 23613
rect 18604 23604 18656 23656
rect 19432 23604 19484 23656
rect 19984 23604 20036 23656
rect 20444 23647 20496 23656
rect 20444 23613 20476 23647
rect 20476 23613 20496 23647
rect 20444 23604 20496 23613
rect 4620 23536 4672 23588
rect 21640 23604 21692 23656
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 22928 23647 22980 23656
rect 22928 23613 22937 23647
rect 22937 23613 22971 23647
rect 22971 23613 22980 23647
rect 22928 23604 22980 23613
rect 29092 23604 29144 23656
rect 31116 23604 31168 23656
rect 2780 23468 2832 23520
rect 5264 23468 5316 23520
rect 5356 23468 5408 23520
rect 26976 23536 27028 23588
rect 9128 23468 9180 23520
rect 13728 23468 13780 23520
rect 13912 23468 13964 23520
rect 16856 23468 16908 23520
rect 19156 23468 19208 23520
rect 20628 23468 20680 23520
rect 20720 23468 20772 23520
rect 23388 23468 23440 23520
rect 23756 23468 23808 23520
rect 25964 23468 26016 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 5264 23264 5316 23316
rect 3976 23128 4028 23180
rect 12256 23128 12308 23180
rect 1952 23060 2004 23112
rect 5540 23060 5592 23112
rect 5632 23060 5684 23112
rect 6736 23060 6788 23112
rect 9588 23060 9640 23112
rect 20536 23264 20588 23316
rect 24768 23264 24820 23316
rect 26976 23264 27028 23316
rect 27252 23264 27304 23316
rect 29828 23307 29880 23316
rect 29828 23273 29837 23307
rect 29837 23273 29871 23307
rect 29871 23273 29880 23307
rect 29828 23264 29880 23273
rect 17224 23196 17276 23248
rect 22100 23196 22152 23248
rect 22284 23196 22336 23248
rect 25136 23196 25188 23248
rect 25688 23196 25740 23248
rect 30840 23196 30892 23248
rect 16488 23128 16540 23180
rect 16856 23128 16908 23180
rect 19248 23128 19300 23180
rect 20536 23171 20588 23180
rect 20536 23137 20545 23171
rect 20545 23137 20579 23171
rect 20579 23137 20588 23171
rect 20536 23128 20588 23137
rect 20996 23128 21048 23180
rect 21916 23128 21968 23180
rect 31116 23171 31168 23180
rect 14280 23103 14332 23112
rect 9496 22992 9548 23044
rect 10784 22992 10836 23044
rect 11704 22992 11756 23044
rect 12256 22992 12308 23044
rect 14280 23069 14289 23103
rect 14289 23069 14323 23103
rect 14323 23069 14332 23103
rect 14280 23060 14332 23069
rect 18512 23060 18564 23112
rect 18972 23060 19024 23112
rect 20720 23060 20772 23112
rect 13820 22992 13872 23044
rect 14556 22992 14608 23044
rect 1860 22924 1912 22976
rect 5540 22924 5592 22976
rect 7012 22924 7064 22976
rect 7564 22924 7616 22976
rect 13728 22924 13780 22976
rect 20812 22992 20864 23044
rect 20996 22992 21048 23044
rect 14740 22924 14792 22976
rect 16580 22924 16632 22976
rect 17408 22924 17460 22976
rect 24400 23060 24452 23112
rect 31116 23137 31125 23171
rect 31125 23137 31159 23171
rect 31159 23137 31168 23171
rect 31116 23128 31168 23137
rect 22652 23035 22704 23044
rect 22652 23001 22661 23035
rect 22661 23001 22695 23035
rect 22695 23001 22704 23035
rect 22652 22992 22704 23001
rect 22744 23035 22796 23044
rect 22744 23001 22753 23035
rect 22753 23001 22787 23035
rect 22787 23001 22796 23035
rect 22744 22992 22796 23001
rect 23020 22992 23072 23044
rect 23940 22992 23992 23044
rect 23480 22924 23532 22976
rect 24768 23035 24820 23044
rect 24768 23001 24777 23035
rect 24777 23001 24811 23035
rect 24811 23001 24820 23035
rect 24768 22992 24820 23001
rect 24400 22924 24452 22976
rect 26424 22967 26476 22976
rect 26424 22933 26433 22967
rect 26433 22933 26467 22967
rect 26467 22933 26476 22967
rect 26424 22924 26476 22933
rect 36084 23060 36136 23112
rect 30288 22992 30340 23044
rect 32128 23035 32180 23044
rect 32128 23001 32137 23035
rect 32137 23001 32171 23035
rect 32171 23001 32180 23035
rect 32128 22992 32180 23001
rect 37648 22924 37700 22976
rect 38016 22924 38068 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 2412 22720 2464 22772
rect 3700 22720 3752 22772
rect 2044 22652 2096 22704
rect 10692 22720 10744 22772
rect 10784 22720 10836 22772
rect 17224 22720 17276 22772
rect 9588 22652 9640 22704
rect 12440 22652 12492 22704
rect 12808 22652 12860 22704
rect 14188 22652 14240 22704
rect 14556 22652 14608 22704
rect 18236 22652 18288 22704
rect 6920 22584 6972 22636
rect 7472 22584 7524 22636
rect 12256 22627 12308 22636
rect 7104 22516 7156 22568
rect 12256 22593 12265 22627
rect 12265 22593 12299 22627
rect 12299 22593 12308 22627
rect 12256 22584 12308 22593
rect 21364 22652 21416 22704
rect 24400 22695 24452 22704
rect 24400 22661 24409 22695
rect 24409 22661 24443 22695
rect 24443 22661 24452 22695
rect 24400 22652 24452 22661
rect 24952 22695 25004 22704
rect 24952 22661 24961 22695
rect 24961 22661 24995 22695
rect 24995 22661 25004 22695
rect 24952 22652 25004 22661
rect 28448 22720 28500 22772
rect 36084 22763 36136 22772
rect 36084 22729 36093 22763
rect 36093 22729 36127 22763
rect 36127 22729 36136 22763
rect 36084 22720 36136 22729
rect 9496 22559 9548 22568
rect 9496 22525 9505 22559
rect 9505 22525 9539 22559
rect 9539 22525 9548 22559
rect 9496 22516 9548 22525
rect 12624 22516 12676 22568
rect 18696 22584 18748 22636
rect 27344 22584 27396 22636
rect 30840 22584 30892 22636
rect 38016 22627 38068 22636
rect 38016 22593 38025 22627
rect 38025 22593 38059 22627
rect 38059 22593 38068 22627
rect 38016 22584 38068 22593
rect 24308 22559 24360 22568
rect 24308 22525 24317 22559
rect 24317 22525 24351 22559
rect 24351 22525 24360 22559
rect 24308 22516 24360 22525
rect 26608 22559 26660 22568
rect 26608 22525 26617 22559
rect 26617 22525 26651 22559
rect 26651 22525 26660 22559
rect 26608 22516 26660 22525
rect 3424 22380 3476 22432
rect 18788 22448 18840 22500
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 17592 22380 17644 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3608 22176 3660 22228
rect 7472 22176 7524 22228
rect 8208 22176 8260 22228
rect 12164 22176 12216 22228
rect 14740 22176 14792 22228
rect 8116 22108 8168 22160
rect 3700 22040 3752 22092
rect 5264 22040 5316 22092
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 11520 22040 11572 22092
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 8392 21972 8444 22024
rect 13820 22108 13872 22160
rect 11796 21972 11848 22024
rect 12348 21972 12400 22024
rect 23388 22040 23440 22092
rect 26884 22108 26936 22160
rect 15108 22015 15160 22024
rect 15108 21981 15117 22015
rect 15117 21981 15151 22015
rect 15151 21981 15160 22015
rect 15108 21972 15160 21981
rect 20076 21972 20128 22024
rect 22100 21972 22152 22024
rect 4712 21904 4764 21956
rect 5540 21904 5592 21956
rect 11520 21904 11572 21956
rect 12716 21904 12768 21956
rect 15384 21947 15436 21956
rect 15384 21913 15393 21947
rect 15393 21913 15427 21947
rect 15427 21913 15436 21947
rect 15384 21904 15436 21913
rect 17592 21904 17644 21956
rect 20168 21904 20220 21956
rect 26424 22040 26476 22092
rect 28172 22040 28224 22092
rect 27436 21972 27488 22024
rect 25964 21947 26016 21956
rect 25964 21913 25973 21947
rect 25973 21913 26007 21947
rect 26007 21913 26016 21947
rect 26884 21947 26936 21956
rect 25964 21904 26016 21913
rect 26884 21913 26893 21947
rect 26893 21913 26927 21947
rect 26927 21913 26936 21947
rect 26884 21904 26936 21913
rect 26976 21904 27028 21956
rect 28448 21972 28500 22024
rect 36636 21972 36688 22024
rect 1768 21879 1820 21888
rect 1768 21845 1777 21879
rect 1777 21845 1811 21879
rect 1811 21845 1820 21879
rect 1768 21836 1820 21845
rect 8116 21836 8168 21888
rect 8760 21836 8812 21888
rect 8944 21836 8996 21888
rect 10416 21836 10468 21888
rect 17316 21836 17368 21888
rect 17868 21836 17920 21888
rect 20628 21836 20680 21888
rect 26240 21836 26292 21888
rect 27988 21836 28040 21888
rect 29828 21879 29880 21888
rect 29828 21845 29837 21879
rect 29837 21845 29871 21879
rect 29871 21845 29880 21879
rect 29828 21836 29880 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4988 21632 5040 21684
rect 5172 21632 5224 21684
rect 5264 21632 5316 21684
rect 7380 21632 7432 21684
rect 7564 21632 7616 21684
rect 8024 21632 8076 21684
rect 8208 21632 8260 21684
rect 7196 21564 7248 21616
rect 9864 21564 9916 21616
rect 1768 21539 1820 21548
rect 1768 21505 1777 21539
rect 1777 21505 1811 21539
rect 1811 21505 1820 21539
rect 1768 21496 1820 21505
rect 3976 21539 4028 21548
rect 3976 21505 3985 21539
rect 3985 21505 4019 21539
rect 4019 21505 4028 21539
rect 3976 21496 4028 21505
rect 5356 21496 5408 21548
rect 4252 21471 4304 21480
rect 4252 21437 4261 21471
rect 4261 21437 4295 21471
rect 4295 21437 4304 21471
rect 4252 21428 4304 21437
rect 4712 21428 4764 21480
rect 4988 21428 5040 21480
rect 6000 21471 6052 21480
rect 6000 21437 6009 21471
rect 6009 21437 6043 21471
rect 6043 21437 6052 21471
rect 6000 21428 6052 21437
rect 6828 21428 6880 21480
rect 7564 21428 7616 21480
rect 8484 21428 8536 21480
rect 10692 21428 10744 21480
rect 12716 21564 12768 21616
rect 15200 21564 15252 21616
rect 17776 21632 17828 21684
rect 25412 21632 25464 21684
rect 29828 21632 29880 21684
rect 25136 21564 25188 21616
rect 25596 21564 25648 21616
rect 27988 21607 28040 21616
rect 27988 21573 27997 21607
rect 27997 21573 28031 21607
rect 28031 21573 28040 21607
rect 27988 21564 28040 21573
rect 14096 21496 14148 21548
rect 15108 21496 15160 21548
rect 16580 21496 16632 21548
rect 20904 21496 20956 21548
rect 23388 21539 23440 21548
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 26700 21496 26752 21548
rect 38292 21539 38344 21548
rect 38292 21505 38301 21539
rect 38301 21505 38335 21539
rect 38335 21505 38344 21539
rect 38292 21496 38344 21505
rect 2228 21292 2280 21344
rect 2504 21292 2556 21344
rect 4896 21292 4948 21344
rect 5724 21292 5776 21344
rect 11796 21360 11848 21412
rect 8668 21335 8720 21344
rect 8668 21301 8677 21335
rect 8677 21301 8711 21335
rect 8711 21301 8720 21335
rect 8668 21292 8720 21301
rect 8760 21292 8812 21344
rect 12348 21292 12400 21344
rect 19248 21428 19300 21480
rect 28080 21428 28132 21480
rect 18512 21292 18564 21344
rect 22008 21360 22060 21412
rect 26424 21360 26476 21412
rect 27804 21360 27856 21412
rect 19892 21292 19944 21344
rect 26332 21335 26384 21344
rect 26332 21301 26341 21335
rect 26341 21301 26375 21335
rect 26375 21301 26384 21335
rect 26332 21292 26384 21301
rect 29736 21292 29788 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 3148 20952 3200 21004
rect 4068 20816 4120 20868
rect 3332 20791 3384 20800
rect 3332 20757 3341 20791
rect 3341 20757 3375 20791
rect 3375 20757 3384 20791
rect 3332 20748 3384 20757
rect 6920 21088 6972 21140
rect 9864 21088 9916 21140
rect 14924 21088 14976 21140
rect 16396 21088 16448 21140
rect 17776 21088 17828 21140
rect 10416 20952 10468 21004
rect 17224 21020 17276 21072
rect 18512 21020 18564 21072
rect 22008 21020 22060 21072
rect 27068 21020 27120 21072
rect 15108 20952 15160 21004
rect 16212 20995 16264 21004
rect 16212 20961 16221 20995
rect 16221 20961 16255 20995
rect 16255 20961 16264 20995
rect 16212 20952 16264 20961
rect 19800 20952 19852 21004
rect 20720 20952 20772 21004
rect 21088 20952 21140 21004
rect 26976 20995 27028 21004
rect 6828 20927 6880 20936
rect 6828 20893 6837 20927
rect 6837 20893 6871 20927
rect 6871 20893 6880 20927
rect 6828 20884 6880 20893
rect 8944 20884 8996 20936
rect 9588 20884 9640 20936
rect 10508 20884 10560 20936
rect 10968 20927 11020 20936
rect 10968 20893 10977 20927
rect 10977 20893 11011 20927
rect 11011 20893 11020 20927
rect 10968 20884 11020 20893
rect 19248 20884 19300 20936
rect 7012 20816 7064 20868
rect 7380 20816 7432 20868
rect 8576 20816 8628 20868
rect 6276 20748 6328 20800
rect 6828 20748 6880 20800
rect 8484 20748 8536 20800
rect 11336 20748 11388 20800
rect 11704 20816 11756 20868
rect 19800 20859 19852 20868
rect 13820 20748 13872 20800
rect 14924 20748 14976 20800
rect 16212 20748 16264 20800
rect 19800 20825 19809 20859
rect 19809 20825 19843 20859
rect 19843 20825 19852 20859
rect 19800 20816 19852 20825
rect 19892 20859 19944 20868
rect 19892 20825 19901 20859
rect 19901 20825 19935 20859
rect 19935 20825 19944 20859
rect 19892 20816 19944 20825
rect 26976 20961 26985 20995
rect 26985 20961 27019 20995
rect 27019 20961 27028 20995
rect 26976 20952 27028 20961
rect 29552 20952 29604 21004
rect 23664 20927 23716 20936
rect 23664 20893 23673 20927
rect 23673 20893 23707 20927
rect 23707 20893 23716 20927
rect 23664 20884 23716 20893
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 37556 20884 37608 20936
rect 38292 20927 38344 20936
rect 38292 20893 38301 20927
rect 38301 20893 38335 20927
rect 38335 20893 38344 20927
rect 38292 20884 38344 20893
rect 25228 20816 25280 20868
rect 26424 20859 26476 20868
rect 26424 20825 26433 20859
rect 26433 20825 26467 20859
rect 26467 20825 26476 20859
rect 26424 20816 26476 20825
rect 28356 20859 28408 20868
rect 28356 20825 28365 20859
rect 28365 20825 28399 20859
rect 28399 20825 28408 20859
rect 28908 20859 28960 20868
rect 28356 20816 28408 20825
rect 28908 20825 28917 20859
rect 28917 20825 28951 20859
rect 28951 20825 28960 20859
rect 28908 20816 28960 20825
rect 25780 20748 25832 20800
rect 30472 20791 30524 20800
rect 30472 20757 30481 20791
rect 30481 20757 30515 20791
rect 30515 20757 30524 20791
rect 30472 20748 30524 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1952 20476 2004 20528
rect 6736 20476 6788 20528
rect 8484 20519 8536 20528
rect 8484 20485 8493 20519
rect 8493 20485 8527 20519
rect 8527 20485 8536 20519
rect 8484 20476 8536 20485
rect 1400 20408 1452 20460
rect 4620 20340 4672 20392
rect 3700 20272 3752 20324
rect 9680 20476 9732 20528
rect 10416 20476 10468 20528
rect 3148 20204 3200 20256
rect 4620 20204 4672 20256
rect 6644 20204 6696 20256
rect 7748 20204 7800 20256
rect 10140 20340 10192 20392
rect 10784 20544 10836 20596
rect 11888 20519 11940 20528
rect 11888 20485 11897 20519
rect 11897 20485 11931 20519
rect 11931 20485 11940 20519
rect 11888 20476 11940 20485
rect 12532 20476 12584 20528
rect 13728 20476 13780 20528
rect 14188 20476 14240 20528
rect 15108 20476 15160 20528
rect 18972 20476 19024 20528
rect 12072 20408 12124 20460
rect 12348 20408 12400 20460
rect 13268 20408 13320 20460
rect 16488 20408 16540 20460
rect 23664 20544 23716 20596
rect 22560 20476 22612 20528
rect 23756 20519 23808 20528
rect 23756 20485 23765 20519
rect 23765 20485 23799 20519
rect 23799 20485 23808 20519
rect 23756 20476 23808 20485
rect 25780 20519 25832 20528
rect 25780 20485 25789 20519
rect 25789 20485 25823 20519
rect 25823 20485 25832 20519
rect 25780 20476 25832 20485
rect 30472 20544 30524 20596
rect 10968 20340 11020 20392
rect 13728 20340 13780 20392
rect 21824 20408 21876 20460
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 24860 20408 24912 20460
rect 9772 20204 9824 20256
rect 10600 20204 10652 20256
rect 10876 20247 10928 20256
rect 10876 20213 10885 20247
rect 10885 20213 10919 20247
rect 10919 20213 10928 20247
rect 10876 20204 10928 20213
rect 13268 20272 13320 20324
rect 22192 20272 22244 20324
rect 16672 20204 16724 20256
rect 16764 20204 16816 20256
rect 20536 20204 20588 20256
rect 22100 20247 22152 20256
rect 22100 20213 22109 20247
rect 22109 20213 22143 20247
rect 22143 20213 22152 20247
rect 23480 20340 23532 20392
rect 24032 20383 24084 20392
rect 24032 20349 24041 20383
rect 24041 20349 24075 20383
rect 24075 20349 24084 20383
rect 24032 20340 24084 20349
rect 26148 20340 26200 20392
rect 27344 20408 27396 20460
rect 29000 20451 29052 20460
rect 29000 20417 29009 20451
rect 29009 20417 29043 20451
rect 29043 20417 29052 20451
rect 29000 20408 29052 20417
rect 26424 20272 26476 20324
rect 29552 20383 29604 20392
rect 29552 20349 29561 20383
rect 29561 20349 29595 20383
rect 29595 20349 29604 20383
rect 29552 20340 29604 20349
rect 30380 20383 30432 20392
rect 30380 20349 30389 20383
rect 30389 20349 30423 20383
rect 30423 20349 30432 20383
rect 30380 20340 30432 20349
rect 22100 20204 22152 20213
rect 29736 20204 29788 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2136 20000 2188 20052
rect 5724 19975 5776 19984
rect 5724 19941 5733 19975
rect 5733 19941 5767 19975
rect 5767 19941 5776 19975
rect 5724 19932 5776 19941
rect 3148 19864 3200 19916
rect 3976 19907 4028 19916
rect 3976 19873 3985 19907
rect 3985 19873 4019 19907
rect 4019 19873 4028 19907
rect 3976 19864 4028 19873
rect 5540 19864 5592 19916
rect 7012 19864 7064 19916
rect 7748 20000 7800 20052
rect 10692 20000 10744 20052
rect 15292 20000 15344 20052
rect 12256 19932 12308 19984
rect 10600 19907 10652 19916
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 10968 19864 11020 19916
rect 11888 19864 11940 19916
rect 15108 19864 15160 19916
rect 28264 20000 28316 20052
rect 21640 19932 21692 19984
rect 22652 19932 22704 19984
rect 24032 19932 24084 19984
rect 28908 19932 28960 19984
rect 16580 19907 16632 19916
rect 16580 19873 16589 19907
rect 16589 19873 16623 19907
rect 16623 19873 16632 19907
rect 16580 19864 16632 19873
rect 16948 19864 17000 19916
rect 20260 19864 20312 19916
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 20904 19907 20956 19916
rect 20904 19873 20913 19907
rect 20913 19873 20947 19907
rect 20947 19873 20956 19907
rect 20904 19864 20956 19873
rect 25688 19864 25740 19916
rect 26148 19907 26200 19916
rect 26148 19873 26157 19907
rect 26157 19873 26191 19907
rect 26191 19873 26200 19907
rect 26148 19864 26200 19873
rect 26608 19907 26660 19916
rect 26608 19873 26617 19907
rect 26617 19873 26651 19907
rect 26651 19873 26660 19907
rect 26608 19864 26660 19873
rect 20352 19839 20404 19848
rect 3240 19728 3292 19780
rect 3332 19728 3384 19780
rect 3608 19660 3660 19712
rect 4712 19728 4764 19780
rect 5172 19660 5224 19712
rect 11336 19728 11388 19780
rect 12256 19728 12308 19780
rect 20352 19805 20361 19839
rect 20361 19805 20395 19839
rect 20395 19805 20404 19839
rect 20352 19796 20404 19805
rect 24952 19839 25004 19848
rect 24952 19805 24961 19839
rect 24961 19805 24995 19839
rect 24995 19805 25004 19839
rect 24952 19796 25004 19805
rect 27436 19796 27488 19848
rect 28448 19796 28500 19848
rect 13176 19771 13228 19780
rect 13176 19737 13185 19771
rect 13185 19737 13219 19771
rect 13219 19737 13228 19771
rect 13176 19728 13228 19737
rect 16488 19728 16540 19780
rect 16948 19728 17000 19780
rect 19432 19728 19484 19780
rect 22744 19771 22796 19780
rect 22744 19737 22753 19771
rect 22753 19737 22787 19771
rect 22787 19737 22796 19771
rect 22744 19728 22796 19737
rect 22836 19771 22888 19780
rect 22836 19737 22845 19771
rect 22845 19737 22879 19771
rect 22879 19737 22888 19771
rect 22836 19728 22888 19737
rect 6828 19660 6880 19712
rect 7840 19660 7892 19712
rect 13728 19660 13780 19712
rect 17132 19660 17184 19712
rect 18328 19703 18380 19712
rect 18328 19669 18337 19703
rect 18337 19669 18371 19703
rect 18371 19669 18380 19703
rect 25044 19703 25096 19712
rect 18328 19660 18380 19669
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 26240 19771 26292 19780
rect 26240 19737 26249 19771
rect 26249 19737 26283 19771
rect 26283 19737 26292 19771
rect 26240 19728 26292 19737
rect 29644 19728 29696 19780
rect 27344 19660 27396 19712
rect 27804 19703 27856 19712
rect 27804 19669 27813 19703
rect 27813 19669 27847 19703
rect 27847 19669 27856 19703
rect 27804 19660 27856 19669
rect 29000 19660 29052 19712
rect 30564 19660 30616 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3700 19456 3752 19508
rect 4896 19456 4948 19508
rect 2872 19388 2924 19440
rect 7472 19456 7524 19508
rect 3976 19320 4028 19372
rect 5816 19320 5868 19372
rect 1676 19116 1728 19168
rect 6000 19252 6052 19304
rect 6460 19252 6512 19304
rect 9772 19456 9824 19508
rect 16672 19456 16724 19508
rect 8944 19388 8996 19440
rect 13636 19388 13688 19440
rect 16764 19388 16816 19440
rect 17776 19388 17828 19440
rect 19248 19456 19300 19508
rect 20352 19499 20404 19508
rect 20352 19465 20361 19499
rect 20361 19465 20395 19499
rect 20395 19465 20404 19499
rect 20352 19456 20404 19465
rect 27436 19456 27488 19508
rect 23112 19431 23164 19440
rect 23112 19397 23121 19431
rect 23121 19397 23155 19431
rect 23155 19397 23164 19431
rect 23112 19388 23164 19397
rect 24768 19388 24820 19440
rect 29000 19431 29052 19440
rect 29000 19397 29009 19431
rect 29009 19397 29043 19431
rect 29043 19397 29052 19431
rect 29000 19388 29052 19397
rect 30380 19456 30432 19508
rect 37648 19456 37700 19508
rect 30564 19431 30616 19440
rect 30564 19397 30573 19431
rect 30573 19397 30607 19431
rect 30607 19397 30616 19431
rect 30564 19388 30616 19397
rect 6000 19116 6052 19168
rect 11060 19252 11112 19304
rect 12164 19295 12216 19304
rect 12164 19261 12173 19295
rect 12173 19261 12207 19295
rect 12207 19261 12216 19295
rect 12164 19252 12216 19261
rect 13728 19320 13780 19372
rect 14096 19363 14148 19372
rect 14096 19329 14105 19363
rect 14105 19329 14139 19363
rect 14139 19329 14148 19363
rect 14096 19320 14148 19329
rect 16580 19320 16632 19372
rect 18880 19320 18932 19372
rect 13820 19116 13872 19168
rect 14372 19116 14424 19168
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 18696 19252 18748 19304
rect 20260 19320 20312 19372
rect 23848 19320 23900 19372
rect 24032 19320 24084 19372
rect 28080 19320 28132 19372
rect 38292 19363 38344 19372
rect 38292 19329 38301 19363
rect 38301 19329 38335 19363
rect 38335 19329 38344 19363
rect 38292 19320 38344 19329
rect 28908 19295 28960 19304
rect 28908 19261 28917 19295
rect 28917 19261 28951 19295
rect 28951 19261 28960 19295
rect 28908 19252 28960 19261
rect 30472 19295 30524 19304
rect 30472 19261 30481 19295
rect 30481 19261 30515 19295
rect 30515 19261 30524 19295
rect 30472 19252 30524 19261
rect 28816 19184 28868 19236
rect 18328 19116 18380 19168
rect 22468 19116 22520 19168
rect 30104 19116 30156 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 6552 18912 6604 18964
rect 9956 18912 10008 18964
rect 10048 18912 10100 18964
rect 12532 18912 12584 18964
rect 13544 18912 13596 18964
rect 15016 18912 15068 18964
rect 19432 18912 19484 18964
rect 22744 18955 22796 18964
rect 22744 18921 22753 18955
rect 22753 18921 22787 18955
rect 22787 18921 22796 18955
rect 22744 18912 22796 18921
rect 23112 18912 23164 18964
rect 30104 18955 30156 18964
rect 3424 18776 3476 18828
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 3056 18708 3108 18760
rect 6828 18751 6880 18760
rect 6828 18717 6837 18751
rect 6837 18717 6871 18751
rect 6871 18717 6880 18751
rect 6828 18708 6880 18717
rect 8208 18708 8260 18760
rect 11336 18819 11388 18828
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11336 18776 11388 18785
rect 14096 18776 14148 18828
rect 20812 18776 20864 18828
rect 8668 18708 8720 18760
rect 11060 18751 11112 18760
rect 11060 18717 11069 18751
rect 11069 18717 11103 18751
rect 11103 18717 11112 18751
rect 11060 18708 11112 18717
rect 16396 18708 16448 18760
rect 4620 18572 4672 18624
rect 5632 18640 5684 18692
rect 11796 18640 11848 18692
rect 15016 18683 15068 18692
rect 15016 18649 15025 18683
rect 15025 18649 15059 18683
rect 15059 18649 15068 18683
rect 15016 18640 15068 18649
rect 15108 18640 15160 18692
rect 19340 18708 19392 18760
rect 19984 18708 20036 18760
rect 21640 18640 21692 18692
rect 5264 18572 5316 18624
rect 5540 18572 5592 18624
rect 6368 18615 6420 18624
rect 6368 18581 6377 18615
rect 6377 18581 6411 18615
rect 6411 18581 6420 18615
rect 6368 18572 6420 18581
rect 6460 18572 6512 18624
rect 9864 18572 9916 18624
rect 13544 18572 13596 18624
rect 18512 18572 18564 18624
rect 22928 18572 22980 18624
rect 30104 18921 30113 18955
rect 30113 18921 30147 18955
rect 30147 18921 30156 18955
rect 30104 18912 30156 18921
rect 25228 18887 25280 18896
rect 25228 18853 25237 18887
rect 25237 18853 25271 18887
rect 25271 18853 25280 18887
rect 25228 18844 25280 18853
rect 37924 18708 37976 18760
rect 25136 18572 25188 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1676 18368 1728 18420
rect 3976 18368 4028 18420
rect 5264 18368 5316 18420
rect 6000 18411 6052 18420
rect 3332 18300 3384 18352
rect 3700 18300 3752 18352
rect 3976 18232 4028 18284
rect 4160 18164 4212 18216
rect 4896 18164 4948 18216
rect 5264 18164 5316 18216
rect 6000 18377 6009 18411
rect 6009 18377 6043 18411
rect 6043 18377 6052 18411
rect 6000 18368 6052 18377
rect 8944 18368 8996 18420
rect 11704 18368 11756 18420
rect 13728 18368 13780 18420
rect 15292 18411 15344 18420
rect 7104 18300 7156 18352
rect 7472 18300 7524 18352
rect 8300 18300 8352 18352
rect 9956 18300 10008 18352
rect 6092 18232 6144 18284
rect 6552 18275 6604 18284
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 9220 18232 9272 18284
rect 6460 18096 6512 18148
rect 6828 18164 6880 18216
rect 7288 18207 7340 18216
rect 7288 18173 7297 18207
rect 7297 18173 7331 18207
rect 7331 18173 7340 18207
rect 7288 18164 7340 18173
rect 7656 18164 7708 18216
rect 10048 18164 10100 18216
rect 12624 18232 12676 18284
rect 14096 18300 14148 18352
rect 15292 18377 15301 18411
rect 15301 18377 15335 18411
rect 15335 18377 15344 18411
rect 15292 18368 15344 18377
rect 18604 18411 18656 18420
rect 18604 18377 18613 18411
rect 18613 18377 18647 18411
rect 18647 18377 18656 18411
rect 18604 18368 18656 18377
rect 18972 18368 19024 18420
rect 17224 18300 17276 18352
rect 18420 18300 18472 18352
rect 16580 18232 16632 18284
rect 13820 18207 13872 18216
rect 11152 18028 11204 18080
rect 11336 18028 11388 18080
rect 13544 18028 13596 18080
rect 13820 18173 13829 18207
rect 13829 18173 13863 18207
rect 13863 18173 13872 18207
rect 13820 18164 13872 18173
rect 22744 18368 22796 18420
rect 24032 18368 24084 18420
rect 36636 18368 36688 18420
rect 20812 18300 20864 18352
rect 21732 18300 21784 18352
rect 21916 18232 21968 18284
rect 22100 18232 22152 18284
rect 24492 18275 24544 18284
rect 24492 18241 24501 18275
rect 24501 18241 24535 18275
rect 24535 18241 24544 18275
rect 24492 18232 24544 18241
rect 38292 18275 38344 18284
rect 38292 18241 38301 18275
rect 38301 18241 38335 18275
rect 38335 18241 38344 18275
rect 38292 18232 38344 18241
rect 19800 18028 19852 18080
rect 21364 18028 21416 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4252 17824 4304 17876
rect 4804 17824 4856 17876
rect 7012 17824 7064 17876
rect 9680 17824 9732 17876
rect 10784 17824 10836 17876
rect 3976 17731 4028 17740
rect 3976 17697 3985 17731
rect 3985 17697 4019 17731
rect 4019 17697 4028 17731
rect 3976 17688 4028 17697
rect 4620 17688 4672 17740
rect 7288 17688 7340 17740
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 15016 17824 15068 17876
rect 1768 17663 1820 17672
rect 1768 17629 1777 17663
rect 1777 17629 1811 17663
rect 1811 17629 1820 17663
rect 1768 17620 1820 17629
rect 2228 17663 2280 17672
rect 2228 17629 2237 17663
rect 2237 17629 2271 17663
rect 2271 17629 2280 17663
rect 2228 17620 2280 17629
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 1768 17484 1820 17536
rect 2044 17484 2096 17536
rect 4160 17484 4212 17536
rect 4896 17552 4948 17604
rect 5816 17552 5868 17604
rect 6460 17484 6512 17536
rect 7104 17552 7156 17604
rect 10508 17552 10560 17604
rect 12716 17552 12768 17604
rect 17040 17824 17092 17876
rect 22744 17824 22796 17876
rect 17592 17756 17644 17808
rect 24860 17756 24912 17808
rect 16580 17688 16632 17740
rect 19800 17731 19852 17740
rect 19800 17697 19809 17731
rect 19809 17697 19843 17731
rect 19843 17697 19852 17731
rect 19800 17688 19852 17697
rect 20812 17731 20864 17740
rect 20812 17697 20821 17731
rect 20821 17697 20855 17731
rect 20855 17697 20864 17731
rect 20812 17688 20864 17697
rect 21364 17688 21416 17740
rect 18052 17620 18104 17672
rect 19340 17620 19392 17672
rect 19432 17620 19484 17672
rect 23020 17620 23072 17672
rect 7564 17484 7616 17536
rect 10692 17484 10744 17536
rect 16672 17552 16724 17604
rect 20812 17552 20864 17604
rect 24032 17552 24084 17604
rect 37280 17552 37332 17604
rect 13820 17484 13872 17536
rect 14832 17484 14884 17536
rect 15200 17484 15252 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1584 17280 1636 17332
rect 7104 17280 7156 17332
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 2964 17144 3016 17196
rect 3792 17212 3844 17264
rect 4068 17212 4120 17264
rect 3424 17144 3476 17196
rect 3516 17076 3568 17128
rect 4252 17144 4304 17196
rect 5356 17212 5408 17264
rect 6552 17212 6604 17264
rect 5448 17187 5500 17196
rect 5448 17153 5457 17187
rect 5457 17153 5491 17187
rect 5491 17153 5500 17187
rect 5448 17144 5500 17153
rect 5540 17144 5592 17196
rect 7932 17144 7984 17196
rect 11060 17280 11112 17332
rect 11980 17280 12032 17332
rect 14188 17280 14240 17332
rect 17776 17323 17828 17332
rect 17776 17289 17785 17323
rect 17785 17289 17819 17323
rect 17819 17289 17828 17323
rect 17776 17280 17828 17289
rect 18420 17323 18472 17332
rect 18420 17289 18429 17323
rect 18429 17289 18463 17323
rect 18463 17289 18472 17323
rect 18420 17280 18472 17289
rect 19432 17280 19484 17332
rect 23112 17280 23164 17332
rect 28908 17280 28960 17332
rect 9680 17212 9732 17264
rect 11888 17255 11940 17264
rect 11888 17221 11897 17255
rect 11897 17221 11931 17255
rect 11931 17221 11940 17255
rect 11888 17212 11940 17221
rect 10968 17144 11020 17196
rect 8392 17076 8444 17128
rect 9772 17076 9824 17128
rect 10876 17076 10928 17128
rect 11060 17076 11112 17128
rect 13176 17076 13228 17128
rect 15936 17144 15988 17196
rect 16488 17144 16540 17196
rect 18052 17144 18104 17196
rect 18144 17144 18196 17196
rect 18420 17144 18472 17196
rect 37556 17212 37608 17264
rect 15292 17076 15344 17128
rect 37740 17144 37792 17196
rect 2596 17008 2648 17060
rect 1492 16940 1544 16992
rect 8484 17008 8536 17060
rect 3792 16983 3844 16992
rect 3792 16949 3801 16983
rect 3801 16949 3835 16983
rect 3835 16949 3844 16983
rect 3792 16940 3844 16949
rect 6644 16940 6696 16992
rect 10140 16940 10192 16992
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 15016 17008 15068 17060
rect 22376 17008 22428 17060
rect 11152 16940 11204 16949
rect 15200 16940 15252 16992
rect 17040 16940 17092 16992
rect 19156 16940 19208 16992
rect 37832 16940 37884 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3516 16736 3568 16788
rect 6184 16736 6236 16788
rect 6552 16736 6604 16788
rect 9588 16736 9640 16788
rect 1676 16532 1728 16584
rect 2964 16600 3016 16652
rect 1768 16464 1820 16516
rect 3976 16532 4028 16584
rect 6092 16668 6144 16720
rect 6276 16668 6328 16720
rect 3424 16464 3476 16516
rect 3700 16464 3752 16516
rect 1952 16396 2004 16448
rect 5632 16600 5684 16652
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 5540 16532 5592 16584
rect 5908 16532 5960 16584
rect 6092 16532 6144 16584
rect 8116 16600 8168 16652
rect 8392 16600 8444 16652
rect 17592 16736 17644 16788
rect 8760 16464 8812 16516
rect 10692 16575 10744 16584
rect 10692 16541 10701 16575
rect 10701 16541 10735 16575
rect 10735 16541 10744 16575
rect 10692 16532 10744 16541
rect 12532 16668 12584 16720
rect 12624 16668 12676 16720
rect 12348 16600 12400 16652
rect 13636 16575 13688 16584
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 14832 16668 14884 16720
rect 25136 16736 25188 16788
rect 13636 16532 13688 16541
rect 15108 16532 15160 16584
rect 15292 16532 15344 16584
rect 16948 16600 17000 16652
rect 18696 16532 18748 16584
rect 22100 16532 22152 16584
rect 16856 16464 16908 16516
rect 17500 16507 17552 16516
rect 17500 16473 17509 16507
rect 17509 16473 17543 16507
rect 17543 16473 17552 16507
rect 17500 16464 17552 16473
rect 19340 16464 19392 16516
rect 20076 16464 20128 16516
rect 26516 16532 26568 16584
rect 37924 16532 37976 16584
rect 5724 16396 5776 16448
rect 5908 16439 5960 16448
rect 5908 16405 5917 16439
rect 5917 16405 5951 16439
rect 5951 16405 5960 16439
rect 5908 16396 5960 16405
rect 6920 16396 6972 16448
rect 7656 16396 7708 16448
rect 10140 16396 10192 16448
rect 11520 16396 11572 16448
rect 11704 16439 11756 16448
rect 11704 16405 11713 16439
rect 11713 16405 11747 16439
rect 11747 16405 11756 16439
rect 11704 16396 11756 16405
rect 16304 16396 16356 16448
rect 16764 16439 16816 16448
rect 16764 16405 16773 16439
rect 16773 16405 16807 16439
rect 16807 16405 16816 16439
rect 16764 16396 16816 16405
rect 22652 16396 22704 16448
rect 22744 16396 22796 16448
rect 23204 16464 23256 16516
rect 38108 16507 38160 16516
rect 38108 16473 38117 16507
rect 38117 16473 38151 16507
rect 38151 16473 38160 16507
rect 38108 16464 38160 16473
rect 37924 16396 37976 16448
rect 38200 16439 38252 16448
rect 38200 16405 38209 16439
rect 38209 16405 38243 16439
rect 38243 16405 38252 16439
rect 38200 16396 38252 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 3332 16235 3384 16244
rect 3332 16201 3341 16235
rect 3341 16201 3375 16235
rect 3375 16201 3384 16235
rect 3332 16192 3384 16201
rect 3424 16192 3476 16244
rect 4160 16167 4212 16176
rect 4160 16133 4169 16167
rect 4169 16133 4203 16167
rect 4203 16133 4212 16167
rect 4160 16124 4212 16133
rect 5908 16124 5960 16176
rect 2596 16099 2648 16108
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 2964 16056 3016 16108
rect 7196 16192 7248 16244
rect 8208 16235 8260 16244
rect 8208 16201 8217 16235
rect 8217 16201 8251 16235
rect 8251 16201 8260 16235
rect 8208 16192 8260 16201
rect 9680 16192 9732 16244
rect 10416 16235 10468 16244
rect 10416 16201 10425 16235
rect 10425 16201 10459 16235
rect 10459 16201 10468 16235
rect 10416 16192 10468 16201
rect 11244 16192 11296 16244
rect 13728 16235 13780 16244
rect 13728 16201 13737 16235
rect 13737 16201 13771 16235
rect 13771 16201 13780 16235
rect 13728 16192 13780 16201
rect 17500 16192 17552 16244
rect 19340 16192 19392 16244
rect 22100 16192 22152 16244
rect 22560 16192 22612 16244
rect 24584 16192 24636 16244
rect 37740 16192 37792 16244
rect 11888 16167 11940 16176
rect 6092 16056 6144 16108
rect 8760 16099 8812 16108
rect 8760 16065 8769 16099
rect 8769 16065 8803 16099
rect 8803 16065 8812 16099
rect 8760 16056 8812 16065
rect 9680 16099 9732 16108
rect 9680 16065 9689 16099
rect 9689 16065 9723 16099
rect 9723 16065 9732 16099
rect 9680 16056 9732 16065
rect 11888 16133 11897 16167
rect 11897 16133 11931 16167
rect 11931 16133 11940 16167
rect 11888 16124 11940 16133
rect 12624 16167 12676 16176
rect 12624 16133 12633 16167
rect 12633 16133 12667 16167
rect 12667 16133 12676 16167
rect 12624 16124 12676 16133
rect 17040 16167 17092 16176
rect 17040 16133 17049 16167
rect 17049 16133 17083 16167
rect 17083 16133 17092 16167
rect 17040 16124 17092 16133
rect 19156 16167 19208 16176
rect 19156 16133 19165 16167
rect 19165 16133 19199 16167
rect 19199 16133 19208 16167
rect 19156 16124 19208 16133
rect 20628 16124 20680 16176
rect 22468 16124 22520 16176
rect 22928 16124 22980 16176
rect 23296 16124 23348 16176
rect 11060 16056 11112 16108
rect 11612 16056 11664 16108
rect 13176 16056 13228 16108
rect 16304 16099 16356 16108
rect 16304 16065 16313 16099
rect 16313 16065 16347 16099
rect 16347 16065 16356 16099
rect 16304 16056 16356 16065
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 4712 15988 4764 16040
rect 5448 15988 5500 16040
rect 8300 15988 8352 16040
rect 8392 15988 8444 16040
rect 7196 15920 7248 15972
rect 10692 15920 10744 15972
rect 11612 15920 11664 15972
rect 18328 15988 18380 16040
rect 18880 15988 18932 16040
rect 19340 16031 19392 16040
rect 19340 15997 19349 16031
rect 19349 15997 19383 16031
rect 19383 15997 19392 16031
rect 19340 15988 19392 15997
rect 20076 15920 20128 15972
rect 20628 15988 20680 16040
rect 23572 16031 23624 16040
rect 21916 15920 21968 15972
rect 23572 15997 23581 16031
rect 23581 15997 23615 16031
rect 23615 15997 23624 16031
rect 23572 15988 23624 15997
rect 26148 15988 26200 16040
rect 37648 16056 37700 16108
rect 38292 16099 38344 16108
rect 38292 16065 38301 16099
rect 38301 16065 38335 16099
rect 38335 16065 38344 16099
rect 38292 16056 38344 16065
rect 36544 15988 36596 16040
rect 23480 15920 23532 15972
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 2596 15852 2648 15904
rect 5356 15852 5408 15904
rect 5540 15852 5592 15904
rect 6092 15852 6144 15904
rect 9680 15852 9732 15904
rect 10232 15852 10284 15904
rect 12072 15852 12124 15904
rect 18788 15852 18840 15904
rect 19340 15852 19392 15904
rect 20628 15852 20680 15904
rect 22928 15852 22980 15904
rect 23112 15852 23164 15904
rect 26424 15920 26476 15972
rect 24860 15852 24912 15904
rect 33324 15895 33376 15904
rect 33324 15861 33333 15895
rect 33333 15861 33367 15895
rect 33367 15861 33376 15895
rect 33324 15852 33376 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8392 15648 8444 15700
rect 10508 15648 10560 15700
rect 3148 15623 3200 15632
rect 3148 15589 3157 15623
rect 3157 15589 3191 15623
rect 3191 15589 3200 15623
rect 3148 15580 3200 15589
rect 16580 15648 16632 15700
rect 18788 15648 18840 15700
rect 22008 15648 22060 15700
rect 22560 15648 22612 15700
rect 22652 15648 22704 15700
rect 10692 15580 10744 15632
rect 12256 15580 12308 15632
rect 13176 15580 13228 15632
rect 20628 15580 20680 15632
rect 23112 15512 23164 15564
rect 26148 15555 26200 15564
rect 26148 15521 26157 15555
rect 26157 15521 26191 15555
rect 26191 15521 26200 15555
rect 26148 15512 26200 15521
rect 34796 15580 34848 15632
rect 27896 15555 27948 15564
rect 27896 15521 27905 15555
rect 27905 15521 27939 15555
rect 27939 15521 27948 15555
rect 27896 15512 27948 15521
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 9680 15444 9732 15496
rect 1768 15351 1820 15360
rect 1768 15317 1777 15351
rect 1777 15317 1811 15351
rect 1811 15317 1820 15351
rect 1768 15308 1820 15317
rect 4160 15376 4212 15428
rect 5264 15376 5316 15428
rect 5356 15419 5408 15428
rect 5356 15385 5365 15419
rect 5365 15385 5399 15419
rect 5399 15385 5408 15419
rect 5356 15376 5408 15385
rect 7012 15376 7064 15428
rect 7656 15419 7708 15428
rect 7656 15385 7665 15419
rect 7665 15385 7699 15419
rect 7699 15385 7708 15419
rect 8576 15419 8628 15428
rect 7656 15376 7708 15385
rect 8576 15385 8585 15419
rect 8585 15385 8619 15419
rect 8619 15385 8628 15419
rect 8576 15376 8628 15385
rect 10048 15419 10100 15428
rect 10048 15385 10057 15419
rect 10057 15385 10091 15419
rect 10091 15385 10100 15419
rect 10048 15376 10100 15385
rect 10140 15419 10192 15428
rect 10140 15385 10149 15419
rect 10149 15385 10183 15419
rect 10183 15385 10192 15419
rect 10140 15376 10192 15385
rect 8024 15308 8076 15360
rect 9864 15308 9916 15360
rect 10416 15308 10468 15360
rect 11520 15419 11572 15428
rect 11520 15385 11529 15419
rect 11529 15385 11563 15419
rect 11563 15385 11572 15419
rect 11520 15376 11572 15385
rect 11888 15376 11940 15428
rect 13176 15487 13228 15496
rect 13176 15453 13185 15487
rect 13185 15453 13219 15487
rect 13219 15453 13228 15487
rect 13176 15444 13228 15453
rect 18052 15444 18104 15496
rect 12348 15376 12400 15428
rect 15660 15376 15712 15428
rect 16856 15419 16908 15428
rect 16856 15385 16865 15419
rect 16865 15385 16899 15419
rect 16899 15385 16908 15419
rect 16856 15376 16908 15385
rect 17868 15419 17920 15428
rect 11612 15308 11664 15360
rect 11704 15308 11756 15360
rect 17868 15385 17877 15419
rect 17877 15385 17911 15419
rect 17911 15385 17920 15419
rect 17868 15376 17920 15385
rect 20260 15444 20312 15496
rect 20996 15444 21048 15496
rect 22468 15444 22520 15496
rect 21364 15376 21416 15428
rect 19432 15308 19484 15360
rect 22008 15308 22060 15360
rect 22928 15419 22980 15428
rect 22928 15385 22937 15419
rect 22937 15385 22971 15419
rect 22971 15385 22980 15419
rect 22928 15376 22980 15385
rect 23112 15376 23164 15428
rect 25044 15376 25096 15428
rect 26056 15376 26108 15428
rect 29828 15419 29880 15428
rect 29828 15385 29837 15419
rect 29837 15385 29871 15419
rect 29871 15385 29880 15419
rect 29828 15376 29880 15385
rect 23480 15308 23532 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 5356 15104 5408 15156
rect 3792 15036 3844 15088
rect 5724 15036 5776 15088
rect 6828 15036 6880 15088
rect 8300 15036 8352 15088
rect 10232 15079 10284 15088
rect 10232 15045 10241 15079
rect 10241 15045 10275 15079
rect 10275 15045 10284 15079
rect 10232 15036 10284 15045
rect 7288 15011 7340 15018
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 7288 14966 7340 14977
rect 7656 14968 7708 15020
rect 9772 14968 9824 15020
rect 3332 14900 3384 14952
rect 3700 14943 3752 14952
rect 3700 14909 3709 14943
rect 3709 14909 3743 14943
rect 3743 14909 3752 14943
rect 3700 14900 3752 14909
rect 1952 14832 2004 14884
rect 5908 14900 5960 14952
rect 6828 14832 6880 14884
rect 8208 14900 8260 14952
rect 8484 14900 8536 14952
rect 9864 14832 9916 14884
rect 10232 14900 10284 14952
rect 11704 15104 11756 15156
rect 12716 15104 12768 15156
rect 16580 15104 16632 15156
rect 11428 15036 11480 15088
rect 16212 15036 16264 15088
rect 16764 15036 16816 15088
rect 17960 15104 18012 15156
rect 21824 15036 21876 15088
rect 22100 15036 22152 15088
rect 23572 15036 23624 15088
rect 24584 15036 24636 15088
rect 11888 14968 11940 15020
rect 12256 14968 12308 15020
rect 14004 14968 14056 15020
rect 16672 14968 16724 15020
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 18788 14968 18840 15020
rect 21364 14968 21416 15020
rect 11980 14900 12032 14952
rect 16580 14900 16632 14952
rect 17224 14943 17276 14952
rect 17224 14909 17233 14943
rect 17233 14909 17267 14943
rect 17267 14909 17276 14943
rect 17224 14900 17276 14909
rect 17592 14900 17644 14952
rect 20904 14900 20956 14952
rect 21916 14900 21968 14952
rect 11888 14832 11940 14884
rect 15016 14832 15068 14884
rect 20996 14832 21048 14884
rect 22928 14900 22980 14952
rect 24860 14900 24912 14952
rect 27712 14900 27764 14952
rect 27988 14900 28040 14952
rect 24308 14875 24360 14884
rect 24308 14841 24317 14875
rect 24317 14841 24351 14875
rect 24351 14841 24360 14875
rect 24308 14832 24360 14841
rect 26884 14832 26936 14884
rect 33600 14832 33652 14884
rect 8116 14807 8168 14816
rect 8116 14773 8125 14807
rect 8125 14773 8159 14807
rect 8159 14773 8168 14807
rect 8116 14764 8168 14773
rect 9404 14764 9456 14816
rect 18328 14764 18380 14816
rect 18420 14764 18472 14816
rect 18696 14764 18748 14816
rect 20168 14764 20220 14816
rect 20628 14764 20680 14816
rect 27712 14764 27764 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2872 14560 2924 14612
rect 3148 14560 3200 14612
rect 4068 14560 4120 14612
rect 5264 14560 5316 14612
rect 5908 14560 5960 14612
rect 6552 14560 6604 14612
rect 7932 14560 7984 14612
rect 8208 14603 8260 14612
rect 8208 14569 8217 14603
rect 8217 14569 8251 14603
rect 8251 14569 8260 14603
rect 8208 14560 8260 14569
rect 11796 14560 11848 14612
rect 16856 14560 16908 14612
rect 17684 14560 17736 14612
rect 24124 14560 24176 14612
rect 24584 14603 24636 14612
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 36544 14560 36596 14612
rect 3700 14492 3752 14544
rect 1676 14356 1728 14408
rect 2412 14399 2464 14408
rect 2412 14365 2421 14399
rect 2421 14365 2455 14399
rect 2455 14365 2464 14399
rect 2412 14356 2464 14365
rect 3792 14356 3844 14408
rect 3884 14356 3936 14408
rect 4804 14288 4856 14340
rect 5632 14356 5684 14408
rect 7380 14424 7432 14476
rect 12532 14424 12584 14476
rect 13268 14492 13320 14544
rect 19248 14492 19300 14544
rect 23664 14492 23716 14544
rect 17592 14424 17644 14476
rect 17868 14424 17920 14476
rect 7656 14356 7708 14408
rect 11060 14356 11112 14408
rect 11704 14356 11756 14408
rect 6552 14288 6604 14340
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 6920 14288 6972 14340
rect 7380 14331 7432 14340
rect 7380 14297 7389 14331
rect 7389 14297 7423 14331
rect 7423 14297 7432 14331
rect 7380 14288 7432 14297
rect 9404 14331 9456 14340
rect 9404 14297 9413 14331
rect 9413 14297 9447 14331
rect 9447 14297 9456 14331
rect 9404 14288 9456 14297
rect 10232 14288 10284 14340
rect 12348 14356 12400 14408
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 11888 14263 11940 14272
rect 11888 14229 11897 14263
rect 11897 14229 11931 14263
rect 11931 14229 11940 14263
rect 11888 14220 11940 14229
rect 11980 14220 12032 14272
rect 15292 14288 15344 14340
rect 17684 14288 17736 14340
rect 18696 14288 18748 14340
rect 19156 14288 19208 14340
rect 20996 14424 21048 14476
rect 29828 14424 29880 14476
rect 20904 14356 20956 14408
rect 21640 14356 21692 14408
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 24400 14356 24452 14408
rect 38292 14399 38344 14408
rect 38292 14365 38301 14399
rect 38301 14365 38335 14399
rect 38335 14365 38344 14399
rect 38292 14356 38344 14365
rect 19340 14220 19392 14272
rect 19432 14220 19484 14272
rect 23572 14288 23624 14340
rect 23388 14220 23440 14272
rect 27620 14263 27672 14272
rect 27620 14229 27629 14263
rect 27629 14229 27663 14263
rect 27663 14229 27672 14263
rect 27620 14220 27672 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4160 14016 4212 14068
rect 5356 14016 5408 14068
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 8116 14016 8168 14068
rect 9864 14016 9916 14068
rect 4712 13948 4764 14000
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 4068 13880 4120 13932
rect 5172 13880 5224 13932
rect 5724 13923 5776 13932
rect 2596 13812 2648 13864
rect 4160 13812 4212 13864
rect 4712 13812 4764 13864
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 6000 13880 6052 13932
rect 5356 13812 5408 13864
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 7104 13880 7156 13932
rect 6828 13812 6880 13821
rect 7656 13812 7708 13864
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 8024 13812 8076 13864
rect 5448 13744 5500 13796
rect 8392 13812 8444 13864
rect 9956 13880 10008 13932
rect 10784 13880 10836 13932
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 11336 13880 11388 13932
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 13820 13948 13872 14000
rect 16212 14016 16264 14068
rect 17132 13948 17184 14000
rect 18420 13991 18472 14000
rect 18420 13957 18429 13991
rect 18429 13957 18463 13991
rect 18463 13957 18472 13991
rect 18420 13948 18472 13957
rect 19248 13948 19300 14000
rect 19892 13948 19944 14000
rect 14004 13880 14056 13932
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 5080 13719 5132 13728
rect 5080 13685 5089 13719
rect 5089 13685 5123 13719
rect 5123 13685 5132 13719
rect 5080 13676 5132 13685
rect 6828 13676 6880 13728
rect 11888 13812 11940 13864
rect 12808 13812 12860 13864
rect 13728 13812 13780 13864
rect 15016 13812 15068 13864
rect 15292 13855 15344 13864
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 17868 13880 17920 13932
rect 20720 14016 20772 14068
rect 24400 14059 24452 14068
rect 24400 14025 24409 14059
rect 24409 14025 24443 14059
rect 24443 14025 24452 14059
rect 24400 14016 24452 14025
rect 26884 13948 26936 14000
rect 27620 13991 27672 14000
rect 27620 13957 27629 13991
rect 27629 13957 27663 13991
rect 27663 13957 27672 13991
rect 27620 13948 27672 13957
rect 27712 13991 27764 14000
rect 27712 13957 27721 13991
rect 27721 13957 27755 13991
rect 27755 13957 27764 13991
rect 27712 13948 27764 13957
rect 16488 13812 16540 13864
rect 19156 13812 19208 13864
rect 19892 13812 19944 13864
rect 22468 13880 22520 13932
rect 24584 13923 24636 13932
rect 24584 13889 24593 13923
rect 24593 13889 24627 13923
rect 24627 13889 24636 13923
rect 24584 13880 24636 13889
rect 26148 13812 26200 13864
rect 27712 13812 27764 13864
rect 27988 13855 28040 13864
rect 27988 13821 27997 13855
rect 27997 13821 28031 13855
rect 28031 13821 28040 13855
rect 27988 13812 28040 13821
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 9772 13676 9824 13685
rect 11244 13744 11296 13796
rect 12164 13744 12216 13796
rect 17960 13744 18012 13796
rect 18052 13744 18104 13796
rect 13360 13719 13412 13728
rect 13360 13685 13369 13719
rect 13369 13685 13403 13719
rect 13403 13685 13412 13719
rect 13360 13676 13412 13685
rect 15660 13676 15712 13728
rect 22284 13676 22336 13728
rect 38200 13676 38252 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2964 13472 3016 13524
rect 6736 13472 6788 13524
rect 7196 13472 7248 13524
rect 12348 13472 12400 13524
rect 12716 13472 12768 13524
rect 13820 13472 13872 13524
rect 2412 13336 2464 13388
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 3424 13379 3476 13388
rect 2780 13336 2832 13345
rect 3424 13345 3433 13379
rect 3433 13345 3467 13379
rect 3467 13345 3476 13379
rect 3424 13336 3476 13345
rect 7288 13404 7340 13456
rect 17224 13472 17276 13524
rect 30380 13472 30432 13524
rect 30564 13472 30616 13524
rect 7012 13379 7064 13388
rect 7012 13345 7021 13379
rect 7021 13345 7055 13379
rect 7055 13345 7064 13379
rect 7012 13336 7064 13345
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 10508 13336 10560 13388
rect 17040 13404 17092 13456
rect 18052 13404 18104 13456
rect 23204 13404 23256 13456
rect 26332 13404 26384 13456
rect 4620 13268 4672 13320
rect 5080 13268 5132 13320
rect 8392 13311 8444 13320
rect 2964 13132 3016 13184
rect 4620 13175 4672 13184
rect 4620 13141 4629 13175
rect 4629 13141 4663 13175
rect 4663 13141 4672 13175
rect 4620 13132 4672 13141
rect 6092 13175 6144 13184
rect 6092 13141 6101 13175
rect 6101 13141 6135 13175
rect 6135 13141 6144 13175
rect 6092 13132 6144 13141
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 6828 13243 6880 13252
rect 6828 13209 6837 13243
rect 6837 13209 6871 13243
rect 6871 13209 6880 13243
rect 6828 13200 6880 13209
rect 9772 13243 9824 13252
rect 9772 13209 9781 13243
rect 9781 13209 9815 13243
rect 9815 13209 9824 13243
rect 9772 13200 9824 13209
rect 9956 13200 10008 13252
rect 10692 13200 10744 13252
rect 12164 13268 12216 13320
rect 15936 13336 15988 13388
rect 16672 13379 16724 13388
rect 16672 13345 16681 13379
rect 16681 13345 16715 13379
rect 16715 13345 16724 13379
rect 16672 13336 16724 13345
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 14648 13268 14700 13320
rect 15660 13311 15712 13320
rect 15660 13277 15669 13311
rect 15669 13277 15703 13311
rect 15703 13277 15712 13311
rect 15660 13268 15712 13277
rect 17040 13268 17092 13320
rect 30472 13336 30524 13388
rect 30564 13379 30616 13388
rect 30564 13345 30573 13379
rect 30573 13345 30607 13379
rect 30607 13345 30616 13379
rect 30564 13336 30616 13345
rect 21456 13268 21508 13320
rect 37280 13311 37332 13320
rect 37280 13277 37289 13311
rect 37289 13277 37323 13311
rect 37323 13277 37332 13311
rect 37280 13268 37332 13277
rect 13268 13200 13320 13252
rect 14740 13200 14792 13252
rect 7472 13132 7524 13184
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 8668 13132 8720 13184
rect 12348 13132 12400 13184
rect 17316 13200 17368 13252
rect 20352 13200 20404 13252
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 17684 13132 17736 13184
rect 20812 13132 20864 13184
rect 23388 13243 23440 13252
rect 23388 13209 23397 13243
rect 23397 13209 23431 13243
rect 23431 13209 23440 13243
rect 23388 13200 23440 13209
rect 25320 13200 25372 13252
rect 26148 13200 26200 13252
rect 26608 13132 26660 13184
rect 37372 13175 37424 13184
rect 37372 13141 37381 13175
rect 37381 13141 37415 13175
rect 37415 13141 37424 13175
rect 37372 13132 37424 13141
rect 38200 13175 38252 13184
rect 38200 13141 38209 13175
rect 38209 13141 38243 13175
rect 38243 13141 38252 13175
rect 38200 13132 38252 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 2964 12928 3016 12980
rect 3056 12928 3108 12980
rect 4896 12928 4948 12980
rect 8300 12928 8352 12980
rect 10600 12928 10652 12980
rect 10692 12928 10744 12980
rect 13544 12928 13596 12980
rect 16948 12928 17000 12980
rect 1676 12860 1728 12912
rect 2044 12792 2096 12844
rect 2504 12792 2556 12844
rect 4804 12860 4856 12912
rect 6644 12860 6696 12912
rect 10140 12860 10192 12912
rect 13360 12860 13412 12912
rect 17776 12860 17828 12912
rect 19064 12860 19116 12912
rect 6552 12792 6604 12844
rect 2596 12724 2648 12776
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 4896 12656 4948 12708
rect 9956 12792 10008 12844
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 1768 12631 1820 12640
rect 1768 12597 1777 12631
rect 1777 12597 1811 12631
rect 1811 12597 1820 12631
rect 1768 12588 1820 12597
rect 8116 12588 8168 12640
rect 10508 12767 10560 12776
rect 10508 12733 10517 12767
rect 10517 12733 10551 12767
rect 10551 12733 10560 12767
rect 10508 12724 10560 12733
rect 11428 12724 11480 12776
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 17316 12792 17368 12844
rect 23112 12928 23164 12980
rect 23296 12860 23348 12912
rect 25780 12835 25832 12844
rect 12532 12724 12584 12733
rect 15568 12724 15620 12776
rect 17592 12724 17644 12776
rect 25780 12801 25789 12835
rect 25789 12801 25823 12835
rect 25823 12801 25832 12835
rect 25780 12792 25832 12801
rect 38016 12835 38068 12844
rect 38016 12801 38025 12835
rect 38025 12801 38059 12835
rect 38059 12801 38068 12835
rect 38016 12792 38068 12801
rect 23296 12767 23348 12776
rect 10600 12656 10652 12708
rect 17684 12656 17736 12708
rect 17868 12656 17920 12708
rect 23296 12733 23305 12767
rect 23305 12733 23339 12767
rect 23339 12733 23348 12767
rect 23296 12724 23348 12733
rect 23572 12767 23624 12776
rect 23572 12733 23581 12767
rect 23581 12733 23615 12767
rect 23615 12733 23624 12767
rect 23572 12724 23624 12733
rect 12256 12588 12308 12640
rect 12716 12588 12768 12640
rect 14648 12588 14700 12640
rect 24860 12656 24912 12708
rect 20076 12588 20128 12640
rect 22100 12631 22152 12640
rect 22100 12597 22109 12631
rect 22109 12597 22143 12631
rect 22143 12597 22152 12631
rect 38200 12631 38252 12640
rect 22100 12588 22152 12597
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2136 12384 2188 12436
rect 3792 12384 3844 12436
rect 6552 12384 6604 12436
rect 2596 12316 2648 12368
rect 4896 12316 4948 12368
rect 2780 12248 2832 12300
rect 3516 12248 3568 12300
rect 5724 12248 5776 12300
rect 1676 12180 1728 12232
rect 4620 12180 4672 12232
rect 5264 12180 5316 12232
rect 7564 12316 7616 12368
rect 6092 12248 6144 12300
rect 16672 12384 16724 12436
rect 17132 12384 17184 12436
rect 26056 12384 26108 12436
rect 38016 12384 38068 12436
rect 8300 12359 8352 12368
rect 8300 12325 8309 12359
rect 8309 12325 8343 12359
rect 8343 12325 8352 12359
rect 8300 12316 8352 12325
rect 10324 12316 10376 12368
rect 12164 12316 12216 12368
rect 8484 12248 8536 12300
rect 9496 12248 9548 12300
rect 17500 12316 17552 12368
rect 18144 12316 18196 12368
rect 24308 12316 24360 12368
rect 15936 12291 15988 12300
rect 15936 12257 15945 12291
rect 15945 12257 15979 12291
rect 15979 12257 15988 12291
rect 15936 12248 15988 12257
rect 17132 12248 17184 12300
rect 22744 12248 22796 12300
rect 23296 12248 23348 12300
rect 8852 12180 8904 12232
rect 14280 12223 14332 12232
rect 5080 12112 5132 12164
rect 7748 12112 7800 12164
rect 8208 12112 8260 12164
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 4896 12044 4948 12096
rect 5172 12044 5224 12096
rect 6000 12044 6052 12096
rect 7104 12044 7156 12096
rect 9404 12112 9456 12164
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 14924 12180 14976 12232
rect 17224 12180 17276 12232
rect 17868 12180 17920 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 22836 12180 22888 12232
rect 25228 12223 25280 12232
rect 25228 12189 25237 12223
rect 25237 12189 25271 12223
rect 25271 12189 25280 12223
rect 25228 12180 25280 12189
rect 28448 12223 28500 12232
rect 28448 12189 28457 12223
rect 28457 12189 28491 12223
rect 28491 12189 28500 12223
rect 28448 12180 28500 12189
rect 37372 12180 37424 12232
rect 10876 12155 10928 12164
rect 10876 12121 10885 12155
rect 10885 12121 10919 12155
rect 10919 12121 10928 12155
rect 10876 12112 10928 12121
rect 12532 12155 12584 12164
rect 12532 12121 12541 12155
rect 12541 12121 12575 12155
rect 12575 12121 12584 12155
rect 12532 12112 12584 12121
rect 13268 12155 13320 12164
rect 13268 12121 13277 12155
rect 13277 12121 13311 12155
rect 13311 12121 13320 12155
rect 13268 12112 13320 12121
rect 15016 12112 15068 12164
rect 19340 12112 19392 12164
rect 20260 12155 20312 12164
rect 20260 12121 20269 12155
rect 20269 12121 20303 12155
rect 20303 12121 20312 12155
rect 20260 12112 20312 12121
rect 22100 12112 22152 12164
rect 22376 12112 22428 12164
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 14648 12044 14700 12096
rect 15292 12044 15344 12096
rect 18420 12044 18472 12096
rect 19984 12044 20036 12096
rect 22744 12044 22796 12096
rect 25688 12087 25740 12096
rect 25688 12053 25697 12087
rect 25697 12053 25731 12087
rect 25731 12053 25740 12087
rect 25688 12044 25740 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 5632 11840 5684 11892
rect 7012 11840 7064 11892
rect 9128 11840 9180 11892
rect 9588 11840 9640 11892
rect 10232 11840 10284 11892
rect 23756 11883 23808 11892
rect 2596 11704 2648 11756
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 6184 11772 6236 11824
rect 4068 11568 4120 11620
rect 6460 11704 6512 11756
rect 8484 11772 8536 11824
rect 7840 11704 7892 11756
rect 5172 11636 5224 11688
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 6368 11636 6420 11688
rect 11336 11772 11388 11824
rect 13452 11815 13504 11824
rect 13452 11781 13461 11815
rect 13461 11781 13495 11815
rect 13495 11781 13504 11815
rect 13452 11772 13504 11781
rect 9772 11704 9824 11756
rect 10416 11704 10468 11756
rect 18144 11772 18196 11824
rect 18420 11815 18472 11824
rect 18420 11781 18429 11815
rect 18429 11781 18463 11815
rect 18463 11781 18472 11815
rect 18420 11772 18472 11781
rect 19984 11815 20036 11824
rect 19984 11781 19993 11815
rect 19993 11781 20027 11815
rect 20027 11781 20036 11815
rect 19984 11772 20036 11781
rect 23756 11849 23765 11883
rect 23765 11849 23799 11883
rect 23799 11849 23808 11883
rect 23756 11840 23808 11849
rect 24768 11840 24820 11892
rect 25228 11840 25280 11892
rect 25688 11840 25740 11892
rect 26240 11772 26292 11824
rect 14648 11747 14700 11756
rect 14648 11713 14657 11747
rect 14657 11713 14691 11747
rect 14691 11713 14700 11747
rect 14648 11704 14700 11713
rect 11152 11636 11204 11688
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 12256 11636 12308 11688
rect 14280 11636 14332 11688
rect 21732 11704 21784 11756
rect 23572 11704 23624 11756
rect 15384 11636 15436 11688
rect 18328 11679 18380 11688
rect 18328 11645 18337 11679
rect 18337 11645 18371 11679
rect 18371 11645 18380 11679
rect 18328 11636 18380 11645
rect 18972 11679 19024 11688
rect 18972 11645 18981 11679
rect 18981 11645 19015 11679
rect 19015 11645 19024 11679
rect 18972 11636 19024 11645
rect 20168 11636 20220 11688
rect 21272 11636 21324 11688
rect 23020 11636 23072 11688
rect 7288 11611 7340 11620
rect 7288 11577 7297 11611
rect 7297 11577 7331 11611
rect 7331 11577 7340 11611
rect 7288 11568 7340 11577
rect 9404 11568 9456 11620
rect 11888 11568 11940 11620
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 2136 11500 2188 11509
rect 2228 11500 2280 11552
rect 5448 11500 5500 11552
rect 7196 11500 7248 11552
rect 8300 11500 8352 11552
rect 8484 11500 8536 11552
rect 10968 11500 11020 11552
rect 11152 11500 11204 11552
rect 15200 11500 15252 11552
rect 20628 11568 20680 11620
rect 22836 11500 22888 11552
rect 24676 11636 24728 11688
rect 25136 11704 25188 11756
rect 25872 11704 25924 11756
rect 27712 11704 27764 11756
rect 23204 11568 23256 11620
rect 25872 11568 25924 11620
rect 26056 11636 26108 11688
rect 26332 11636 26384 11688
rect 26976 11636 27028 11688
rect 27344 11679 27396 11688
rect 27344 11645 27353 11679
rect 27353 11645 27387 11679
rect 27387 11645 27396 11679
rect 27344 11636 27396 11645
rect 31852 11568 31904 11620
rect 24952 11500 25004 11552
rect 26516 11500 26568 11552
rect 34428 11500 34480 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1584 11296 1636 11348
rect 2044 11296 2096 11348
rect 4068 11296 4120 11348
rect 5632 11296 5684 11348
rect 6552 11296 6604 11348
rect 11060 11296 11112 11348
rect 11980 11296 12032 11348
rect 12532 11296 12584 11348
rect 4988 11228 5040 11280
rect 7840 11228 7892 11280
rect 2228 11092 2280 11144
rect 2688 11092 2740 11144
rect 4068 11092 4120 11144
rect 4712 11160 4764 11212
rect 4252 11092 4304 11144
rect 5356 11160 5408 11212
rect 5540 11160 5592 11212
rect 10048 11228 10100 11280
rect 14740 11228 14792 11280
rect 15660 11228 15712 11280
rect 9496 11160 9548 11212
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 23204 11228 23256 11280
rect 19984 11160 20036 11212
rect 20352 11203 20404 11212
rect 20352 11169 20361 11203
rect 20361 11169 20395 11203
rect 20395 11169 20404 11203
rect 20352 11160 20404 11169
rect 7380 11092 7432 11144
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9312 11135 9364 11144
rect 9312 11101 9321 11135
rect 9321 11101 9355 11135
rect 9355 11101 9364 11135
rect 9312 11092 9364 11101
rect 9588 11092 9640 11144
rect 15200 11092 15252 11144
rect 20996 11092 21048 11144
rect 21732 11092 21784 11144
rect 22468 11092 22520 11144
rect 23756 11092 23808 11144
rect 5356 11067 5408 11076
rect 5356 11033 5365 11067
rect 5365 11033 5399 11067
rect 5399 11033 5408 11067
rect 5356 11024 5408 11033
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 6460 11024 6512 11076
rect 8208 11024 8260 11076
rect 10416 11067 10468 11076
rect 10416 11033 10425 11067
rect 10425 11033 10459 11067
rect 10459 11033 10468 11067
rect 10416 11024 10468 11033
rect 11060 11067 11112 11076
rect 11060 11033 11069 11067
rect 11069 11033 11103 11067
rect 11103 11033 11112 11067
rect 11060 11024 11112 11033
rect 11152 11067 11204 11076
rect 11152 11033 11161 11067
rect 11161 11033 11195 11067
rect 11195 11033 11204 11067
rect 11152 11024 11204 11033
rect 11704 11024 11756 11076
rect 12164 11024 12216 11076
rect 12624 11067 12676 11076
rect 12624 11033 12633 11067
rect 12633 11033 12667 11067
rect 12667 11033 12676 11067
rect 12624 11024 12676 11033
rect 12716 11067 12768 11076
rect 12716 11033 12725 11067
rect 12725 11033 12759 11067
rect 12759 11033 12768 11067
rect 15568 11067 15620 11076
rect 12716 11024 12768 11033
rect 15568 11033 15577 11067
rect 15577 11033 15611 11067
rect 15611 11033 15620 11067
rect 15568 11024 15620 11033
rect 15660 11067 15712 11076
rect 15660 11033 15669 11067
rect 15669 11033 15703 11067
rect 15703 11033 15712 11067
rect 16212 11067 16264 11076
rect 15660 11024 15712 11033
rect 16212 11033 16221 11067
rect 16221 11033 16255 11067
rect 16255 11033 16264 11067
rect 16212 11024 16264 11033
rect 20076 11024 20128 11076
rect 23848 11067 23900 11076
rect 23848 11033 23857 11067
rect 23857 11033 23891 11067
rect 23891 11033 23900 11067
rect 23848 11024 23900 11033
rect 24952 11296 25004 11348
rect 26056 11296 26108 11348
rect 27344 11296 27396 11348
rect 24216 11228 24268 11280
rect 37464 11228 37516 11280
rect 24676 11203 24728 11212
rect 24676 11169 24685 11203
rect 24685 11169 24719 11203
rect 24719 11169 24728 11203
rect 24676 11160 24728 11169
rect 26976 11203 27028 11212
rect 26976 11169 26985 11203
rect 26985 11169 27019 11203
rect 27019 11169 27028 11203
rect 26976 11160 27028 11169
rect 26516 11135 26568 11144
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 27988 11135 28040 11144
rect 27988 11101 27997 11135
rect 27997 11101 28031 11135
rect 28031 11101 28040 11135
rect 27988 11092 28040 11101
rect 31852 11135 31904 11144
rect 31852 11101 31861 11135
rect 31861 11101 31895 11135
rect 31895 11101 31904 11135
rect 31852 11092 31904 11101
rect 37188 11092 37240 11144
rect 2320 10956 2372 11008
rect 3240 10956 3292 11008
rect 7196 10956 7248 11008
rect 9680 10956 9732 11008
rect 10784 10956 10836 11008
rect 14372 10956 14424 11008
rect 14832 10999 14884 11008
rect 14832 10965 14841 10999
rect 14841 10965 14875 10999
rect 14875 10965 14884 10999
rect 14832 10956 14884 10965
rect 14924 10956 14976 11008
rect 17224 10956 17276 11008
rect 17316 10956 17368 11008
rect 19432 10956 19484 11008
rect 21180 10999 21232 11008
rect 21180 10965 21189 10999
rect 21189 10965 21223 10999
rect 21223 10965 21232 10999
rect 21180 10956 21232 10965
rect 25044 11024 25096 11076
rect 25320 11067 25372 11076
rect 25320 11033 25329 11067
rect 25329 11033 25363 11067
rect 25363 11033 25372 11067
rect 25320 11024 25372 11033
rect 28080 11024 28132 11076
rect 32588 11024 32640 11076
rect 33140 10956 33192 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 3424 10752 3476 10804
rect 5356 10795 5408 10804
rect 5356 10761 5365 10795
rect 5365 10761 5399 10795
rect 5399 10761 5408 10795
rect 5356 10752 5408 10761
rect 9312 10752 9364 10804
rect 2596 10727 2648 10736
rect 2596 10693 2605 10727
rect 2605 10693 2639 10727
rect 2639 10693 2648 10727
rect 2596 10684 2648 10693
rect 3516 10727 3568 10736
rect 3516 10693 3525 10727
rect 3525 10693 3559 10727
rect 3559 10693 3568 10727
rect 3516 10684 3568 10693
rect 7012 10684 7064 10736
rect 7104 10684 7156 10736
rect 9680 10727 9732 10736
rect 9680 10693 9689 10727
rect 9689 10693 9723 10727
rect 9723 10693 9732 10727
rect 10876 10752 10928 10804
rect 9680 10684 9732 10693
rect 11888 10727 11940 10736
rect 11888 10693 11897 10727
rect 11897 10693 11931 10727
rect 11931 10693 11940 10727
rect 11888 10684 11940 10693
rect 4804 10616 4856 10668
rect 6000 10616 6052 10668
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 11244 10616 11296 10668
rect 2412 10480 2464 10532
rect 7288 10548 7340 10600
rect 8484 10548 8536 10600
rect 11796 10591 11848 10600
rect 8300 10480 8352 10532
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 13452 10752 13504 10804
rect 14096 10684 14148 10736
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 17224 10752 17276 10804
rect 17960 10727 18012 10736
rect 17960 10693 17969 10727
rect 17969 10693 18003 10727
rect 18003 10693 18012 10727
rect 17960 10684 18012 10693
rect 18328 10752 18380 10804
rect 20260 10752 20312 10804
rect 23480 10752 23532 10804
rect 25320 10684 25372 10736
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 14832 10616 14884 10668
rect 17316 10616 17368 10668
rect 14556 10548 14608 10600
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 17868 10548 17920 10557
rect 16212 10480 16264 10532
rect 1768 10412 1820 10464
rect 3516 10412 3568 10464
rect 5172 10412 5224 10464
rect 7012 10412 7064 10464
rect 11336 10412 11388 10464
rect 14740 10412 14792 10464
rect 15200 10412 15252 10464
rect 15384 10412 15436 10464
rect 17408 10412 17460 10464
rect 18236 10548 18288 10600
rect 20904 10616 20956 10668
rect 21180 10616 21232 10668
rect 22468 10616 22520 10668
rect 24676 10616 24728 10668
rect 24860 10616 24912 10668
rect 20168 10548 20220 10600
rect 20628 10548 20680 10600
rect 22284 10548 22336 10600
rect 23848 10548 23900 10600
rect 21180 10455 21232 10464
rect 21180 10421 21189 10455
rect 21189 10421 21223 10455
rect 21223 10421 21232 10455
rect 21180 10412 21232 10421
rect 23112 10455 23164 10464
rect 23112 10421 23121 10455
rect 23121 10421 23155 10455
rect 23155 10421 23164 10455
rect 23112 10412 23164 10421
rect 24860 10455 24912 10464
rect 24860 10421 24869 10455
rect 24869 10421 24903 10455
rect 24903 10421 24912 10455
rect 24860 10412 24912 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 8852 10208 8904 10260
rect 12624 10208 12676 10260
rect 17868 10208 17920 10260
rect 8484 10140 8536 10192
rect 17960 10140 18012 10192
rect 2320 10115 2372 10124
rect 2320 10081 2329 10115
rect 2329 10081 2363 10115
rect 2363 10081 2372 10115
rect 2320 10072 2372 10081
rect 2964 10072 3016 10124
rect 3424 10072 3476 10124
rect 4896 10072 4948 10124
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 5080 10004 5132 10056
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 9128 10072 9180 10124
rect 19340 10140 19392 10192
rect 19984 10208 20036 10260
rect 22284 10251 22336 10260
rect 22284 10217 22293 10251
rect 22293 10217 22327 10251
rect 22327 10217 22336 10251
rect 22284 10208 22336 10217
rect 25044 10208 25096 10260
rect 23020 10140 23072 10192
rect 9864 10004 9916 10056
rect 11152 10004 11204 10056
rect 2136 9936 2188 9988
rect 11428 9936 11480 9988
rect 11796 9936 11848 9988
rect 20444 10072 20496 10124
rect 12992 10004 13044 10056
rect 22008 10004 22060 10056
rect 23112 10004 23164 10056
rect 24584 10004 24636 10056
rect 14832 9936 14884 9988
rect 17408 9979 17460 9988
rect 17408 9945 17417 9979
rect 17417 9945 17451 9979
rect 17451 9945 17460 9979
rect 36452 10004 36504 10056
rect 17408 9936 17460 9945
rect 1492 9868 1544 9920
rect 4988 9911 5040 9920
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 9220 9868 9272 9920
rect 16488 9868 16540 9920
rect 38200 9911 38252 9920
rect 38200 9877 38209 9911
rect 38209 9877 38243 9911
rect 38243 9877 38252 9911
rect 38200 9868 38252 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2596 9664 2648 9716
rect 14740 9664 14792 9716
rect 20628 9664 20680 9716
rect 21180 9664 21232 9716
rect 8208 9639 8260 9648
rect 2596 9528 2648 9580
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 5264 9528 5316 9580
rect 6460 9528 6512 9580
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 8208 9605 8217 9639
rect 8217 9605 8251 9639
rect 8251 9605 8260 9639
rect 8208 9596 8260 9605
rect 9220 9639 9272 9648
rect 9220 9605 9229 9639
rect 9229 9605 9263 9639
rect 9263 9605 9272 9639
rect 9220 9596 9272 9605
rect 10416 9596 10468 9648
rect 30380 9596 30432 9648
rect 6552 9528 6604 9537
rect 10232 9571 10284 9580
rect 7104 9460 7156 9512
rect 5816 9392 5868 9444
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 24124 9528 24176 9580
rect 34244 9528 34296 9580
rect 11060 9460 11112 9512
rect 12072 9460 12124 9512
rect 20444 9460 20496 9512
rect 20812 9460 20864 9512
rect 34336 9503 34388 9512
rect 34336 9469 34345 9503
rect 34345 9469 34379 9503
rect 34379 9469 34388 9503
rect 34336 9460 34388 9469
rect 8484 9392 8536 9444
rect 36452 9392 36504 9444
rect 3792 9367 3844 9376
rect 3792 9333 3801 9367
rect 3801 9333 3835 9367
rect 3835 9333 3844 9367
rect 3792 9324 3844 9333
rect 6644 9367 6696 9376
rect 6644 9333 6653 9367
rect 6653 9333 6687 9367
rect 6687 9333 6696 9367
rect 6644 9324 6696 9333
rect 11796 9324 11848 9376
rect 19340 9324 19392 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 6828 9120 6880 9172
rect 10140 9120 10192 9172
rect 11612 9120 11664 9172
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 26332 9163 26384 9172
rect 26332 9129 26341 9163
rect 26341 9129 26375 9163
rect 26375 9129 26384 9163
rect 26332 9120 26384 9129
rect 2504 9052 2556 9104
rect 3424 9052 3476 9104
rect 2872 8984 2924 9036
rect 20444 9027 20496 9036
rect 20444 8993 20453 9027
rect 20453 8993 20487 9027
rect 20487 8993 20496 9027
rect 20444 8984 20496 8993
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 4988 8916 5040 8968
rect 6644 8916 6696 8968
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 13176 8916 13228 8968
rect 23848 8916 23900 8968
rect 26332 8959 26384 8968
rect 26332 8925 26341 8959
rect 26341 8925 26375 8959
rect 26375 8925 26384 8959
rect 26332 8916 26384 8925
rect 32588 8959 32640 8968
rect 32588 8925 32597 8959
rect 32597 8925 32631 8959
rect 32631 8925 32640 8959
rect 32588 8916 32640 8925
rect 2872 8823 2924 8832
rect 2872 8789 2881 8823
rect 2881 8789 2915 8823
rect 2915 8789 2924 8823
rect 2872 8780 2924 8789
rect 3056 8780 3108 8832
rect 4620 8823 4672 8832
rect 4620 8789 4629 8823
rect 4629 8789 4663 8823
rect 4663 8789 4672 8823
rect 4620 8780 4672 8789
rect 24768 8780 24820 8832
rect 34152 8780 34204 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1952 8576 2004 8628
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 5172 8576 5224 8628
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 4620 8440 4672 8492
rect 15200 8440 15252 8492
rect 20996 8483 21048 8492
rect 20996 8449 21005 8483
rect 21005 8449 21039 8483
rect 21039 8449 21048 8483
rect 20996 8440 21048 8449
rect 27068 8440 27120 8492
rect 38108 8483 38160 8492
rect 38108 8449 38117 8483
rect 38117 8449 38151 8483
rect 38151 8449 38160 8483
rect 38108 8440 38160 8449
rect 3792 8372 3844 8424
rect 13268 8372 13320 8424
rect 12440 8304 12492 8356
rect 28908 8304 28960 8356
rect 20996 8236 21048 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3332 8032 3384 8084
rect 14832 8075 14884 8084
rect 14832 8041 14841 8075
rect 14841 8041 14875 8075
rect 14875 8041 14884 8075
rect 14832 8032 14884 8041
rect 20812 8075 20864 8084
rect 20812 8041 20821 8075
rect 20821 8041 20855 8075
rect 20855 8041 20864 8075
rect 20812 8032 20864 8041
rect 9128 7896 9180 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 3516 7828 3568 7880
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 12440 7828 12492 7880
rect 14740 7871 14792 7880
rect 14740 7837 14749 7871
rect 14749 7837 14783 7871
rect 14783 7837 14792 7871
rect 14740 7828 14792 7837
rect 19340 7828 19392 7880
rect 20996 7871 21048 7880
rect 20996 7837 21005 7871
rect 21005 7837 21039 7871
rect 21039 7837 21048 7871
rect 20996 7828 21048 7837
rect 24768 7871 24820 7880
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 24768 7828 24820 7837
rect 28908 7828 28960 7880
rect 33140 7828 33192 7880
rect 34152 7828 34204 7880
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 6828 7692 6880 7744
rect 17500 7692 17552 7744
rect 25964 7692 26016 7744
rect 31668 7692 31720 7744
rect 34796 7692 34848 7744
rect 38200 7735 38252 7744
rect 38200 7701 38209 7735
rect 38209 7701 38243 7735
rect 38243 7701 38252 7735
rect 38200 7692 38252 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1860 7420 1912 7472
rect 2872 7420 2924 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 3240 7352 3292 7404
rect 9128 7352 9180 7404
rect 21088 7352 21140 7404
rect 34428 7352 34480 7404
rect 2964 7259 3016 7268
rect 2964 7225 2973 7259
rect 2973 7225 3007 7259
rect 3007 7225 3016 7259
rect 2964 7216 3016 7225
rect 12900 7216 12952 7268
rect 19984 7216 20036 7268
rect 4620 7148 4672 7200
rect 17040 7148 17092 7200
rect 37740 7148 37792 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 34796 6740 34848 6792
rect 2780 6672 2832 6724
rect 2136 6604 2188 6656
rect 38016 6604 38068 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 15200 6239 15252 6248
rect 15200 6205 15209 6239
rect 15209 6205 15243 6239
rect 15243 6205 15252 6239
rect 15200 6196 15252 6205
rect 24492 6196 24544 6248
rect 37464 6239 37516 6248
rect 37464 6205 37473 6239
rect 37473 6205 37507 6239
rect 37507 6205 37516 6239
rect 37464 6196 37516 6205
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 2872 5856 2924 5865
rect 14556 5788 14608 5840
rect 15200 5763 15252 5772
rect 15200 5729 15209 5763
rect 15209 5729 15243 5763
rect 15243 5729 15252 5763
rect 15200 5720 15252 5729
rect 1492 5652 1544 5704
rect 3608 5652 3660 5704
rect 5448 5652 5500 5704
rect 15292 5627 15344 5636
rect 15292 5593 15301 5627
rect 15301 5593 15335 5627
rect 15335 5593 15344 5627
rect 15292 5584 15344 5593
rect 1768 5559 1820 5568
rect 1768 5525 1777 5559
rect 1777 5525 1811 5559
rect 1811 5525 1820 5559
rect 1768 5516 1820 5525
rect 4712 5516 4764 5568
rect 24768 5516 24820 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4712 5219 4764 5228
rect 4712 5185 4721 5219
rect 4721 5185 4755 5219
rect 4755 5185 4764 5219
rect 4712 5176 4764 5185
rect 11704 5176 11756 5228
rect 24768 5219 24820 5228
rect 24768 5185 24777 5219
rect 24777 5185 24811 5219
rect 24811 5185 24820 5219
rect 24768 5176 24820 5185
rect 38016 5219 38068 5228
rect 38016 5185 38025 5219
rect 38025 5185 38059 5219
rect 38059 5185 38068 5219
rect 38016 5176 38068 5185
rect 4620 4972 4672 5024
rect 11704 4972 11756 5024
rect 30472 4972 30524 5024
rect 38200 5015 38252 5024
rect 38200 4981 38209 5015
rect 38209 4981 38243 5015
rect 38243 4981 38252 5015
rect 38200 4972 38252 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 32128 4564 32180 4616
rect 37740 4564 37792 4616
rect 1676 4539 1728 4548
rect 1676 4505 1685 4539
rect 1685 4505 1719 4539
rect 1719 4505 1728 4539
rect 1676 4496 1728 4505
rect 12164 4428 12216 4480
rect 35348 4471 35400 4480
rect 35348 4437 35357 4471
rect 35357 4437 35391 4471
rect 35391 4437 35400 4471
rect 35348 4428 35400 4437
rect 38200 4471 38252 4480
rect 38200 4437 38209 4471
rect 38209 4437 38243 4471
rect 38243 4437 38252 4471
rect 38200 4428 38252 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 37924 4088 37976 4140
rect 39304 3884 39356 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2228 3680 2280 3732
rect 37832 3544 37884 3596
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 37924 3476 37976 3528
rect 27988 3340 28040 3392
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3976 3136 4028 3188
rect 34244 3136 34296 3188
rect 4620 3068 4672 3120
rect 13176 3068 13228 3120
rect 1952 3000 2004 3052
rect 3240 3000 3292 3052
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 25780 3043 25832 3052
rect 25780 3009 25789 3043
rect 25789 3009 25823 3043
rect 25823 3009 25832 3043
rect 37280 3068 37332 3120
rect 25780 3000 25832 3009
rect 36728 3000 36780 3052
rect 11612 2932 11664 2984
rect 28448 2932 28500 2984
rect 37464 2975 37516 2984
rect 37464 2941 37473 2975
rect 37473 2941 37507 2975
rect 37507 2941 37516 2975
rect 37464 2932 37516 2941
rect 11152 2864 11204 2916
rect 664 2796 716 2848
rect 16856 2839 16908 2848
rect 16856 2805 16865 2839
rect 16865 2805 16899 2839
rect 16899 2805 16908 2839
rect 16856 2796 16908 2805
rect 20628 2796 20680 2848
rect 25228 2796 25280 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 7104 2592 7156 2644
rect 10232 2592 10284 2644
rect 14740 2592 14792 2644
rect 18236 2635 18288 2644
rect 18236 2601 18245 2635
rect 18245 2601 18279 2635
rect 18279 2601 18288 2635
rect 18236 2592 18288 2601
rect 22008 2635 22060 2644
rect 22008 2601 22017 2635
rect 22017 2601 22051 2635
rect 22051 2601 22060 2635
rect 22008 2592 22060 2601
rect 24676 2592 24728 2644
rect 26332 2592 26384 2644
rect 27436 2592 27488 2644
rect 20 2524 72 2576
rect 4712 2456 4764 2508
rect 22284 2524 22336 2576
rect 31576 2524 31628 2576
rect 8484 2456 8536 2508
rect 13176 2499 13228 2508
rect 1676 2363 1728 2372
rect 1676 2329 1685 2363
rect 1685 2329 1719 2363
rect 1719 2329 1728 2363
rect 1676 2320 1728 2329
rect 3424 2320 3476 2372
rect 6460 2388 6512 2440
rect 7104 2388 7156 2440
rect 8392 2388 8444 2440
rect 9680 2388 9732 2440
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 13176 2465 13185 2499
rect 13185 2465 13219 2499
rect 13219 2465 13228 2499
rect 13176 2456 13228 2465
rect 20628 2456 20680 2508
rect 14188 2388 14240 2440
rect 6828 2320 6880 2372
rect 1768 2295 1820 2304
rect 1768 2261 1777 2295
rect 1777 2261 1811 2295
rect 1811 2261 1820 2295
rect 1768 2252 1820 2261
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 3884 2252 3936 2304
rect 5172 2252 5224 2304
rect 9036 2252 9088 2304
rect 11336 2320 11388 2372
rect 16856 2388 16908 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18052 2388 18104 2440
rect 19340 2388 19392 2440
rect 19984 2388 20036 2440
rect 21916 2388 21968 2440
rect 24860 2456 24912 2508
rect 23848 2388 23900 2440
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 25964 2431 26016 2440
rect 25964 2397 25973 2431
rect 25973 2397 26007 2431
rect 26007 2397 26016 2431
rect 25964 2388 26016 2397
rect 27068 2388 27120 2440
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 30472 2431 30524 2440
rect 30472 2397 30481 2431
rect 30481 2397 30515 2431
rect 30515 2397 30524 2431
rect 30472 2388 30524 2397
rect 31668 2388 31720 2440
rect 33324 2388 33376 2440
rect 37280 2456 37332 2508
rect 35348 2388 35400 2440
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 27804 2320 27856 2372
rect 28356 2320 28408 2372
rect 10968 2252 11020 2304
rect 14832 2252 14884 2304
rect 16120 2252 16172 2304
rect 17408 2252 17460 2304
rect 20628 2252 20680 2304
rect 22560 2252 22612 2304
rect 25136 2252 25188 2304
rect 25780 2252 25832 2304
rect 29644 2252 29696 2304
rect 30288 2252 30340 2304
rect 31576 2252 31628 2304
rect 32864 2252 32916 2304
rect 33508 2252 33560 2304
rect 34796 2252 34848 2304
rect 36084 2252 36136 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 9036 2048 9088 2100
rect 12992 2048 13044 2100
rect 1768 1980 1820 2032
rect 15016 1980 15068 2032
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 2594 39200 2650 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14186 39200 14242 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 17406 39200 17462 39800
rect 18694 39200 18750 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 21914 39200 21970 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25134 39200 25190 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 28354 39200 28410 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 34256 39222 34468 39250
rect 32 36174 60 39200
rect 1320 36786 1348 39200
rect 1766 38856 1822 38865
rect 1766 38791 1822 38800
rect 1780 37466 1808 38791
rect 1768 37460 1820 37466
rect 1768 37402 1820 37408
rect 2320 37256 2372 37262
rect 2320 37198 2372 37204
rect 2608 37210 2636 39200
rect 2870 38176 2926 38185
rect 2870 38111 2926 38120
rect 2780 37256 2832 37262
rect 2608 37204 2780 37210
rect 2608 37198 2832 37204
rect 1308 36780 1360 36786
rect 1308 36722 1360 36728
rect 1860 36576 1912 36582
rect 1860 36518 1912 36524
rect 20 36168 72 36174
rect 20 36110 72 36116
rect 1676 35692 1728 35698
rect 1676 35634 1728 35640
rect 1492 35488 1544 35494
rect 1688 35465 1716 35634
rect 1492 35430 1544 35436
rect 1674 35456 1730 35465
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1412 23225 1440 24754
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1400 20460 1452 20466
rect 1400 20402 1452 20408
rect 1412 19145 1440 20402
rect 1398 19136 1454 19145
rect 1398 19071 1454 19080
rect 1504 16998 1532 35430
rect 1674 35391 1730 35400
rect 1766 34776 1822 34785
rect 1766 34711 1822 34720
rect 1780 34610 1808 34711
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1766 33416 1822 33425
rect 1766 33351 1768 33360
rect 1820 33351 1822 33360
rect 1768 33322 1820 33328
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1780 32065 1808 32166
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 1872 31822 1900 36518
rect 2044 32428 2096 32434
rect 2044 32370 2096 32376
rect 1860 31816 1912 31822
rect 1860 31758 1912 31764
rect 1766 31376 1822 31385
rect 1766 31311 1768 31320
rect 1820 31311 1822 31320
rect 1768 31282 1820 31288
rect 2056 30258 2084 32370
rect 1860 30252 1912 30258
rect 1860 30194 1912 30200
rect 2044 30252 2096 30258
rect 2044 30194 2096 30200
rect 1766 30016 1822 30025
rect 1766 29951 1822 29960
rect 1780 29646 1808 29951
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1584 28960 1636 28966
rect 1584 28902 1636 28908
rect 1596 27674 1624 28902
rect 1780 28665 1808 29106
rect 1872 29102 1900 30194
rect 2332 29782 2360 37198
rect 2608 37182 2820 37198
rect 2688 36576 2740 36582
rect 2688 36518 2740 36524
rect 2596 35488 2648 35494
rect 2596 35430 2648 35436
rect 2608 35018 2636 35430
rect 2700 35034 2728 36518
rect 2884 36174 2912 38111
rect 2964 37256 3016 37262
rect 2964 37198 3016 37204
rect 2872 36168 2924 36174
rect 2872 36110 2924 36116
rect 2596 35012 2648 35018
rect 2700 35006 2820 35034
rect 2596 34954 2648 34960
rect 2688 34944 2740 34950
rect 2688 34886 2740 34892
rect 2700 34542 2728 34886
rect 2688 34536 2740 34542
rect 2688 34478 2740 34484
rect 2700 33590 2728 34478
rect 2792 33590 2820 35006
rect 2872 34604 2924 34610
rect 2872 34546 2924 34552
rect 2688 33584 2740 33590
rect 2688 33526 2740 33532
rect 2780 33584 2832 33590
rect 2780 33526 2832 33532
rect 2700 32994 2728 33526
rect 2608 32978 2728 32994
rect 2596 32972 2728 32978
rect 2648 32966 2728 32972
rect 2596 32914 2648 32920
rect 2700 31890 2728 32966
rect 2884 32842 2912 34546
rect 2872 32836 2924 32842
rect 2872 32778 2924 32784
rect 2976 32026 3004 37198
rect 3252 37126 3280 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37262 4660 37726
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 5828 37210 5856 39200
rect 6092 37392 6144 37398
rect 6092 37334 6144 37340
rect 5828 37182 6040 37210
rect 6012 37126 6040 37182
rect 3240 37120 3292 37126
rect 3240 37062 3292 37068
rect 5724 37120 5776 37126
rect 5724 37062 5776 37068
rect 6000 37120 6052 37126
rect 6000 37062 6052 37068
rect 3514 36816 3570 36825
rect 5736 36786 5764 37062
rect 6104 36854 6132 37334
rect 6472 37262 6500 39200
rect 7760 37262 7788 39200
rect 6460 37256 6512 37262
rect 6460 37198 6512 37204
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 6564 36922 6592 37198
rect 8024 37120 8076 37126
rect 8024 37062 8076 37068
rect 6552 36916 6604 36922
rect 6552 36858 6604 36864
rect 6092 36848 6144 36854
rect 6092 36790 6144 36796
rect 3514 36751 3570 36760
rect 4712 36780 4764 36786
rect 3424 36644 3476 36650
rect 3424 36586 3476 36592
rect 3436 35698 3464 36586
rect 3424 35692 3476 35698
rect 3424 35634 3476 35640
rect 3148 35284 3200 35290
rect 3148 35226 3200 35232
rect 3160 33454 3188 35226
rect 3332 35080 3384 35086
rect 3332 35022 3384 35028
rect 3344 34746 3372 35022
rect 3332 34740 3384 34746
rect 3332 34682 3384 34688
rect 3436 33998 3464 35634
rect 3424 33992 3476 33998
rect 3424 33934 3476 33940
rect 3148 33448 3200 33454
rect 3148 33390 3200 33396
rect 2964 32020 3016 32026
rect 2964 31962 3016 31968
rect 2688 31884 2740 31890
rect 2688 31826 2740 31832
rect 2412 31816 2464 31822
rect 2412 31758 2464 31764
rect 3148 31816 3200 31822
rect 3148 31758 3200 31764
rect 2320 29776 2372 29782
rect 2320 29718 2372 29724
rect 1952 29504 2004 29510
rect 1952 29446 2004 29452
rect 1860 29096 1912 29102
rect 1860 29038 1912 29044
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 1872 28558 1900 29038
rect 1860 28552 1912 28558
rect 1860 28494 1912 28500
rect 1768 28076 1820 28082
rect 1768 28018 1820 28024
rect 1584 27668 1636 27674
rect 1584 27610 1636 27616
rect 1780 27305 1808 28018
rect 1766 27296 1822 27305
rect 1766 27231 1822 27240
rect 1676 26988 1728 26994
rect 1676 26930 1728 26936
rect 1688 26625 1716 26930
rect 1860 26852 1912 26858
rect 1860 26794 1912 26800
rect 1674 26616 1730 26625
rect 1674 26551 1730 26560
rect 1872 26489 1900 26794
rect 1858 26480 1914 26489
rect 1858 26415 1914 26424
rect 1584 25288 1636 25294
rect 1584 25230 1636 25236
rect 1766 25256 1822 25265
rect 1596 24993 1624 25230
rect 1766 25191 1822 25200
rect 1780 25158 1808 25191
rect 1768 25152 1820 25158
rect 1768 25094 1820 25100
rect 1582 24984 1638 24993
rect 1582 24919 1638 24928
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1780 23905 1808 24006
rect 1766 23896 1822 23905
rect 1766 23831 1822 23840
rect 1964 23118 1992 29446
rect 2228 27872 2280 27878
rect 2228 27814 2280 27820
rect 2240 27713 2268 27814
rect 2226 27704 2282 27713
rect 2226 27639 2282 27648
rect 2424 26450 2452 31758
rect 3160 31482 3188 31758
rect 3148 31476 3200 31482
rect 3148 31418 3200 31424
rect 3436 31346 3464 33934
rect 3424 31340 3476 31346
rect 3424 31282 3476 31288
rect 3148 29028 3200 29034
rect 3148 28970 3200 28976
rect 2872 28416 2924 28422
rect 2872 28358 2924 28364
rect 2412 26444 2464 26450
rect 2412 26386 2464 26392
rect 2884 26314 2912 28358
rect 3160 27402 3188 28970
rect 3332 28484 3384 28490
rect 3332 28426 3384 28432
rect 3148 27396 3200 27402
rect 3148 27338 3200 27344
rect 2872 26308 2924 26314
rect 2872 26250 2924 26256
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 1952 23112 2004 23118
rect 1952 23054 2004 23060
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1596 17338 1624 21966
rect 1768 21888 1820 21894
rect 1766 21856 1768 21865
rect 1820 21856 1822 21865
rect 1766 21791 1822 21800
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1780 20505 1808 21490
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1688 18766 1716 19110
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1688 18426 1716 18702
rect 1766 18456 1822 18465
rect 1676 18420 1728 18426
rect 1766 18391 1822 18400
rect 1676 18362 1728 18368
rect 1780 17678 1808 18391
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1688 17105 1716 17138
rect 1674 17096 1730 17105
rect 1674 17031 1730 17040
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1688 14414 1716 16526
rect 1780 16522 1808 17478
rect 1768 16516 1820 16522
rect 1768 16458 1820 16464
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1780 15065 1808 15302
rect 1766 15056 1822 15065
rect 1766 14991 1822 15000
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1596 11354 1624 13874
rect 1688 12918 1716 14350
rect 1768 13728 1820 13734
rect 1766 13696 1768 13705
rect 1820 13696 1822 13705
rect 1766 13631 1822 13640
rect 1676 12912 1728 12918
rect 1676 12854 1728 12860
rect 1688 12238 1716 12854
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 12345 1808 12582
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10062 1808 10406
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 5710 1532 9862
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7585 1624 7822
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1872 7478 1900 22918
rect 2424 22778 2452 23598
rect 2412 22772 2464 22778
rect 2412 22714 2464 22720
rect 2044 22704 2096 22710
rect 2044 22646 2096 22652
rect 1952 20528 2004 20534
rect 1952 20470 2004 20476
rect 1964 16454 1992 20470
rect 2056 17542 2084 22646
rect 2228 21344 2280 21350
rect 2228 21286 2280 21292
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2136 20052 2188 20058
rect 2136 19994 2188 20000
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 1964 8634 1992 14826
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2056 11354 2084 12786
rect 2148 12442 2176 19994
rect 2240 17678 2268 21286
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 13394 2452 14350
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2516 12850 2544 21286
rect 2596 17060 2648 17066
rect 2596 17002 2648 17008
rect 2608 16697 2636 17002
rect 2594 16688 2650 16697
rect 2594 16623 2650 16632
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2608 15910 2636 16050
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2608 12782 2636 13806
rect 2596 12776 2648 12782
rect 2516 12724 2596 12730
rect 2516 12718 2648 12724
rect 2516 12702 2636 12718
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2148 9994 2176 11494
rect 2240 11150 2268 11494
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2332 10130 2360 10950
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 2226 9616 2282 9625
rect 2226 9551 2282 9560
rect 2240 8974 2268 9551
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2424 8786 2452 10474
rect 2516 9110 2544 12702
rect 2608 12653 2636 12702
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2608 11762 2636 12310
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2700 11150 2728 24550
rect 3344 24138 3372 28426
rect 3528 27402 3556 36751
rect 4712 36722 4764 36728
rect 5724 36780 5776 36786
rect 5724 36722 5776 36728
rect 7656 36780 7708 36786
rect 7656 36722 7708 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4724 36378 4752 36722
rect 6460 36576 6512 36582
rect 6460 36518 6512 36524
rect 4712 36372 4764 36378
rect 4712 36314 4764 36320
rect 6472 36242 6500 36518
rect 7668 36310 7696 36722
rect 7748 36576 7800 36582
rect 7746 36544 7748 36553
rect 7800 36544 7802 36553
rect 7746 36479 7802 36488
rect 7656 36304 7708 36310
rect 7656 36246 7708 36252
rect 6460 36236 6512 36242
rect 6460 36178 6512 36184
rect 6552 36100 6604 36106
rect 6552 36042 6604 36048
rect 6828 36100 6880 36106
rect 6828 36042 6880 36048
rect 3608 35692 3660 35698
rect 3608 35634 3660 35640
rect 3620 35290 3648 35634
rect 4068 35624 4120 35630
rect 4068 35566 4120 35572
rect 3976 35488 4028 35494
rect 3976 35430 4028 35436
rect 3608 35284 3660 35290
rect 3608 35226 3660 35232
rect 3988 34678 4016 35430
rect 4080 35290 4108 35566
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 35284 4120 35290
rect 4068 35226 4120 35232
rect 4896 35284 4948 35290
rect 4896 35226 4948 35232
rect 3976 34672 4028 34678
rect 4080 34649 4108 35226
rect 4620 34944 4672 34950
rect 4620 34886 4672 34892
rect 3976 34614 4028 34620
rect 4066 34640 4122 34649
rect 4066 34575 4122 34584
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 34202 4660 34886
rect 4620 34196 4672 34202
rect 4620 34138 4672 34144
rect 4804 33652 4856 33658
rect 4804 33594 4856 33600
rect 4620 33312 4672 33318
rect 4620 33254 4672 33260
rect 4712 33312 4764 33318
rect 4712 33254 4764 33260
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4160 31884 4212 31890
rect 4080 31844 4160 31872
rect 4080 31482 4108 31844
rect 4160 31826 4212 31832
rect 4068 31476 4120 31482
rect 4068 31418 4120 31424
rect 3884 31136 3936 31142
rect 3884 31078 3936 31084
rect 3792 29164 3844 29170
rect 3792 29106 3844 29112
rect 3516 27396 3568 27402
rect 3516 27338 3568 27344
rect 3422 26344 3478 26353
rect 3422 26279 3424 26288
rect 3476 26279 3478 26288
rect 3424 26250 3476 26256
rect 3804 25906 3832 29106
rect 3896 25974 3924 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 3976 28552 4028 28558
rect 3976 28494 4028 28500
rect 3988 28014 4016 28494
rect 3976 28008 4028 28014
rect 3976 27950 4028 27956
rect 3988 27538 4016 27950
rect 3976 27532 4028 27538
rect 3976 27474 4028 27480
rect 4080 27418 4108 29242
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3988 27390 4108 27418
rect 3988 27062 4016 27390
rect 3976 27056 4028 27062
rect 3976 26998 4028 27004
rect 3884 25968 3936 25974
rect 3884 25910 3936 25916
rect 3792 25900 3844 25906
rect 3792 25842 3844 25848
rect 3700 25696 3752 25702
rect 3700 25638 3752 25644
rect 3608 25288 3660 25294
rect 3608 25230 3660 25236
rect 3620 24750 3648 25230
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3620 24274 3648 24686
rect 3608 24268 3660 24274
rect 3608 24210 3660 24216
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 2780 23792 2832 23798
rect 2780 23734 2832 23740
rect 2792 23526 2820 23734
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 3620 22760 3648 24210
rect 3712 23798 3740 25638
rect 3700 23792 3752 23798
rect 3700 23734 3752 23740
rect 3700 22772 3752 22778
rect 3620 22732 3700 22760
rect 3700 22714 3752 22720
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3160 20262 3188 20946
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3160 19922 3188 20198
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3344 19786 3372 20742
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 3332 19780 3384 19786
rect 3332 19722 3384 19728
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 2884 14618 2912 19382
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2976 16658 3004 17138
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2976 16114 3004 16594
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2976 13530 3004 15438
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2792 12306 2820 13330
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2976 12986 3004 13126
rect 3068 12986 3096 18702
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 3160 14618 3188 15574
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2870 11656 2926 11665
rect 2870 11591 2926 11600
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2608 9722 2636 10678
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2594 9616 2650 9625
rect 2792 9586 2820 10231
rect 2594 9551 2596 9560
rect 2648 9551 2650 9560
rect 2780 9580 2832 9586
rect 2596 9522 2648 9528
rect 2780 9522 2832 9528
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2884 9042 2912 11591
rect 3252 11014 3280 19722
rect 3436 18834 3464 22374
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3620 19718 3648 22170
rect 3712 22098 3740 22714
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 3804 22001 3832 25842
rect 3988 25820 4016 26998
rect 4068 26784 4120 26790
rect 4068 26726 4120 26732
rect 4080 25838 4108 26726
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3896 25792 4016 25820
rect 4068 25832 4120 25838
rect 3790 21992 3846 22001
rect 3790 21927 3846 21936
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3332 18352 3384 18358
rect 3332 18294 3384 18300
rect 3344 16250 3372 18294
rect 3436 17202 3464 18770
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3528 16794 3556 17070
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3424 16516 3476 16522
rect 3424 16458 3476 16464
rect 3436 16250 3464 16458
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2332 8758 2452 8786
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1688 6905 1716 7346
rect 1674 6896 1730 6905
rect 1674 6831 1730 6840
rect 2148 6662 2176 8434
rect 2332 6866 2360 8758
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1768 5568 1820 5574
rect 1766 5536 1768 5545
rect 1820 5536 1822 5545
rect 1766 5471 1822 5480
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1688 4185 1716 4490
rect 1674 4176 1730 4185
rect 1674 4111 1730 4120
rect 2240 3738 2268 6734
rect 2792 6730 2820 8871
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8498 2912 8774
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2884 5914 2912 7414
rect 2976 7274 3004 10066
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8498 3096 8774
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3344 8090 3372 14894
rect 3422 14240 3478 14249
rect 3422 14175 3478 14184
rect 3436 13394 3464 14175
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3436 10810 3464 13330
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3528 11762 3556 12242
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3514 10976 3570 10985
rect 3514 10911 3570 10920
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3436 10130 3464 10746
rect 3528 10742 3556 10911
rect 3516 10736 3568 10742
rect 3516 10678 3568 10684
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7410 3280 7686
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 1768 3528 1820 3534
rect 1766 3496 1768 3505
rect 1820 3496 1822 3505
rect 1766 3431 1822 3440
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 676 800 704 2790
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 18 200 74 800
rect 662 200 718 800
rect 1688 785 1716 2314
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1780 2038 1808 2246
rect 1768 2032 1820 2038
rect 1768 1974 1820 1980
rect 1964 800 1992 2994
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 2145 2544 2246
rect 2502 2136 2558 2145
rect 2502 2071 2558 2080
rect 3252 800 3280 2994
rect 3436 2378 3464 9046
rect 3528 8634 3556 10406
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3528 7886 3556 8570
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3620 5710 3648 19654
rect 3712 19514 3740 20266
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 3712 16522 3740 18294
rect 3804 17270 3832 21927
rect 3792 17264 3844 17270
rect 3792 17206 3844 17212
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3804 15094 3832 16934
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14550 3740 14894
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3896 14414 3924 25792
rect 4068 25774 4120 25780
rect 4528 25832 4580 25838
rect 4632 25820 4660 33254
rect 4724 32910 4752 33254
rect 4816 33114 4844 33594
rect 4804 33108 4856 33114
rect 4804 33050 4856 33056
rect 4712 32904 4764 32910
rect 4712 32846 4764 32852
rect 4908 32774 4936 35226
rect 5356 35148 5408 35154
rect 5356 35090 5408 35096
rect 5368 34746 5396 35090
rect 6564 34746 6592 36042
rect 5356 34740 5408 34746
rect 5356 34682 5408 34688
rect 6552 34740 6604 34746
rect 6552 34682 6604 34688
rect 5724 34604 5776 34610
rect 5724 34546 5776 34552
rect 6276 34604 6328 34610
rect 6276 34546 6328 34552
rect 5540 33448 5592 33454
rect 5540 33390 5592 33396
rect 5552 32978 5580 33390
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 4896 32768 4948 32774
rect 4896 32710 4948 32716
rect 4908 31278 4936 32710
rect 5632 32224 5684 32230
rect 5632 32166 5684 32172
rect 5354 31376 5410 31385
rect 5354 31311 5356 31320
rect 5408 31311 5410 31320
rect 5356 31282 5408 31288
rect 4896 31272 4948 31278
rect 4896 31214 4948 31220
rect 4712 30048 4764 30054
rect 4712 29990 4764 29996
rect 4724 27062 4752 29990
rect 5644 29238 5672 32166
rect 5632 29232 5684 29238
rect 5632 29174 5684 29180
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4816 27470 4844 29038
rect 5632 28484 5684 28490
rect 5632 28426 5684 28432
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 5448 28008 5500 28014
rect 5448 27950 5500 27956
rect 4896 27600 4948 27606
rect 4896 27542 4948 27548
rect 4804 27464 4856 27470
rect 4804 27406 4856 27412
rect 4712 27056 4764 27062
rect 4712 26998 4764 27004
rect 4580 25792 4844 25820
rect 4528 25774 4580 25780
rect 4080 25294 4108 25774
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4620 24880 4672 24886
rect 4620 24822 4672 24828
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 23866 4660 24822
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4724 23866 4752 24142
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4620 23588 4672 23594
rect 4620 23530 4672 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 23180 4028 23186
rect 3976 23122 4028 23128
rect 3988 21554 4016 23122
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3988 19922 4016 21490
rect 4252 21480 4304 21486
rect 4250 21448 4252 21457
rect 4304 21448 4306 21457
rect 4250 21383 4306 21392
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 20868 4120 20874
rect 4068 20810 4120 20816
rect 3976 19916 4028 19922
rect 3976 19858 4028 19864
rect 3988 19378 4016 19858
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3988 18426 4016 19314
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3988 18290 4016 18362
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3988 17746 4016 18226
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 4080 17270 4108 20810
rect 4632 20398 4660 23530
rect 4712 21956 4764 21962
rect 4712 21898 4764 21904
rect 4724 21486 4752 21898
rect 4712 21480 4764 21486
rect 4712 21422 4764 21428
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18952 4660 20198
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4540 18924 4660 18952
rect 4160 18216 4212 18222
rect 4158 18184 4160 18193
rect 4540 18193 4568 18924
rect 4620 18624 4672 18630
rect 4620 18566 4672 18572
rect 4212 18184 4214 18193
rect 4158 18119 4214 18128
rect 4526 18184 4582 18193
rect 4526 18119 4582 18128
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4172 16980 4200 17478
rect 4264 17202 4292 17818
rect 4632 17746 4660 18566
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4080 16952 4200 16980
rect 4080 16708 4108 16952
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4080 16680 4200 16708
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3988 16153 4016 16526
rect 4172 16182 4200 16680
rect 4160 16176 4212 16182
rect 3974 16144 4030 16153
rect 4160 16118 4212 16124
rect 3974 16079 4030 16088
rect 4172 15892 4200 16118
rect 4080 15864 4200 15892
rect 4080 15586 4108 15864
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4080 15558 4200 15586
rect 4172 15434 4200 15558
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3804 12442 3832 14350
rect 4080 13938 4108 14554
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4172 13870 4200 14010
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13326 4660 17682
rect 4724 16046 4752 19722
rect 4816 17882 4844 25792
rect 4908 23662 4936 27542
rect 4896 23656 4948 23662
rect 4896 23598 4948 23604
rect 5000 21706 5028 27950
rect 5264 27464 5316 27470
rect 5264 27406 5316 27412
rect 5276 23730 5304 27406
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 5368 24274 5396 26726
rect 5460 26586 5488 27950
rect 5448 26580 5500 26586
rect 5448 26522 5500 26528
rect 5644 25226 5672 28426
rect 5632 25220 5684 25226
rect 5632 25162 5684 25168
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 5368 24154 5396 24210
rect 5368 24126 5488 24154
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4908 21690 5028 21706
rect 4908 21684 5040 21690
rect 4908 21678 4988 21684
rect 4908 21350 4936 21678
rect 4988 21626 5040 21632
rect 5000 21595 5028 21626
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4908 18222 4936 19450
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4896 17604 4948 17610
rect 4896 17546 4948 17552
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4724 14006 4752 14214
rect 4712 14000 4764 14006
rect 4712 13942 4764 13948
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 4632 12238 4660 13126
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4080 11354 4108 11562
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4724 11218 4752 13806
rect 4816 12918 4844 14282
rect 4908 12986 4936 17546
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4894 12880 4950 12889
rect 4894 12815 4950 12824
rect 4908 12714 4936 12815
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4908 12374 4936 12650
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4068 11144 4120 11150
rect 4252 11144 4304 11150
rect 4120 11104 4252 11132
rect 4068 11086 4120 11092
rect 4252 11086 4304 11092
rect 4816 10674 4844 12038
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4908 10130 4936 12038
rect 5000 11286 5028 21422
rect 5092 13818 5120 23598
rect 5276 23526 5304 23666
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 5356 23520 5408 23526
rect 5356 23462 5408 23468
rect 5276 23322 5304 23462
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 5264 22092 5316 22098
rect 5184 22052 5264 22080
rect 5184 21690 5212 22052
rect 5264 22034 5316 22040
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5276 21457 5304 21626
rect 5368 21554 5396 23462
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5262 21448 5318 21457
rect 5262 21383 5318 21392
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 16590 5212 19654
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5276 18426 5304 18566
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5276 15586 5304 18158
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 5368 15910 5396 17206
rect 5460 17202 5488 24126
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5552 23118 5580 23802
rect 5644 23118 5672 25162
rect 5736 23866 5764 34546
rect 6288 34474 6316 34546
rect 6276 34468 6328 34474
rect 6276 34410 6328 34416
rect 6458 34096 6514 34105
rect 6458 34031 6514 34040
rect 6184 33516 6236 33522
rect 6184 33458 6236 33464
rect 6196 32910 6224 33458
rect 6184 32904 6236 32910
rect 6182 32872 6184 32881
rect 6236 32872 6238 32881
rect 6182 32807 6238 32816
rect 6472 31822 6500 34031
rect 6840 33046 6868 36042
rect 7840 35488 7892 35494
rect 7840 35430 7892 35436
rect 7748 34944 7800 34950
rect 7748 34886 7800 34892
rect 7760 34610 7788 34886
rect 7748 34604 7800 34610
rect 7748 34546 7800 34552
rect 7852 33590 7880 35430
rect 7840 33584 7892 33590
rect 7840 33526 7892 33532
rect 7472 33448 7524 33454
rect 7472 33390 7524 33396
rect 6828 33040 6880 33046
rect 6828 32982 6880 32988
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 6552 32360 6604 32366
rect 6552 32302 6604 32308
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6000 31680 6052 31686
rect 6000 31622 6052 31628
rect 6012 31278 6040 31622
rect 6564 31482 6592 32302
rect 6840 32026 6868 32846
rect 6920 32768 6972 32774
rect 6920 32710 6972 32716
rect 6828 32020 6880 32026
rect 6828 31962 6880 31968
rect 6552 31476 6604 31482
rect 6552 31418 6604 31424
rect 6932 31346 6960 32710
rect 7484 32502 7512 33390
rect 7564 32768 7616 32774
rect 7564 32710 7616 32716
rect 7576 32570 7604 32710
rect 7564 32564 7616 32570
rect 7564 32506 7616 32512
rect 7472 32496 7524 32502
rect 7472 32438 7524 32444
rect 7484 31890 7512 32438
rect 7472 31884 7524 31890
rect 7472 31826 7524 31832
rect 7852 31822 7880 33526
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 7840 31816 7892 31822
rect 7840 31758 7892 31764
rect 6920 31340 6972 31346
rect 6920 31282 6972 31288
rect 6000 31272 6052 31278
rect 6000 31214 6052 31220
rect 6012 28626 6040 31214
rect 7116 30394 7144 31758
rect 7104 30388 7156 30394
rect 7104 30330 7156 30336
rect 6552 29096 6604 29102
rect 6552 29038 6604 29044
rect 6000 28620 6052 28626
rect 6000 28562 6052 28568
rect 6564 28558 6592 29038
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6000 28416 6052 28422
rect 6000 28358 6052 28364
rect 6012 28150 6040 28358
rect 6000 28144 6052 28150
rect 6000 28086 6052 28092
rect 6564 28082 6592 28494
rect 6552 28076 6604 28082
rect 7116 28064 7144 30330
rect 7116 28036 7420 28064
rect 6552 28018 6604 28024
rect 7012 27328 7064 27334
rect 7012 27270 7064 27276
rect 6092 26376 6144 26382
rect 6092 26318 6144 26324
rect 6104 25838 6132 26318
rect 7024 26314 7052 27270
rect 6644 26308 6696 26314
rect 6644 26250 6696 26256
rect 7012 26308 7064 26314
rect 7012 26250 7064 26256
rect 6092 25832 6144 25838
rect 6092 25774 6144 25780
rect 6104 25362 6132 25774
rect 6656 25702 6684 26250
rect 6644 25696 6696 25702
rect 6644 25638 6696 25644
rect 6092 25356 6144 25362
rect 6092 25298 6144 25304
rect 6368 25220 6420 25226
rect 6368 25162 6420 25168
rect 6380 25129 6408 25162
rect 6366 25120 6422 25129
rect 6366 25055 6422 25064
rect 5724 23860 5776 23866
rect 5724 23802 5776 23808
rect 5736 23730 5764 23802
rect 5724 23724 5776 23730
rect 5724 23666 5776 23672
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5632 23112 5684 23118
rect 5632 23054 5684 23060
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 5552 21962 5580 22918
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 5724 21344 5776 21350
rect 5724 21286 5776 21292
rect 5736 19990 5764 21286
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5552 18630 5580 19858
rect 5632 18692 5684 18698
rect 5632 18634 5684 18640
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5552 16590 5580 17138
rect 5644 16658 5672 18634
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5540 16584 5592 16590
rect 5736 16538 5764 19926
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5828 17762 5856 19314
rect 6012 19310 6040 21422
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 18426 6040 19110
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5828 17734 5948 17762
rect 5816 17604 5868 17610
rect 5816 17546 5868 17552
rect 5540 16526 5592 16532
rect 5644 16510 5764 16538
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5184 15558 5304 15586
rect 5184 13938 5212 15558
rect 5264 15428 5316 15434
rect 5264 15370 5316 15376
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5276 14618 5304 15370
rect 5368 15162 5396 15370
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5368 14074 5396 15098
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5356 13864 5408 13870
rect 5092 13790 5304 13818
rect 5356 13806 5408 13812
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 5092 13326 5120 13670
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5276 12434 5304 13790
rect 5184 12406 5304 12434
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 5092 10062 5120 12106
rect 5184 12102 5212 12406
rect 5368 12322 5396 13806
rect 5460 13802 5488 15982
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 12782 5488 13738
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5552 12628 5580 15846
rect 5644 14414 5672 16510
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 15094 5764 16390
rect 5828 15502 5856 17546
rect 5920 16590 5948 17734
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5920 16182 5948 16390
rect 5908 16176 5960 16182
rect 5908 16118 5960 16124
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5920 14618 5948 14894
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5632 14408 5684 14414
rect 5684 14368 5856 14396
rect 5632 14350 5684 14356
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5276 12294 5396 12322
rect 5460 12600 5580 12628
rect 5276 12238 5304 12294
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5184 10470 5212 11630
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3804 8430 3832 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5000 8974 5028 9862
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4632 8498 4660 8774
rect 5184 8634 5212 10406
rect 5276 9586 5304 12174
rect 5460 11642 5488 12600
rect 5736 12306 5764 13874
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5644 11694 5672 11834
rect 5368 11614 5488 11642
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5368 11218 5396 11614
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5460 11082 5488 11494
rect 5644 11354 5672 11630
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5368 10810 5396 11018
rect 5552 10962 5580 11154
rect 5460 10934 5580 10962
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3988 3194 4016 7822
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5114 4660 7142
rect 5460 5710 5488 10934
rect 5828 9450 5856 14368
rect 6012 13938 6040 18362
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 6104 16726 6132 18226
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 6104 16590 6132 16662
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6104 15910 6132 16050
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6104 12306 6132 13126
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 10674 6040 12038
rect 6196 11830 6224 16730
rect 6288 16726 6316 20742
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6472 18630 6500 19246
rect 6564 18970 6592 23666
rect 6656 20262 6684 25638
rect 7104 25152 7156 25158
rect 6826 25120 6882 25129
rect 7104 25094 7156 25100
rect 6826 25055 6882 25064
rect 6840 24698 6868 25055
rect 6840 24670 6960 24698
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 6840 24410 6868 24550
rect 6932 24410 6960 24670
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6748 23118 6776 24074
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6748 20534 6776 23054
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6828 22092 6880 22098
rect 6932 22080 6960 22578
rect 6880 22052 6960 22080
rect 6828 22034 6880 22040
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6840 20942 6868 21422
rect 6932 21146 6960 22052
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6840 20806 6868 20878
rect 7024 20874 7052 22918
rect 7116 22574 7144 25094
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6840 19718 6868 20742
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6380 11694 6408 18566
rect 6564 18290 6592 18906
rect 6840 18766 6868 19654
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6840 18222 6868 18702
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6460 18148 6512 18154
rect 6460 18090 6512 18096
rect 6472 17542 6500 18090
rect 7024 17882 7052 19858
rect 7116 18358 7144 22510
rect 7196 21616 7248 21622
rect 7196 21558 7248 21564
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6472 11762 6500 17478
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 6564 16794 6592 17206
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6564 15502 6592 16730
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6564 14346 6592 14554
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6564 12850 6592 14282
rect 6656 12918 6684 16934
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6840 14890 6868 15030
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6932 14346 6960 16390
rect 7024 15586 7052 17818
rect 7104 17604 7156 17610
rect 7104 17546 7156 17552
rect 7116 17338 7144 17546
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7208 16250 7236 21558
rect 7300 18306 7328 23598
rect 7392 21690 7420 28036
rect 7932 26444 7984 26450
rect 7932 26386 7984 26392
rect 7472 25832 7524 25838
rect 7472 25774 7524 25780
rect 7484 24274 7512 25774
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7472 24268 7524 24274
rect 7472 24210 7524 24216
rect 7484 23730 7512 24210
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7484 22642 7512 23666
rect 7760 23662 7788 24754
rect 7748 23656 7800 23662
rect 7748 23598 7800 23604
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7380 20868 7432 20874
rect 7380 20810 7432 20816
rect 7392 19394 7420 20810
rect 7484 19514 7512 22170
rect 7576 21690 7604 22918
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 7576 21486 7604 21626
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7760 20058 7788 20198
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7392 19366 7604 19394
rect 7472 18352 7524 18358
rect 7300 18278 7420 18306
rect 7472 18294 7524 18300
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7300 17746 7328 18158
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7024 15558 7144 15586
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6828 13864 6880 13870
rect 6748 13824 6828 13852
rect 6748 13530 6776 13824
rect 6828 13806 6880 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6840 13258 6868 13670
rect 7024 13512 7052 15370
rect 7116 13938 7144 15558
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7208 13530 7236 15914
rect 7288 15018 7340 15024
rect 7288 14960 7340 14966
rect 7300 14328 7328 14960
rect 7392 14482 7420 18278
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7380 14340 7432 14346
rect 7300 14300 7380 14328
rect 7300 14249 7328 14300
rect 7380 14282 7432 14288
rect 7286 14240 7342 14249
rect 7286 14175 7342 14184
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 6932 13484 7052 13512
rect 7196 13524 7248 13530
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6932 12594 6960 13484
rect 7196 13466 7248 13472
rect 7300 13462 7328 14010
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6656 12566 6960 12594
rect 6552 12436 6604 12442
rect 6656 12434 6684 12566
rect 6656 12406 6960 12434
rect 6552 12378 6604 12384
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6564 11354 6592 12378
rect 6932 11778 6960 12406
rect 7024 11898 7052 13330
rect 7484 13190 7512 18294
rect 7576 17542 7604 19366
rect 7656 18216 7708 18222
rect 7852 18170 7880 19654
rect 7708 18164 7880 18170
rect 7656 18158 7880 18164
rect 7668 18142 7880 18158
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12434 7512 13126
rect 7392 12406 7512 12434
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6932 11750 7052 11778
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6472 9586 6500 11018
rect 6564 9586 6592 11290
rect 7024 10742 7052 11750
rect 7116 10742 7144 12038
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7208 11014 7236 11494
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7024 10470 7052 10678
rect 7300 10606 7328 11562
rect 7392 11150 7420 12406
rect 7576 12374 7604 17478
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7668 15434 7696 16390
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 7654 15328 7710 15337
rect 7654 15263 7710 15272
rect 7668 15026 7696 15263
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7668 13870 7696 14350
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7760 12170 7788 18142
rect 7944 17202 7972 26386
rect 8036 25362 8064 37062
rect 9048 36786 9076 39200
rect 9692 37262 9720 39200
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 10980 37210 11008 39200
rect 12268 37330 12296 39200
rect 12256 37324 12308 37330
rect 12256 37266 12308 37272
rect 10980 37182 11100 37210
rect 13556 37194 13584 39200
rect 14200 37262 14228 39200
rect 14004 37256 14056 37262
rect 14004 37198 14056 37204
rect 14188 37256 14240 37262
rect 14188 37198 14240 37204
rect 11072 37126 11100 37182
rect 13544 37188 13596 37194
rect 13544 37130 13596 37136
rect 9496 37120 9548 37126
rect 9496 37062 9548 37068
rect 10876 37120 10928 37126
rect 10876 37062 10928 37068
rect 11060 37120 11112 37126
rect 11060 37062 11112 37068
rect 9310 36816 9366 36825
rect 9036 36780 9088 36786
rect 9310 36751 9366 36760
rect 9036 36722 9088 36728
rect 8668 36712 8720 36718
rect 8668 36654 8720 36660
rect 8680 36378 8708 36654
rect 9128 36576 9180 36582
rect 9128 36518 9180 36524
rect 8668 36372 8720 36378
rect 8668 36314 8720 36320
rect 9140 36310 9168 36518
rect 8116 36304 8168 36310
rect 8116 36246 8168 36252
rect 9128 36304 9180 36310
rect 9128 36246 9180 36252
rect 8128 33998 8156 36246
rect 9140 36106 9168 36246
rect 9128 36100 9180 36106
rect 9128 36042 9180 36048
rect 9324 35766 9352 36751
rect 9312 35760 9364 35766
rect 9312 35702 9364 35708
rect 8208 35148 8260 35154
rect 8208 35090 8260 35096
rect 8220 34202 8248 35090
rect 9508 35057 9536 37062
rect 10888 36922 10916 37062
rect 10140 36916 10192 36922
rect 10140 36858 10192 36864
rect 10876 36916 10928 36922
rect 10876 36858 10928 36864
rect 12900 36916 12952 36922
rect 12900 36858 12952 36864
rect 13912 36916 13964 36922
rect 13912 36858 13964 36864
rect 9588 36236 9640 36242
rect 9640 36196 9996 36224
rect 9588 36178 9640 36184
rect 9968 36106 9996 36196
rect 9772 36100 9824 36106
rect 9772 36042 9824 36048
rect 9956 36100 10008 36106
rect 9956 36042 10008 36048
rect 9784 35290 9812 36042
rect 9588 35284 9640 35290
rect 9588 35226 9640 35232
rect 9772 35284 9824 35290
rect 9772 35226 9824 35232
rect 9494 35048 9550 35057
rect 9494 34983 9550 34992
rect 9600 34610 9628 35226
rect 9588 34604 9640 34610
rect 9588 34546 9640 34552
rect 8208 34196 8260 34202
rect 8208 34138 8260 34144
rect 8116 33992 8168 33998
rect 8116 33934 8168 33940
rect 8220 33454 8248 34138
rect 8944 34060 8996 34066
rect 8944 34002 8996 34008
rect 8208 33448 8260 33454
rect 8208 33390 8260 33396
rect 8956 32910 8984 34002
rect 9404 33448 9456 33454
rect 9404 33390 9456 33396
rect 8944 32904 8996 32910
rect 8944 32846 8996 32852
rect 8956 32434 8984 32846
rect 8300 32428 8352 32434
rect 8300 32370 8352 32376
rect 8944 32428 8996 32434
rect 8944 32370 8996 32376
rect 8312 31414 8340 32370
rect 8956 31822 8984 32370
rect 8944 31816 8996 31822
rect 8944 31758 8996 31764
rect 8300 31408 8352 31414
rect 8300 31350 8352 31356
rect 9220 26920 9272 26926
rect 9220 26862 9272 26868
rect 8024 25356 8076 25362
rect 8024 25298 8076 25304
rect 8116 24064 8168 24070
rect 8116 24006 8168 24012
rect 8128 22166 8156 24006
rect 9232 23866 9260 26862
rect 9416 24410 9444 33390
rect 10152 31142 10180 36858
rect 11980 36848 12032 36854
rect 11980 36790 12032 36796
rect 10416 36712 10468 36718
rect 10416 36654 10468 36660
rect 10324 36576 10376 36582
rect 10324 36518 10376 36524
rect 10336 36281 10364 36518
rect 10322 36272 10378 36281
rect 10232 36236 10284 36242
rect 10428 36242 10456 36654
rect 11888 36644 11940 36650
rect 11888 36586 11940 36592
rect 10322 36207 10378 36216
rect 10416 36236 10468 36242
rect 10232 36178 10284 36184
rect 10416 36178 10468 36184
rect 10244 35601 10272 36178
rect 11900 36174 11928 36586
rect 11992 36242 12020 36790
rect 12440 36712 12492 36718
rect 12440 36654 12492 36660
rect 11980 36236 12032 36242
rect 11980 36178 12032 36184
rect 10876 36168 10928 36174
rect 10876 36110 10928 36116
rect 11888 36168 11940 36174
rect 11888 36110 11940 36116
rect 10888 35834 10916 36110
rect 11060 36032 11112 36038
rect 11060 35974 11112 35980
rect 11520 36032 11572 36038
rect 11520 35974 11572 35980
rect 11612 36032 11664 36038
rect 11612 35974 11664 35980
rect 10876 35828 10928 35834
rect 10876 35770 10928 35776
rect 10230 35592 10286 35601
rect 10230 35527 10286 35536
rect 10244 32842 10272 35527
rect 10508 35080 10560 35086
rect 10508 35022 10560 35028
rect 10520 34746 10548 35022
rect 10508 34740 10560 34746
rect 10508 34682 10560 34688
rect 11072 34066 11100 35974
rect 11532 35698 11560 35974
rect 11520 35692 11572 35698
rect 11520 35634 11572 35640
rect 11060 34060 11112 34066
rect 11060 34002 11112 34008
rect 11072 33969 11100 34002
rect 11058 33960 11114 33969
rect 10324 33924 10376 33930
rect 10324 33866 10376 33872
rect 10600 33924 10652 33930
rect 11058 33895 11114 33904
rect 11334 33960 11390 33969
rect 11334 33895 11390 33904
rect 10600 33866 10652 33872
rect 10232 32836 10284 32842
rect 10232 32778 10284 32784
rect 10232 32224 10284 32230
rect 10232 32166 10284 32172
rect 10244 31890 10272 32166
rect 10336 31958 10364 33866
rect 10612 33658 10640 33866
rect 10600 33652 10652 33658
rect 10600 33594 10652 33600
rect 10692 32224 10744 32230
rect 10692 32166 10744 32172
rect 10324 31952 10376 31958
rect 10324 31894 10376 31900
rect 10232 31884 10284 31890
rect 10232 31826 10284 31832
rect 10244 31686 10272 31826
rect 10232 31680 10284 31686
rect 10232 31622 10284 31628
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 9876 30598 9904 31078
rect 9864 30592 9916 30598
rect 9864 30534 9916 30540
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9692 28762 9720 28902
rect 9680 28756 9732 28762
rect 9680 28698 9732 28704
rect 9956 27872 10008 27878
rect 9956 27814 10008 27820
rect 9968 25838 9996 27814
rect 9956 25832 10008 25838
rect 9956 25774 10008 25780
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9128 23520 9180 23526
rect 9128 23462 9180 23468
rect 8208 22228 8260 22234
rect 8208 22170 8260 22176
rect 8116 22160 8168 22166
rect 8116 22102 8168 22108
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 8024 21684 8076 21690
rect 8024 21626 8076 21632
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 8036 15450 8064 21626
rect 8128 16658 8156 21830
rect 8220 21690 8248 22170
rect 8392 22024 8444 22030
rect 8390 21992 8392 22001
rect 8444 21992 8446 22001
rect 8390 21927 8446 21936
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8484 21480 8536 21486
rect 8484 21422 8536 21428
rect 8496 20806 8524 21422
rect 8772 21350 8800 21830
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8576 20868 8628 20874
rect 8576 20810 8628 20816
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8496 20534 8524 20742
rect 8484 20528 8536 20534
rect 8484 20470 8536 20476
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8220 16250 8248 18702
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8312 16046 8340 18294
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8404 16658 8432 17070
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8404 15706 8432 15982
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 7944 15422 8064 15450
rect 7944 14618 7972 15422
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8036 13870 8064 15302
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 14074 8156 14758
rect 8220 14618 8248 14894
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7852 11762 7880 13806
rect 8312 12986 8340 15030
rect 8496 14958 8524 17002
rect 8588 15434 8616 20810
rect 8680 18766 8708 21286
rect 8956 20942 8984 21830
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8944 19440 8996 19446
rect 8944 19382 8996 19388
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8404 13326 8432 13806
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8312 12782 8340 12922
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8128 12434 8156 12582
rect 8128 12406 8248 12434
rect 8220 12170 8248 12406
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 8312 11558 8340 12310
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7852 10674 7880 11222
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 8974 6684 9318
rect 6840 9178 6868 9998
rect 8220 9654 8248 11018
rect 8312 10538 8340 11494
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5234 4752 5510
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4632 5086 4752 5114
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4632 3126 4660 4966
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4724 2514 4752 5086
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 3896 800 3924 2246
rect 5184 800 5212 2246
rect 6472 800 6500 2382
rect 6840 2378 6868 7686
rect 7116 2650 7144 9454
rect 8404 2774 8432 13262
rect 8680 13190 8708 18702
rect 8956 18426 8984 19382
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8760 16516 8812 16522
rect 8760 16458 8812 16464
rect 8772 16153 8800 16458
rect 8758 16144 8814 16153
rect 8758 16079 8760 16088
rect 8812 16079 8814 16088
rect 8760 16050 8812 16056
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8496 12306 8524 13126
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8496 11558 8524 11766
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8496 10198 8524 10542
rect 8864 10266 8892 12174
rect 9140 11898 9168 23462
rect 9232 18290 9260 23802
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9508 22574 9536 22986
rect 9600 22710 9628 23054
rect 9588 22704 9640 22710
rect 9588 22646 9640 22652
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9600 20942 9628 22646
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 9876 21146 9904 21558
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9600 17241 9628 20878
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9692 17882 9720 20470
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9784 19514 9812 20198
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9680 17264 9732 17270
rect 9586 17232 9642 17241
rect 9680 17206 9732 17212
rect 9586 17167 9642 17176
rect 9600 16794 9628 17167
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9692 16250 9720 17206
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9678 16144 9734 16153
rect 9678 16079 9680 16088
rect 9732 16079 9734 16088
rect 9680 16050 9732 16056
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15502 9720 15846
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9784 15026 9812 17070
rect 9876 15366 9904 18566
rect 9968 18358 9996 18906
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 10060 18222 10088 18906
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10060 17746 10088 18158
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10152 16998 10180 20334
rect 10140 16992 10192 16998
rect 9968 16952 10140 16980
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9862 14920 9918 14929
rect 9862 14855 9864 14864
rect 9916 14855 9918 14864
rect 9864 14826 9916 14832
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 14346 9444 14758
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9784 13258 9812 13670
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9416 11626 9444 12106
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9508 11218 9536 12242
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9600 11744 9628 11834
rect 9772 11756 9824 11762
rect 9600 11716 9772 11744
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9600 11150 9628 11716
rect 9772 11698 9824 11704
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8496 9450 8524 10134
rect 9140 10130 9168 11086
rect 9324 10810 9352 11086
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9692 10742 9720 10950
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9876 10062 9904 14010
rect 9968 13938 9996 16952
rect 10140 16934 10192 16940
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10152 15434 10180 16390
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 10060 14940 10088 15370
rect 10244 15094 10272 15846
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10232 14952 10284 14958
rect 10060 14912 10232 14940
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9968 12850 9996 13194
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 10060 12764 10088 14912
rect 10232 14894 10284 14900
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10244 13394 10272 14282
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10140 12912 10192 12918
rect 10192 12860 10272 12866
rect 10140 12854 10272 12860
rect 10152 12838 10272 12854
rect 10060 12736 10180 12764
rect 10046 12608 10102 12617
rect 10046 12543 10102 12552
rect 10060 11286 10088 12543
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9654 9260 9862
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 10152 9178 10180 12736
rect 10244 11898 10272 12838
rect 10336 12374 10364 31894
rect 10704 31278 10732 32166
rect 11348 31754 11376 33895
rect 11428 33856 11480 33862
rect 11428 33798 11480 33804
rect 11440 32910 11468 33798
rect 11428 32904 11480 32910
rect 11428 32846 11480 32852
rect 11440 32745 11468 32846
rect 11624 32842 11652 35974
rect 12452 35630 12480 36654
rect 12912 36310 12940 36858
rect 12992 36712 13044 36718
rect 12992 36654 13044 36660
rect 13004 36310 13032 36654
rect 12900 36304 12952 36310
rect 12900 36246 12952 36252
rect 12992 36304 13044 36310
rect 12992 36246 13044 36252
rect 13544 36168 13596 36174
rect 13544 36110 13596 36116
rect 13556 36009 13584 36110
rect 13542 36000 13598 36009
rect 13542 35935 13598 35944
rect 12440 35624 12492 35630
rect 12440 35566 12492 35572
rect 12808 35624 12860 35630
rect 12808 35566 12860 35572
rect 12256 35488 12308 35494
rect 12256 35430 12308 35436
rect 12268 35222 12296 35430
rect 12256 35216 12308 35222
rect 12256 35158 12308 35164
rect 12452 35154 12480 35566
rect 12532 35488 12584 35494
rect 12532 35430 12584 35436
rect 12544 35290 12572 35430
rect 12532 35284 12584 35290
rect 12532 35226 12584 35232
rect 12440 35148 12492 35154
rect 12440 35090 12492 35096
rect 12624 34944 12676 34950
rect 12624 34886 12676 34892
rect 12716 34944 12768 34950
rect 12716 34886 12768 34892
rect 12636 34610 12664 34886
rect 12728 34610 12756 34886
rect 12440 34604 12492 34610
rect 12440 34546 12492 34552
rect 12624 34604 12676 34610
rect 12624 34546 12676 34552
rect 12716 34604 12768 34610
rect 12716 34546 12768 34552
rect 11704 33856 11756 33862
rect 11704 33798 11756 33804
rect 11716 33522 11744 33798
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 11612 32836 11664 32842
rect 11612 32778 11664 32784
rect 11426 32736 11482 32745
rect 11426 32671 11482 32680
rect 11796 31816 11848 31822
rect 11796 31758 11848 31764
rect 11152 31748 11204 31754
rect 11348 31726 11468 31754
rect 11152 31690 11204 31696
rect 10968 31680 11020 31686
rect 11020 31628 11100 31634
rect 10968 31622 11100 31628
rect 10980 31606 11100 31622
rect 10692 31272 10744 31278
rect 10692 31214 10744 31220
rect 11072 29238 11100 31606
rect 11164 30802 11192 31690
rect 11244 31680 11296 31686
rect 11244 31622 11296 31628
rect 11256 31210 11284 31622
rect 11244 31204 11296 31210
rect 11244 31146 11296 31152
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11060 29232 11112 29238
rect 11060 29174 11112 29180
rect 11244 29096 11296 29102
rect 11244 29038 11296 29044
rect 11152 29028 11204 29034
rect 11152 28970 11204 28976
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10520 26314 10548 27338
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 10508 26308 10560 26314
rect 10508 26250 10560 26256
rect 10782 26208 10838 26217
rect 10782 26143 10838 26152
rect 10796 26042 10824 26143
rect 10784 26036 10836 26042
rect 10784 25978 10836 25984
rect 11072 25226 11100 26726
rect 11164 26314 11192 28970
rect 11256 28558 11284 29038
rect 11244 28552 11296 28558
rect 11244 28494 11296 28500
rect 11256 26994 11284 28494
rect 11244 26988 11296 26994
rect 11244 26930 11296 26936
rect 11152 26308 11204 26314
rect 11152 26250 11204 26256
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10796 22778 10824 22986
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 10428 21010 10456 21830
rect 10704 21486 10732 22714
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 10416 20528 10468 20534
rect 10416 20470 10468 20476
rect 10428 16250 10456 20470
rect 10520 19802 10548 20878
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10612 19922 10640 20198
rect 10796 20074 10824 20538
rect 10980 20398 11008 20878
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10704 20058 10824 20074
rect 10692 20052 10824 20058
rect 10744 20046 10824 20052
rect 10692 19994 10744 20000
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10520 19774 10640 19802
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10520 15706 10548 17546
rect 10612 16402 10640 19774
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 16590 10732 17478
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10612 16374 10732 16402
rect 10704 15978 10732 16374
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10704 15638 10732 15914
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10428 15201 10456 15302
rect 10414 15192 10470 15201
rect 10414 15127 10470 15136
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10428 11762 10456 15127
rect 10796 13938 10824 17818
rect 10888 17134 10916 20198
rect 10980 19922 11008 20334
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 10980 19802 11008 19858
rect 10980 19774 11100 19802
rect 11072 19310 11100 19774
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11072 18766 11100 19246
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 17338 11100 18702
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 10966 17232 11022 17241
rect 10966 17167 10968 17176
rect 11020 17167 11022 17176
rect 10968 17138 11020 17144
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11072 16114 11100 17070
rect 11164 16998 11192 18022
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 14414 11100 16050
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10520 12782 10548 13330
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10704 12986 10732 13194
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10520 12617 10548 12718
rect 10612 12714 10640 12922
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10506 12608 10562 12617
rect 10506 12543 10562 12552
rect 10980 12434 11008 13874
rect 10796 12406 11008 12434
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10428 9654 10456 11018
rect 10796 11014 10824 12406
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10888 10810 10916 12106
rect 11164 11694 11192 16934
rect 11256 16250 11284 23598
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 11348 19786 11376 20742
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11348 18086 11376 18770
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11440 15094 11468 31726
rect 11808 31346 11836 31758
rect 12452 31414 12480 34546
rect 12532 33924 12584 33930
rect 12532 33866 12584 33872
rect 12348 31408 12400 31414
rect 12348 31350 12400 31356
rect 12440 31408 12492 31414
rect 12440 31350 12492 31356
rect 11796 31340 11848 31346
rect 11796 31282 11848 31288
rect 11612 30184 11664 30190
rect 11612 30126 11664 30132
rect 11624 29646 11652 30126
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11624 29102 11652 29582
rect 11796 29572 11848 29578
rect 11796 29514 11848 29520
rect 11612 29096 11664 29102
rect 11612 29038 11664 29044
rect 11612 28484 11664 28490
rect 11612 28426 11664 28432
rect 11520 27328 11572 27334
rect 11520 27270 11572 27276
rect 11532 24138 11560 27270
rect 11624 26217 11652 28426
rect 11610 26208 11666 26217
rect 11610 26143 11666 26152
rect 11520 24132 11572 24138
rect 11520 24074 11572 24080
rect 11704 23044 11756 23050
rect 11704 22986 11756 22992
rect 11520 22092 11572 22098
rect 11716 22094 11744 22986
rect 11520 22034 11572 22040
rect 11624 22066 11744 22094
rect 11532 21962 11560 22034
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11532 15434 11560 16390
rect 11624 16114 11652 22066
rect 11808 22030 11836 29514
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 12268 25906 12296 26386
rect 12256 25900 12308 25906
rect 12256 25842 12308 25848
rect 12268 24274 12296 25842
rect 12256 24268 12308 24274
rect 12256 24210 12308 24216
rect 11888 24132 11940 24138
rect 11888 24074 11940 24080
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 11796 21412 11848 21418
rect 11796 21354 11848 21360
rect 11704 20868 11756 20874
rect 11704 20810 11756 20816
rect 11716 18426 11744 20810
rect 11808 20346 11836 21354
rect 11900 20534 11928 24074
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 12084 20466 12112 23666
rect 12268 23186 12296 24210
rect 12256 23180 12308 23186
rect 12256 23122 12308 23128
rect 12256 23044 12308 23050
rect 12256 22986 12308 22992
rect 12268 22642 12296 22986
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12164 22228 12216 22234
rect 12164 22170 12216 22176
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 11808 20318 12112 20346
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 11624 15366 11652 15914
rect 11716 15366 11744 16390
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10968 11552 11020 11558
rect 11152 11552 11204 11558
rect 11020 11500 11100 11506
rect 10968 11494 11100 11500
rect 11152 11494 11204 11500
rect 10980 11478 11100 11494
rect 11072 11354 11100 11478
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11164 11082 11192 11494
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9140 7954 9168 8910
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9140 7410 9168 7890
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8404 2746 8524 2774
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 8496 2514 8524 2746
rect 10244 2650 10272 9522
rect 11072 9518 11100 11018
rect 11256 10674 11284 13738
rect 11348 11830 11376 13874
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11348 10470 11376 11154
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11164 2922 11192 9998
rect 11440 9994 11468 12718
rect 11624 12434 11652 15302
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11716 14414 11744 15098
rect 11808 14618 11836 18634
rect 11900 17270 11928 19858
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11992 17338 12020 17614
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11900 16182 11928 17206
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11900 15434 11928 16118
rect 12084 15910 12112 20318
rect 12176 19310 12204 22170
rect 12360 22094 12388 31350
rect 12544 28694 12572 33866
rect 12716 32020 12768 32026
rect 12716 31962 12768 31968
rect 12532 28688 12584 28694
rect 12532 28630 12584 28636
rect 12728 28642 12756 31962
rect 12820 31754 12848 35566
rect 13358 35184 13414 35193
rect 13176 35148 13228 35154
rect 13358 35119 13360 35128
rect 13176 35090 13228 35096
rect 13412 35119 13414 35128
rect 13360 35090 13412 35096
rect 13188 34406 13216 35090
rect 13268 35080 13320 35086
rect 13268 35022 13320 35028
rect 13280 34678 13308 35022
rect 13268 34672 13320 34678
rect 13268 34614 13320 34620
rect 13176 34400 13228 34406
rect 13176 34342 13228 34348
rect 13188 34048 13216 34342
rect 13728 34196 13780 34202
rect 13728 34138 13780 34144
rect 13268 34060 13320 34066
rect 13188 34020 13268 34048
rect 13188 33522 13216 34020
rect 13268 34002 13320 34008
rect 13740 33590 13768 34138
rect 13728 33584 13780 33590
rect 13728 33526 13780 33532
rect 13176 33516 13228 33522
rect 13176 33458 13228 33464
rect 13084 32768 13136 32774
rect 13084 32710 13136 32716
rect 13096 32502 13124 32710
rect 13084 32496 13136 32502
rect 13084 32438 13136 32444
rect 13544 32496 13596 32502
rect 13544 32438 13596 32444
rect 12820 31726 13032 31754
rect 13004 30122 13032 31726
rect 13452 30252 13504 30258
rect 13452 30194 13504 30200
rect 13464 30122 13492 30194
rect 12992 30116 13044 30122
rect 12992 30058 13044 30064
rect 13452 30116 13504 30122
rect 13452 30058 13504 30064
rect 12728 28614 13032 28642
rect 13004 28422 13032 28614
rect 12532 28416 12584 28422
rect 12532 28358 12584 28364
rect 12992 28416 13044 28422
rect 12992 28358 13044 28364
rect 12544 25820 12572 28358
rect 12808 28076 12860 28082
rect 12808 28018 12860 28024
rect 12820 27538 12848 28018
rect 13004 27674 13032 28358
rect 12992 27668 13044 27674
rect 12992 27610 13044 27616
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 13004 26586 13032 27270
rect 13556 27044 13584 32438
rect 13726 32056 13782 32065
rect 13726 31991 13782 32000
rect 13740 29578 13768 31991
rect 13924 31210 13952 36858
rect 14016 36378 14044 37198
rect 15488 37126 15516 39200
rect 15568 37256 15620 37262
rect 15568 37198 15620 37204
rect 14096 37120 14148 37126
rect 14096 37062 14148 37068
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 14924 37120 14976 37126
rect 14924 37062 14976 37068
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 14004 36372 14056 36378
rect 14004 36314 14056 36320
rect 14004 33448 14056 33454
rect 14004 33390 14056 33396
rect 14016 33046 14044 33390
rect 14004 33040 14056 33046
rect 14004 32982 14056 32988
rect 13912 31204 13964 31210
rect 13912 31146 13964 31152
rect 13912 30048 13964 30054
rect 13912 29990 13964 29996
rect 13728 29572 13780 29578
rect 13728 29514 13780 29520
rect 13924 29306 13952 29990
rect 14016 29782 14044 32982
rect 14004 29776 14056 29782
rect 14004 29718 14056 29724
rect 13912 29300 13964 29306
rect 13912 29242 13964 29248
rect 14108 28762 14136 37062
rect 14292 36038 14320 37062
rect 14936 36922 14964 37062
rect 14832 36916 14884 36922
rect 14832 36858 14884 36864
rect 14924 36916 14976 36922
rect 14924 36858 14976 36864
rect 14844 36802 14872 36858
rect 15028 36802 15056 37062
rect 14844 36774 15056 36802
rect 15016 36576 15068 36582
rect 15016 36518 15068 36524
rect 14646 36136 14702 36145
rect 14646 36071 14648 36080
rect 14700 36071 14702 36080
rect 14648 36042 14700 36048
rect 14280 36032 14332 36038
rect 14280 35974 14332 35980
rect 14648 35624 14700 35630
rect 14648 35566 14700 35572
rect 14188 35488 14240 35494
rect 14188 35430 14240 35436
rect 14200 34241 14228 35430
rect 14660 35154 14688 35566
rect 14648 35148 14700 35154
rect 14648 35090 14700 35096
rect 14372 34672 14424 34678
rect 14372 34614 14424 34620
rect 14186 34232 14242 34241
rect 14186 34167 14242 34176
rect 14200 32978 14228 34167
rect 14384 33114 14412 34614
rect 14660 34406 14688 35090
rect 14832 35012 14884 35018
rect 14832 34954 14884 34960
rect 14844 34649 14872 34954
rect 14830 34640 14886 34649
rect 14830 34575 14886 34584
rect 14648 34400 14700 34406
rect 14648 34342 14700 34348
rect 14660 34066 14688 34342
rect 14648 34060 14700 34066
rect 14648 34002 14700 34008
rect 14372 33108 14424 33114
rect 14372 33050 14424 33056
rect 14188 32972 14240 32978
rect 14188 32914 14240 32920
rect 15028 30122 15056 36518
rect 15580 36242 15608 37198
rect 16776 36854 16804 39200
rect 17420 37126 17448 39200
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 17868 37256 17920 37262
rect 18708 37210 18736 39200
rect 17868 37198 17920 37204
rect 17224 37120 17276 37126
rect 17224 37062 17276 37068
rect 17408 37120 17460 37126
rect 17408 37062 17460 37068
rect 16764 36848 16816 36854
rect 16764 36790 16816 36796
rect 17236 36718 17264 37062
rect 17408 36848 17460 36854
rect 17408 36790 17460 36796
rect 16764 36712 16816 36718
rect 16764 36654 16816 36660
rect 17224 36712 17276 36718
rect 17420 36689 17448 36790
rect 17224 36654 17276 36660
rect 17406 36680 17462 36689
rect 16580 36644 16632 36650
rect 16580 36586 16632 36592
rect 16672 36644 16724 36650
rect 16672 36586 16724 36592
rect 16396 36304 16448 36310
rect 16396 36246 16448 36252
rect 15568 36236 15620 36242
rect 15568 36178 15620 36184
rect 15568 36100 15620 36106
rect 15568 36042 15620 36048
rect 15580 34746 15608 36042
rect 16408 35222 16436 36246
rect 16592 35329 16620 36586
rect 16578 35320 16634 35329
rect 16578 35255 16634 35264
rect 16396 35216 16448 35222
rect 16396 35158 16448 35164
rect 15568 34740 15620 34746
rect 15568 34682 15620 34688
rect 15580 34082 15608 34682
rect 16304 34468 16356 34474
rect 16304 34410 16356 34416
rect 15844 34400 15896 34406
rect 15844 34342 15896 34348
rect 16026 34368 16082 34377
rect 15856 34134 15884 34342
rect 16026 34303 16082 34312
rect 15844 34128 15896 34134
rect 15580 34054 15792 34082
rect 15844 34070 15896 34076
rect 15384 33992 15436 33998
rect 15384 33934 15436 33940
rect 15108 33380 15160 33386
rect 15108 33322 15160 33328
rect 15120 32774 15148 33322
rect 15396 32842 15424 33934
rect 15660 33312 15712 33318
rect 15660 33254 15712 33260
rect 15384 32836 15436 32842
rect 15384 32778 15436 32784
rect 15108 32768 15160 32774
rect 15108 32710 15160 32716
rect 15292 32768 15344 32774
rect 15292 32710 15344 32716
rect 15304 32502 15332 32710
rect 15292 32496 15344 32502
rect 15292 32438 15344 32444
rect 15396 31958 15424 32778
rect 15672 32434 15700 33254
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 15384 31952 15436 31958
rect 15384 31894 15436 31900
rect 15396 31346 15424 31894
rect 15384 31340 15436 31346
rect 15384 31282 15436 31288
rect 15764 30870 15792 34054
rect 16040 33862 16068 34303
rect 16212 33924 16264 33930
rect 16212 33866 16264 33872
rect 16028 33856 16080 33862
rect 16028 33798 16080 33804
rect 16224 33658 16252 33866
rect 15844 33652 15896 33658
rect 15844 33594 15896 33600
rect 16212 33652 16264 33658
rect 16212 33594 16264 33600
rect 15752 30864 15804 30870
rect 15752 30806 15804 30812
rect 15016 30116 15068 30122
rect 15016 30058 15068 30064
rect 14188 29504 14240 29510
rect 14188 29446 14240 29452
rect 14200 29238 14228 29446
rect 14188 29232 14240 29238
rect 14188 29174 14240 29180
rect 14372 28960 14424 28966
rect 14372 28902 14424 28908
rect 14004 28756 14056 28762
rect 14004 28698 14056 28704
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 13820 28552 13872 28558
rect 13820 28494 13872 28500
rect 13636 28416 13688 28422
rect 13636 28358 13688 28364
rect 13648 28150 13676 28358
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 13728 27056 13780 27062
rect 13556 27024 13728 27044
rect 13780 27024 13782 27033
rect 13556 27016 13726 27024
rect 13084 26988 13136 26994
rect 13726 26959 13782 26968
rect 13084 26930 13136 26936
rect 13096 26586 13124 26930
rect 12992 26580 13044 26586
rect 12992 26522 13044 26528
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 12624 25832 12676 25838
rect 12544 25792 12624 25820
rect 12900 25832 12952 25838
rect 12676 25792 12756 25820
rect 12624 25774 12676 25780
rect 12440 22704 12492 22710
rect 12492 22652 12664 22658
rect 12440 22646 12664 22652
rect 12452 22630 12664 22646
rect 12636 22574 12664 22630
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 12728 22386 12756 25792
rect 12900 25774 12952 25780
rect 12808 22704 12860 22710
rect 12912 22658 12940 25774
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 13280 24138 13308 24686
rect 13268 24132 13320 24138
rect 13268 24074 13320 24080
rect 13280 23662 13308 24074
rect 13268 23656 13320 23662
rect 13268 23598 13320 23604
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 12860 22652 12940 22658
rect 12808 22646 12940 22652
rect 12820 22630 12940 22646
rect 12268 22066 12388 22094
rect 12544 22358 12756 22386
rect 12268 19990 12296 22066
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12360 21350 12388 21966
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 12544 20534 12572 22358
rect 12912 22216 12940 22630
rect 12636 22188 12940 22216
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12256 19984 12308 19990
rect 12256 19926 12308 19932
rect 12268 19786 12296 19926
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14890 11928 14962
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11900 14498 11928 14826
rect 11808 14470 11928 14498
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11532 12406 11652 12434
rect 11532 10724 11560 12406
rect 11716 11082 11744 14350
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11808 10962 11836 14470
rect 11992 14278 12020 14894
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11900 13870 11928 14214
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 12176 13802 12204 19246
rect 12360 16658 12388 20402
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12544 16726 12572 18906
rect 12636 18442 12664 22188
rect 12716 21956 12768 21962
rect 12716 21898 12768 21904
rect 12728 21622 12756 21898
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 13280 20466 13308 23598
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 13176 19780 13228 19786
rect 13176 19722 13228 19728
rect 12636 18414 12848 18442
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12636 16726 12664 18226
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12636 16182 12664 16662
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12256 15632 12308 15638
rect 12256 15574 12308 15580
rect 12268 15026 12296 15574
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12360 14414 12388 15370
rect 12728 15162 12756 17546
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12164 13320 12216 13326
rect 12216 13280 12296 13308
rect 12164 13262 12216 13268
rect 12268 12646 12296 13280
rect 12360 13190 12388 13466
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12544 12782 12572 14418
rect 12820 13870 12848 18414
rect 13188 17134 13216 19722
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13188 15638 13216 16050
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 13188 15502 13216 15574
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13280 14550 13308 20266
rect 13556 18970 13584 23598
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13740 22982 13768 23462
rect 13832 23050 13860 28494
rect 14016 28422 14044 28698
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 13924 23526 13952 23802
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13832 22166 13860 22986
rect 14200 22710 14228 24686
rect 14292 24274 14320 25230
rect 14280 24268 14332 24274
rect 14280 24210 14332 24216
rect 14292 23118 14320 24210
rect 14384 23866 14412 28902
rect 14556 28688 14608 28694
rect 14556 28630 14608 28636
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 14372 23860 14424 23866
rect 14372 23802 14424 23808
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14188 22704 14240 22710
rect 14188 22646 14240 22652
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 14200 22094 14228 22646
rect 14016 22066 14228 22094
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13728 20528 13780 20534
rect 13728 20470 13780 20476
rect 13740 20398 13768 20470
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13636 19440 13688 19446
rect 13636 19382 13688 19388
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13556 18086 13584 18566
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13648 16590 13676 19382
rect 13740 19378 13768 19654
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13832 19174 13860 20742
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13740 16250 13768 18362
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13832 17542 13860 18158
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 14016 15026 14044 22066
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14108 19378 14136 21490
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14108 18834 14136 19314
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 14108 18358 14136 18770
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 14200 17338 14228 20470
rect 14372 19168 14424 19174
rect 14292 19116 14372 19122
rect 14292 19110 14424 19116
rect 14292 19094 14412 19110
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13280 13938 13308 14486
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12728 13326 12756 13466
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12176 11694 12204 12310
rect 12268 11694 12296 12582
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11716 10934 11836 10962
rect 11532 10696 11652 10724
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11624 9178 11652 10696
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 7116 800 7144 2382
rect 8404 800 8432 2382
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9048 2106 9076 2246
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 9692 800 9720 2382
rect 11348 2378 11376 8910
rect 11716 5234 11744 10934
rect 11900 10742 11928 11562
rect 12544 11354 12572 12106
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11808 9994 11836 10542
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11808 9382 11836 9930
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11336 2372 11388 2378
rect 11336 2314 11388 2320
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 800 11008 2246
rect 11624 800 11652 2926
rect 11716 2446 11744 4966
rect 11992 3058 12020 11290
rect 12728 11082 12756 12582
rect 13280 12170 13308 13194
rect 13372 12918 13400 13670
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13556 12986 13584 13262
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13740 12850 13768 13806
rect 13832 13530 13860 13942
rect 14016 13938 14044 14962
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 14292 12238 14320 19094
rect 14476 12434 14504 28494
rect 14568 28082 14596 28630
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 15016 28144 15068 28150
rect 15016 28086 15068 28092
rect 14556 28076 14608 28082
rect 14556 28018 14608 28024
rect 14568 27878 14596 28018
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 15028 24750 15056 28086
rect 15212 28014 15240 28494
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 15764 28121 15792 28426
rect 15856 28393 15884 33594
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15948 32570 15976 32778
rect 15936 32564 15988 32570
rect 15936 32506 15988 32512
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 15948 31754 15976 31962
rect 15936 31748 15988 31754
rect 15936 31690 15988 31696
rect 16212 30728 16264 30734
rect 16212 30670 16264 30676
rect 16224 30394 16252 30670
rect 16212 30388 16264 30394
rect 16212 30330 16264 30336
rect 16316 29889 16344 34410
rect 16408 30394 16436 35158
rect 16488 35148 16540 35154
rect 16488 35090 16540 35096
rect 16500 34474 16528 35090
rect 16488 34468 16540 34474
rect 16488 34410 16540 34416
rect 16592 32842 16620 35255
rect 16684 34746 16712 36586
rect 16776 36174 16804 36654
rect 17406 36615 17462 36624
rect 16948 36576 17000 36582
rect 16948 36518 17000 36524
rect 17132 36576 17184 36582
rect 17132 36518 17184 36524
rect 16960 36417 16988 36518
rect 16946 36408 17002 36417
rect 16946 36343 17002 36352
rect 16764 36168 16816 36174
rect 16764 36110 16816 36116
rect 16776 35680 16804 36110
rect 16948 35828 17000 35834
rect 16948 35770 17000 35776
rect 16776 35652 16896 35680
rect 16868 35086 16896 35652
rect 16960 35465 16988 35770
rect 16946 35456 17002 35465
rect 16946 35391 17002 35400
rect 17144 35154 17172 36518
rect 17224 35624 17276 35630
rect 17224 35566 17276 35572
rect 17132 35148 17184 35154
rect 17132 35090 17184 35096
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 16672 34740 16724 34746
rect 16672 34682 16724 34688
rect 16684 34406 16712 34682
rect 16868 34542 16896 35022
rect 16948 34944 17000 34950
rect 16946 34912 16948 34921
rect 17000 34912 17002 34921
rect 16946 34847 17002 34856
rect 17236 34542 17264 35566
rect 17500 35148 17552 35154
rect 17500 35090 17552 35096
rect 17408 34672 17460 34678
rect 17512 34660 17540 35090
rect 17460 34632 17540 34660
rect 17408 34614 17460 34620
rect 16856 34536 16908 34542
rect 16856 34478 16908 34484
rect 17224 34536 17276 34542
rect 17224 34478 17276 34484
rect 16672 34400 16724 34406
rect 16672 34342 16724 34348
rect 16868 34066 16896 34478
rect 16948 34400 17000 34406
rect 16948 34342 17000 34348
rect 16960 34066 16988 34342
rect 16856 34060 16908 34066
rect 16856 34002 16908 34008
rect 16948 34060 17000 34066
rect 16948 34002 17000 34008
rect 17408 34060 17460 34066
rect 17408 34002 17460 34008
rect 16868 33454 16896 34002
rect 17420 33658 17448 34002
rect 17684 33856 17736 33862
rect 17684 33798 17736 33804
rect 17408 33652 17460 33658
rect 17408 33594 17460 33600
rect 17500 33652 17552 33658
rect 17500 33594 17552 33600
rect 17132 33584 17184 33590
rect 17184 33544 17356 33572
rect 17132 33526 17184 33532
rect 17328 33538 17356 33544
rect 17512 33538 17540 33594
rect 17328 33510 17540 33538
rect 16856 33448 16908 33454
rect 16856 33390 16908 33396
rect 16764 32972 16816 32978
rect 16764 32914 16816 32920
rect 16580 32836 16632 32842
rect 16580 32778 16632 32784
rect 16776 32756 16804 32914
rect 16868 32910 16896 33390
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 17040 32836 17092 32842
rect 17040 32778 17092 32784
rect 16776 32728 16896 32756
rect 16764 32428 16816 32434
rect 16764 32370 16816 32376
rect 16776 31890 16804 32370
rect 16764 31884 16816 31890
rect 16764 31826 16816 31832
rect 16868 31754 16896 32728
rect 17052 31754 17080 32778
rect 16592 31726 16896 31754
rect 16948 31748 17000 31754
rect 16396 30388 16448 30394
rect 16396 30330 16448 30336
rect 16302 29880 16358 29889
rect 16302 29815 16358 29824
rect 16120 29096 16172 29102
rect 16120 29038 16172 29044
rect 16132 28966 16160 29038
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 16120 28960 16172 28966
rect 16120 28902 16172 28908
rect 15948 28762 15976 28902
rect 15936 28756 15988 28762
rect 15936 28698 15988 28704
rect 15842 28384 15898 28393
rect 15842 28319 15898 28328
rect 15750 28112 15806 28121
rect 15750 28047 15806 28056
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 15212 27538 15240 27950
rect 15200 27532 15252 27538
rect 15200 27474 15252 27480
rect 15382 26752 15438 26761
rect 15382 26687 15438 26696
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 15212 24070 15240 24754
rect 15200 24064 15252 24070
rect 15200 24006 15252 24012
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 14568 22710 14596 22986
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14752 22234 14780 22918
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 14936 20806 14964 21082
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14844 16726 14872 17478
rect 14832 16720 14884 16726
rect 14832 16662 14884 16668
rect 14646 13424 14702 13433
rect 14646 13359 14702 13368
rect 14660 13326 14688 13359
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14660 12646 14688 13262
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14384 12406 14504 12434
rect 14280 12232 14332 12238
rect 13358 12200 13414 12209
rect 13268 12164 13320 12170
rect 14280 12174 14332 12180
rect 13358 12135 13414 12144
rect 13268 12106 13320 12112
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12084 9178 12112 9454
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12176 4486 12204 11018
rect 12636 10266 12664 11018
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12452 7886 12480 8298
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12912 7274 12940 10610
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12912 800 12940 2382
rect 13004 2106 13032 9998
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13188 3126 13216 8910
rect 13280 8430 13308 12106
rect 13372 12102 13400 12135
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13464 10810 13492 11766
rect 14292 11694 14320 12174
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14384 11506 14412 12406
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11762 14688 12038
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14292 11478 14412 11506
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 14096 10736 14148 10742
rect 14292 10724 14320 11478
rect 14752 11286 14780 13194
rect 14936 12238 14964 20742
rect 15028 18970 15056 23802
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 15120 21554 15148 21966
rect 15212 21622 15240 24006
rect 15396 21962 15424 26687
rect 15764 26518 15792 28047
rect 15752 26512 15804 26518
rect 15752 26454 15804 26460
rect 15856 22094 15884 28319
rect 16132 27520 16160 28902
rect 16592 28558 16620 31726
rect 17052 31748 17184 31754
rect 17052 31726 17132 31748
rect 16948 31690 17000 31696
rect 17132 31690 17184 31696
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16672 31272 16724 31278
rect 16672 31214 16724 31220
rect 16684 30326 16712 31214
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16762 30288 16818 30297
rect 16868 30258 16896 31282
rect 16960 30308 16988 31690
rect 17408 31408 17460 31414
rect 17460 31368 17632 31396
rect 17408 31350 17460 31356
rect 17604 31142 17632 31368
rect 17696 31249 17724 33798
rect 17788 31754 17816 37198
rect 17880 36582 17908 37198
rect 18616 37194 18736 37210
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 18604 37188 18736 37194
rect 18656 37182 18736 37188
rect 18604 37130 18656 37136
rect 18788 37120 18840 37126
rect 18788 37062 18840 37068
rect 18420 36848 18472 36854
rect 18420 36790 18472 36796
rect 18236 36780 18288 36786
rect 18236 36722 18288 36728
rect 18144 36644 18196 36650
rect 18144 36586 18196 36592
rect 17868 36576 17920 36582
rect 17868 36518 17920 36524
rect 18156 36174 18184 36586
rect 18248 36310 18276 36722
rect 18326 36408 18382 36417
rect 18432 36378 18460 36790
rect 18800 36378 18828 37062
rect 19444 36802 19472 37198
rect 19996 37126 20024 39200
rect 21284 37330 21312 39200
rect 21272 37324 21324 37330
rect 21272 37266 21324 37272
rect 20996 37256 21048 37262
rect 20732 37194 20944 37210
rect 20996 37198 21048 37204
rect 20720 37188 20956 37194
rect 20772 37182 20904 37188
rect 20720 37130 20772 37136
rect 20904 37130 20956 37136
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20534 36952 20590 36961
rect 20076 36916 20128 36922
rect 21008 36922 21036 37198
rect 21928 37194 21956 39200
rect 23216 37330 23244 39200
rect 23204 37324 23256 37330
rect 23204 37266 23256 37272
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 23112 37256 23164 37262
rect 23388 37256 23440 37262
rect 23112 37198 23164 37204
rect 23216 37204 23388 37210
rect 23216 37198 23440 37204
rect 21916 37188 21968 37194
rect 21916 37130 21968 37136
rect 20534 36887 20590 36896
rect 20628 36916 20680 36922
rect 20076 36858 20128 36864
rect 19340 36780 19392 36786
rect 19444 36774 19748 36802
rect 20088 36786 20116 36858
rect 19340 36722 19392 36728
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 19260 36417 19288 36654
rect 19246 36408 19302 36417
rect 18326 36343 18382 36352
rect 18420 36372 18472 36378
rect 18236 36304 18288 36310
rect 18236 36246 18288 36252
rect 18340 36174 18368 36343
rect 18420 36314 18472 36320
rect 18788 36372 18840 36378
rect 19246 36343 19302 36352
rect 18788 36314 18840 36320
rect 18144 36168 18196 36174
rect 18144 36110 18196 36116
rect 18328 36168 18380 36174
rect 18328 36110 18380 36116
rect 18512 36032 18564 36038
rect 18696 36032 18748 36038
rect 18512 35974 18564 35980
rect 18694 36000 18696 36009
rect 18748 36000 18750 36009
rect 18524 35737 18552 35974
rect 18694 35935 18750 35944
rect 18510 35728 18566 35737
rect 18510 35663 18566 35672
rect 17868 35624 17920 35630
rect 17868 35566 17920 35572
rect 17880 34746 17908 35566
rect 18420 35556 18472 35562
rect 18420 35498 18472 35504
rect 17958 34912 18014 34921
rect 17958 34847 18014 34856
rect 17972 34746 18000 34847
rect 17868 34740 17920 34746
rect 17868 34682 17920 34688
rect 17960 34740 18012 34746
rect 17960 34682 18012 34688
rect 18144 34468 18196 34474
rect 18144 34410 18196 34416
rect 18156 34377 18184 34410
rect 18142 34368 18198 34377
rect 18142 34303 18198 34312
rect 18432 34066 18460 35498
rect 18524 35494 18552 35663
rect 18512 35488 18564 35494
rect 18512 35430 18564 35436
rect 19352 35222 19380 36722
rect 19720 36174 19748 36774
rect 20076 36780 20128 36786
rect 20076 36722 20128 36728
rect 20548 36718 20576 36887
rect 20628 36858 20680 36864
rect 20996 36916 21048 36922
rect 20996 36858 21048 36864
rect 21916 36916 21968 36922
rect 21916 36858 21968 36864
rect 20536 36712 20588 36718
rect 20536 36654 20588 36660
rect 20260 36576 20312 36582
rect 20260 36518 20312 36524
rect 20272 36242 20300 36518
rect 20536 36372 20588 36378
rect 20536 36314 20588 36320
rect 20260 36236 20312 36242
rect 20260 36178 20312 36184
rect 19708 36168 19760 36174
rect 19708 36110 19760 36116
rect 20076 36168 20128 36174
rect 20076 36110 20128 36116
rect 19432 36100 19484 36106
rect 19432 36042 19484 36048
rect 19340 35216 19392 35222
rect 19340 35158 19392 35164
rect 19444 35086 19472 36042
rect 19708 36032 19760 36038
rect 19760 35992 20024 36020
rect 19708 35974 19760 35980
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35698 20024 35992
rect 20088 35873 20116 36110
rect 20548 36106 20576 36314
rect 20168 36100 20220 36106
rect 20168 36042 20220 36048
rect 20536 36100 20588 36106
rect 20536 36042 20588 36048
rect 20074 35864 20130 35873
rect 20074 35799 20130 35808
rect 19984 35692 20036 35698
rect 19984 35634 20036 35640
rect 20180 35630 20208 36042
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 20168 35624 20220 35630
rect 20168 35566 20220 35572
rect 19984 35216 20036 35222
rect 19984 35158 20036 35164
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 18604 34944 18656 34950
rect 18604 34886 18656 34892
rect 18512 34400 18564 34406
rect 18616 34388 18644 34886
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19996 34746 20024 35158
rect 20180 35086 20208 35566
rect 20168 35080 20220 35086
rect 20168 35022 20220 35028
rect 20260 35080 20312 35086
rect 20260 35022 20312 35028
rect 20168 34944 20220 34950
rect 20168 34886 20220 34892
rect 19984 34740 20036 34746
rect 19984 34682 20036 34688
rect 18564 34360 18644 34388
rect 18512 34342 18564 34348
rect 18616 34134 18644 34360
rect 18512 34128 18564 34134
rect 18512 34070 18564 34076
rect 18604 34128 18656 34134
rect 18604 34070 18656 34076
rect 18420 34060 18472 34066
rect 18420 34002 18472 34008
rect 17868 33856 17920 33862
rect 17868 33798 17920 33804
rect 17880 33454 17908 33798
rect 17868 33448 17920 33454
rect 17868 33390 17920 33396
rect 18524 33318 18552 34070
rect 19156 33992 19208 33998
rect 19156 33934 19208 33940
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 19168 33114 19196 33934
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19246 33144 19302 33153
rect 18972 33108 19024 33114
rect 18972 33050 19024 33056
rect 19156 33108 19208 33114
rect 19246 33079 19302 33088
rect 19156 33050 19208 33056
rect 18880 33040 18932 33046
rect 18708 32988 18880 32994
rect 18708 32982 18932 32988
rect 18708 32966 18920 32982
rect 18708 32910 18736 32966
rect 18696 32904 18748 32910
rect 18696 32846 18748 32852
rect 18880 32904 18932 32910
rect 18880 32846 18932 32852
rect 18892 32570 18920 32846
rect 18984 32570 19012 33050
rect 18880 32564 18932 32570
rect 18880 32506 18932 32512
rect 18972 32564 19024 32570
rect 18972 32506 19024 32512
rect 19260 32502 19288 33079
rect 19432 33040 19484 33046
rect 19484 33000 19564 33028
rect 19432 32982 19484 32988
rect 19536 32960 19564 33000
rect 19616 32972 19668 32978
rect 19536 32932 19616 32960
rect 19616 32914 19668 32920
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19248 32496 19300 32502
rect 19248 32438 19300 32444
rect 18512 32428 18564 32434
rect 18512 32370 18564 32376
rect 18524 31890 18552 32370
rect 18972 32360 19024 32366
rect 18972 32302 19024 32308
rect 18696 32292 18748 32298
rect 18696 32234 18748 32240
rect 18512 31884 18564 31890
rect 18432 31844 18512 31872
rect 17788 31726 17908 31754
rect 17682 31240 17738 31249
rect 17682 31175 17738 31184
rect 17500 31136 17552 31142
rect 17500 31078 17552 31084
rect 17592 31136 17644 31142
rect 17592 31078 17644 31084
rect 17316 30320 17368 30326
rect 16960 30280 17172 30308
rect 16762 30223 16764 30232
rect 16816 30223 16818 30232
rect 16856 30252 16908 30258
rect 16764 30194 16816 30200
rect 16856 30194 16908 30200
rect 16868 29730 16896 30194
rect 16946 30152 17002 30161
rect 16946 30087 16948 30096
rect 17000 30087 17002 30096
rect 16948 30058 17000 30064
rect 16776 29714 16896 29730
rect 16764 29708 16896 29714
rect 16816 29702 16896 29708
rect 17040 29708 17092 29714
rect 16764 29650 16816 29656
rect 17040 29650 17092 29656
rect 16672 29572 16724 29578
rect 16672 29514 16724 29520
rect 16684 29034 16712 29514
rect 16776 29306 16804 29650
rect 16764 29300 16816 29306
rect 16764 29242 16816 29248
rect 17052 29186 17080 29650
rect 16776 29158 17080 29186
rect 16672 29028 16724 29034
rect 16672 28970 16724 28976
rect 16776 28642 16804 29158
rect 16856 29096 16908 29102
rect 16856 29038 16908 29044
rect 16684 28614 16804 28642
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16304 27940 16356 27946
rect 16304 27882 16356 27888
rect 16212 27532 16264 27538
rect 16132 27492 16212 27520
rect 16212 27474 16264 27480
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 16040 25430 16068 25774
rect 16028 25424 16080 25430
rect 16028 25366 16080 25372
rect 16316 24954 16344 27882
rect 16486 27568 16542 27577
rect 16486 27503 16488 27512
rect 16540 27503 16542 27512
rect 16488 27474 16540 27480
rect 16396 27396 16448 27402
rect 16684 27384 16712 28614
rect 16868 28558 16896 29038
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16764 28484 16816 28490
rect 16764 28426 16816 28432
rect 16776 28082 16804 28426
rect 16764 28076 16816 28082
rect 16764 28018 16816 28024
rect 16868 28014 16896 28494
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16856 28008 16908 28014
rect 16856 27950 16908 27956
rect 16448 27356 16712 27384
rect 16396 27338 16448 27344
rect 16868 26994 16896 27950
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16868 26450 16896 26930
rect 16856 26444 16908 26450
rect 16960 26432 16988 28358
rect 17144 27606 17172 30280
rect 17316 30262 17368 30268
rect 17224 29232 17276 29238
rect 17224 29174 17276 29180
rect 17236 28694 17264 29174
rect 17224 28688 17276 28694
rect 17224 28630 17276 28636
rect 17236 28150 17264 28630
rect 17224 28144 17276 28150
rect 17224 28086 17276 28092
rect 17132 27600 17184 27606
rect 17132 27542 17184 27548
rect 17144 27062 17172 27542
rect 17132 27056 17184 27062
rect 17132 26998 17184 27004
rect 16960 26404 17080 26432
rect 16856 26386 16908 26392
rect 16946 26344 17002 26353
rect 16580 26308 16632 26314
rect 16946 26279 16948 26288
rect 16580 26250 16632 26256
rect 17000 26279 17002 26288
rect 16948 26250 17000 26256
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16500 24886 16528 25094
rect 16488 24880 16540 24886
rect 16488 24822 16540 24828
rect 16500 23186 16528 24822
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 16592 22982 16620 26250
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16868 24732 16896 25774
rect 16948 24744 17000 24750
rect 16868 24704 16948 24732
rect 16868 24274 16896 24704
rect 16948 24686 17000 24692
rect 17052 24562 17080 26404
rect 16960 24534 17080 24562
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16776 23866 16804 24074
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16868 23730 16896 24210
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16868 23186 16896 23462
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 15856 22066 15976 22094
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15200 21616 15252 21622
rect 15200 21558 15252 21564
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 15120 21010 15148 21490
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15120 19922 15148 20470
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 15028 17882 15056 18634
rect 15016 17876 15068 17882
rect 15016 17818 15068 17824
rect 15028 17066 15056 17818
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 15120 16590 15148 18634
rect 15304 18426 15332 19994
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15212 16998 15240 17478
rect 15304 17134 15332 18362
rect 15948 17202 15976 22066
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16224 20806 16252 20946
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16408 18766 16436 21082
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16500 19786 16528 20402
rect 16592 19922 16620 21490
rect 16684 20318 16896 20346
rect 16684 20262 16712 20318
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16500 17202 16528 19722
rect 16592 19378 16620 19858
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16592 18290 16620 19314
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16592 17746 16620 18226
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16684 17610 16712 19450
rect 16776 19446 16804 20198
rect 16868 19768 16896 20318
rect 16960 19922 16988 24534
rect 17144 22094 17172 26998
rect 17328 26450 17356 30262
rect 17512 28490 17540 31078
rect 17604 30938 17632 31078
rect 17592 30932 17644 30938
rect 17592 30874 17644 30880
rect 17500 28484 17552 28490
rect 17500 28426 17552 28432
rect 17408 27396 17460 27402
rect 17408 27338 17460 27344
rect 17316 26444 17368 26450
rect 17316 26386 17368 26392
rect 17420 26353 17448 27338
rect 17406 26344 17462 26353
rect 17406 26279 17462 26288
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17236 25974 17264 26182
rect 17224 25968 17276 25974
rect 17224 25910 17276 25916
rect 17512 24818 17540 28426
rect 17696 28014 17724 31175
rect 17776 30864 17828 30870
rect 17776 30806 17828 30812
rect 17788 30598 17816 30806
rect 17776 30592 17828 30598
rect 17776 30534 17828 30540
rect 17774 29880 17830 29889
rect 17774 29815 17776 29824
rect 17828 29815 17830 29824
rect 17776 29786 17828 29792
rect 17880 29730 17908 31726
rect 18432 30802 18460 31844
rect 18512 31826 18564 31832
rect 18708 31754 18736 32234
rect 18984 32230 19012 32302
rect 18972 32224 19024 32230
rect 18972 32166 19024 32172
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 18788 31816 18840 31822
rect 18788 31758 18840 31764
rect 18524 31726 18736 31754
rect 18420 30796 18472 30802
rect 18420 30738 18472 30744
rect 18236 30592 18288 30598
rect 18236 30534 18288 30540
rect 17960 30184 18012 30190
rect 18012 30144 18184 30172
rect 17960 30126 18012 30132
rect 18156 29753 18184 30144
rect 17788 29702 17908 29730
rect 18142 29744 18198 29753
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17788 27441 17816 29702
rect 18142 29679 18198 29688
rect 18156 29102 18184 29679
rect 18248 29646 18276 30534
rect 18326 30152 18382 30161
rect 18326 30087 18328 30096
rect 18380 30087 18382 30096
rect 18328 30058 18380 30064
rect 18420 29844 18472 29850
rect 18420 29786 18472 29792
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 18432 29578 18460 29786
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 17868 29096 17920 29102
rect 18144 29096 18196 29102
rect 17920 29044 18000 29050
rect 17868 29038 18000 29044
rect 18144 29038 18196 29044
rect 17880 29022 18000 29038
rect 17972 28506 18000 29022
rect 17972 28478 18368 28506
rect 17868 28416 17920 28422
rect 17866 28384 17868 28393
rect 17920 28384 17922 28393
rect 17866 28319 17922 28328
rect 17866 28112 17922 28121
rect 17866 28047 17922 28056
rect 17880 28014 17908 28047
rect 17868 28008 17920 28014
rect 17868 27950 17920 27956
rect 18236 27940 18288 27946
rect 18236 27882 18288 27888
rect 17868 27872 17920 27878
rect 18144 27872 18196 27878
rect 17920 27820 18092 27826
rect 17868 27814 18092 27820
rect 18144 27814 18196 27820
rect 17880 27798 18092 27814
rect 17958 27704 18014 27713
rect 18064 27674 18092 27798
rect 17958 27639 17960 27648
rect 18012 27639 18014 27648
rect 18052 27668 18104 27674
rect 17960 27610 18012 27616
rect 18052 27610 18104 27616
rect 17774 27432 17830 27441
rect 17774 27367 17830 27376
rect 18064 25294 18092 27610
rect 18156 25838 18184 27814
rect 18248 27470 18276 27882
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18052 25288 18104 25294
rect 18052 25230 18104 25236
rect 18156 24954 18184 25774
rect 18340 25770 18368 28478
rect 18524 27554 18552 31726
rect 18604 31136 18656 31142
rect 18604 31078 18656 31084
rect 18616 28762 18644 31078
rect 18696 30048 18748 30054
rect 18696 29990 18748 29996
rect 18604 28756 18656 28762
rect 18604 28698 18656 28704
rect 18708 27674 18736 29990
rect 18800 29646 18828 31758
rect 19248 30728 19300 30734
rect 19248 30670 19300 30676
rect 19260 30546 19288 30670
rect 19352 30666 19380 32166
rect 19444 31113 19472 32846
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19984 32496 20036 32502
rect 19984 32438 20036 32444
rect 19996 31754 20024 32438
rect 19996 31726 20116 31754
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19430 31104 19486 31113
rect 19430 31039 19486 31048
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 19340 30660 19392 30666
rect 19340 30602 19392 30608
rect 19260 30518 19380 30546
rect 18880 30388 18932 30394
rect 18880 30330 18932 30336
rect 18892 29850 18920 30330
rect 19352 30258 19380 30518
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19708 30252 19760 30258
rect 19708 30194 19760 30200
rect 19720 30161 19748 30194
rect 19706 30152 19762 30161
rect 19706 30087 19762 30096
rect 19064 30048 19116 30054
rect 19064 29990 19116 29996
rect 18880 29844 18932 29850
rect 18880 29786 18932 29792
rect 18788 29640 18840 29646
rect 18788 29582 18840 29588
rect 19076 29306 19104 29990
rect 19338 29608 19394 29617
rect 19338 29543 19394 29552
rect 19432 29572 19484 29578
rect 19064 29300 19116 29306
rect 19064 29242 19116 29248
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 19168 28082 19196 29242
rect 19352 28694 19380 29543
rect 19432 29514 19484 29520
rect 19444 29209 19472 29514
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19430 29200 19486 29209
rect 19430 29135 19486 29144
rect 19340 28688 19392 28694
rect 19340 28630 19392 28636
rect 19432 28688 19484 28694
rect 19432 28630 19484 28636
rect 19444 28422 19472 28630
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19064 28076 19116 28082
rect 19064 28018 19116 28024
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 18786 27704 18842 27713
rect 18696 27668 18748 27674
rect 18786 27639 18788 27648
rect 18696 27610 18748 27616
rect 18840 27639 18842 27648
rect 18788 27610 18840 27616
rect 18524 27526 18920 27554
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 18512 26988 18564 26994
rect 18512 26930 18564 26936
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18432 25838 18460 25978
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 18328 25764 18380 25770
rect 18328 25706 18380 25712
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18326 25664 18382 25673
rect 18248 25294 18276 25638
rect 18326 25599 18382 25608
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18052 24948 18104 24954
rect 18052 24890 18104 24896
rect 18144 24948 18196 24954
rect 18144 24890 18196 24896
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17684 24744 17736 24750
rect 17604 24704 17684 24732
rect 17604 24698 17632 24704
rect 17512 24670 17632 24698
rect 17684 24686 17736 24692
rect 17512 24614 17540 24670
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 18064 24018 18092 24890
rect 18340 24818 18368 25599
rect 18524 25378 18552 26930
rect 18616 25702 18644 27406
rect 18788 26784 18840 26790
rect 18786 26752 18788 26761
rect 18840 26752 18842 26761
rect 18786 26687 18842 26696
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18800 26217 18828 26318
rect 18786 26208 18842 26217
rect 18786 26143 18842 26152
rect 18788 25900 18840 25906
rect 18788 25842 18840 25848
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 18696 25696 18748 25702
rect 18696 25638 18748 25644
rect 18616 25498 18644 25638
rect 18604 25492 18656 25498
rect 18604 25434 18656 25440
rect 18524 25350 18644 25378
rect 18328 24812 18380 24818
rect 18248 24772 18328 24800
rect 18144 24064 18196 24070
rect 18064 24012 18144 24018
rect 18064 24006 18196 24012
rect 18064 23990 18184 24006
rect 17224 23248 17276 23254
rect 17224 23190 17276 23196
rect 17236 22778 17264 23190
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17052 22066 17172 22094
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16948 19780 17000 19786
rect 16868 19740 16948 19768
rect 16948 19722 17000 19728
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15304 16590 15332 17070
rect 16960 16658 16988 19722
rect 17052 17882 17080 22066
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17144 19310 17172 19654
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17236 18358 17264 21014
rect 17224 18352 17276 18358
rect 17224 18294 17276 18300
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16316 16114 16344 16390
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15016 14884 15068 14890
rect 15016 14826 15068 14832
rect 15028 14414 15056 14826
rect 15016 14408 15068 14414
rect 15068 14368 15148 14396
rect 15016 14350 15068 14356
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15028 12170 15056 13806
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14148 10696 14320 10724
rect 14096 10678 14148 10684
rect 14384 10674 14412 10950
rect 14844 10674 14872 10950
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14936 10606 14964 10950
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 14568 5846 14596 10542
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 9722 14780 10406
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14844 8090 14872 9930
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14556 5840 14608 5846
rect 14556 5782 14608 5788
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13188 2514 13216 3062
rect 14752 2650 14780 7822
rect 15120 6914 15148 14368
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15304 13870 15332 14282
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15672 13734 15700 15370
rect 16592 15162 16620 15642
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16224 14074 16252 15030
rect 16592 14958 16620 15098
rect 16776 15094 16804 16390
rect 16868 15434 16896 16458
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16764 15088 16816 15094
rect 16670 15056 16726 15065
rect 16764 15030 16816 15036
rect 16670 14991 16672 15000
rect 16724 14991 16726 15000
rect 16672 14962 16724 14968
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16868 14618 16896 15370
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15658 13560 15714 13569
rect 15658 13495 15714 13504
rect 15672 13326 15700 13495
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11150 15240 11494
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 8498 15240 10406
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15028 6886 15148 6914
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 12992 2100 13044 2106
rect 12992 2042 13044 2048
rect 14200 800 14228 2382
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 800 14872 2246
rect 15028 2038 15056 6886
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15212 5778 15240 6190
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15304 5642 15332 12038
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 10470 15424 11630
rect 15580 11082 15608 12718
rect 15948 12306 15976 13330
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15672 11082 15700 11222
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16224 10538 16252 11018
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 16500 9926 16528 13806
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16684 12442 16712 13330
rect 16960 12986 16988 16594
rect 17052 16182 17080 16934
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 17052 13326 17080 13398
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17144 12442 17172 13942
rect 17236 13530 17264 14894
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17328 13410 17356 21830
rect 17236 13382 17356 13410
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17144 12306 17172 12378
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17236 12238 17264 13382
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17328 12850 17356 13194
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17420 12434 17448 22918
rect 18248 22710 18276 24772
rect 18328 24754 18380 24760
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 18432 23798 18460 24550
rect 18616 24426 18644 25350
rect 18524 24398 18644 24426
rect 18420 23792 18472 23798
rect 18420 23734 18472 23740
rect 18524 23118 18552 24398
rect 18708 24342 18736 25638
rect 18696 24336 18748 24342
rect 18696 24278 18748 24284
rect 18696 24200 18748 24206
rect 18800 24188 18828 25842
rect 18748 24160 18828 24188
rect 18696 24142 18748 24148
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18236 22704 18288 22710
rect 18236 22646 18288 22652
rect 17592 22432 17644 22438
rect 17592 22374 17644 22380
rect 17604 21962 17632 22374
rect 17592 21956 17644 21962
rect 17592 21898 17644 21904
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17788 21146 17816 21626
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17604 16794 17632 17750
rect 17788 17338 17816 19382
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 17512 16250 17540 16458
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17880 15586 17908 21830
rect 18248 19334 18276 22646
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18524 21078 18552 21286
rect 18512 21072 18564 21078
rect 18512 21014 18564 21020
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18156 19306 18276 19334
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 18064 17202 18092 17614
rect 18156 17202 18184 19306
rect 18340 19174 18368 19654
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18432 17338 18460 18294
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 17788 15558 17908 15586
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17604 14482 17632 14894
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17696 14346 17724 14554
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17696 13274 17724 14282
rect 17328 12406 17448 12434
rect 17512 13246 17724 13274
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17328 11014 17356 12406
rect 17512 12374 17540 13246
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17604 12782 17632 13126
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17696 12714 17724 13126
rect 17788 12918 17816 15558
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17880 14482 17908 15370
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 13938 17908 14418
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 17972 13802 18000 15098
rect 18064 15065 18092 15438
rect 18050 15056 18106 15065
rect 18050 14991 18106 15000
rect 18340 14822 18368 15982
rect 18432 15201 18460 17138
rect 18418 15192 18474 15201
rect 18418 15127 18474 15136
rect 18432 15026 18460 15127
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18524 14906 18552 18566
rect 18616 18426 18644 23598
rect 18708 22642 18736 24142
rect 18892 24070 18920 27526
rect 18972 26988 19024 26994
rect 18972 26930 19024 26936
rect 18984 26858 19012 26930
rect 18972 26852 19024 26858
rect 18972 26794 19024 26800
rect 19076 25430 19104 28018
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19248 27600 19300 27606
rect 19248 27542 19300 27548
rect 19156 27056 19208 27062
rect 19156 26998 19208 27004
rect 19168 26042 19196 26998
rect 19260 26994 19288 27542
rect 19444 27470 19472 27814
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 19248 26512 19300 26518
rect 19248 26454 19300 26460
rect 19260 26314 19288 26454
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 19156 26036 19208 26042
rect 19156 25978 19208 25984
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19168 25673 19196 25842
rect 19154 25664 19210 25673
rect 19154 25599 19210 25608
rect 19064 25424 19116 25430
rect 19064 25366 19116 25372
rect 19156 25424 19208 25430
rect 19156 25366 19208 25372
rect 19168 24138 19196 25366
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 19260 24342 19288 25094
rect 19352 24750 19380 26998
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19248 24336 19300 24342
rect 19248 24278 19300 24284
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19156 24132 19208 24138
rect 19156 24074 19208 24080
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18800 22506 18828 24006
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18788 22500 18840 22506
rect 18788 22442 18840 22448
rect 18984 20534 19012 23054
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18708 16590 18736 19246
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18892 16046 18920 19314
rect 18984 18426 19012 20470
rect 19168 19334 19196 23462
rect 19260 23186 19288 24142
rect 19444 23662 19472 27406
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19892 26920 19944 26926
rect 19996 26908 20024 30670
rect 20088 28558 20116 31726
rect 20180 30802 20208 34886
rect 20272 33998 20300 35022
rect 20364 34921 20392 35634
rect 20536 35556 20588 35562
rect 20536 35498 20588 35504
rect 20444 34944 20496 34950
rect 20350 34912 20406 34921
rect 20444 34886 20496 34892
rect 20350 34847 20406 34856
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20272 32842 20300 33934
rect 20260 32836 20312 32842
rect 20260 32778 20312 32784
rect 20272 32434 20300 32778
rect 20260 32428 20312 32434
rect 20260 32370 20312 32376
rect 20168 30796 20220 30802
rect 20168 30738 20220 30744
rect 20272 30734 20300 32370
rect 20456 31754 20484 34886
rect 20548 34678 20576 35498
rect 20536 34672 20588 34678
rect 20536 34614 20588 34620
rect 20640 33046 20668 36858
rect 20720 36780 20772 36786
rect 20772 36740 20852 36768
rect 20720 36722 20772 36728
rect 20718 36680 20774 36689
rect 20718 36615 20774 36624
rect 20732 35834 20760 36615
rect 20824 36378 20852 36740
rect 21638 36680 21694 36689
rect 21638 36615 21694 36624
rect 21652 36378 21680 36615
rect 21928 36582 21956 36858
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22190 36680 22246 36689
rect 22100 36644 22152 36650
rect 22190 36615 22192 36624
rect 22100 36586 22152 36592
rect 22244 36615 22246 36624
rect 22192 36586 22244 36592
rect 21916 36576 21968 36582
rect 21916 36518 21968 36524
rect 22008 36576 22060 36582
rect 22008 36518 22060 36524
rect 20812 36372 20864 36378
rect 20812 36314 20864 36320
rect 21640 36372 21692 36378
rect 21640 36314 21692 36320
rect 21088 36236 21140 36242
rect 21088 36178 21140 36184
rect 20904 36100 20956 36106
rect 20904 36042 20956 36048
rect 20916 35834 20944 36042
rect 20720 35828 20772 35834
rect 20720 35770 20772 35776
rect 20904 35828 20956 35834
rect 20904 35770 20956 35776
rect 20720 35692 20772 35698
rect 20720 35634 20772 35640
rect 20732 35086 20760 35634
rect 20996 35488 21048 35494
rect 20810 35456 20866 35465
rect 20810 35391 20866 35400
rect 20994 35456 20996 35465
rect 21048 35456 21050 35465
rect 20994 35391 21050 35400
rect 20720 35080 20772 35086
rect 20720 35022 20772 35028
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20628 33040 20680 33046
rect 20628 32982 20680 32988
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20548 32434 20576 32846
rect 20536 32428 20588 32434
rect 20536 32370 20588 32376
rect 20628 31952 20680 31958
rect 20732 31906 20760 34886
rect 20824 34542 20852 35391
rect 20996 34944 21048 34950
rect 20916 34892 20996 34898
rect 20916 34886 21048 34892
rect 20916 34870 21036 34886
rect 20812 34536 20864 34542
rect 20812 34478 20864 34484
rect 20680 31900 20760 31906
rect 20628 31894 20760 31900
rect 20640 31878 20760 31894
rect 20824 31754 20852 34478
rect 20916 33658 20944 34870
rect 21100 33658 21128 36178
rect 21180 35828 21232 35834
rect 21180 35770 21232 35776
rect 21192 35494 21220 35770
rect 21548 35760 21600 35766
rect 21548 35702 21600 35708
rect 21272 35624 21324 35630
rect 21272 35566 21324 35572
rect 21180 35488 21232 35494
rect 21180 35430 21232 35436
rect 21192 34542 21220 35430
rect 21180 34536 21232 34542
rect 21180 34478 21232 34484
rect 21180 33856 21232 33862
rect 21180 33798 21232 33804
rect 21192 33658 21220 33798
rect 20904 33652 20956 33658
rect 20904 33594 20956 33600
rect 21088 33652 21140 33658
rect 21088 33594 21140 33600
rect 21180 33652 21232 33658
rect 21180 33594 21232 33600
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 21008 32745 21036 33458
rect 21100 32842 21128 33594
rect 21088 32836 21140 32842
rect 21088 32778 21140 32784
rect 21180 32836 21232 32842
rect 21180 32778 21232 32784
rect 20994 32736 21050 32745
rect 20994 32671 21050 32680
rect 21192 32609 21220 32778
rect 21178 32600 21234 32609
rect 21178 32535 21234 32544
rect 21088 32224 21140 32230
rect 21088 32166 21140 32172
rect 21100 32065 21128 32166
rect 21086 32056 21142 32065
rect 21086 31991 21142 32000
rect 20456 31726 20668 31754
rect 20824 31726 21036 31754
rect 20352 31340 20404 31346
rect 20352 31282 20404 31288
rect 20260 30728 20312 30734
rect 20260 30670 20312 30676
rect 20168 30592 20220 30598
rect 20168 30534 20220 30540
rect 20180 30326 20208 30534
rect 20168 30320 20220 30326
rect 20168 30262 20220 30268
rect 20364 29646 20392 31282
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 20168 29640 20220 29646
rect 20352 29640 20404 29646
rect 20220 29588 20300 29594
rect 20168 29582 20300 29588
rect 20352 29582 20404 29588
rect 20180 29566 20300 29582
rect 20076 28552 20128 28558
rect 20076 28494 20128 28500
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 20088 28150 20116 28358
rect 20076 28144 20128 28150
rect 20076 28086 20128 28092
rect 19944 26880 20024 26908
rect 19892 26862 19944 26868
rect 19984 26512 20036 26518
rect 19984 26454 20036 26460
rect 20074 26480 20130 26489
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19892 25424 19944 25430
rect 19890 25392 19892 25401
rect 19944 25392 19946 25401
rect 19890 25327 19946 25336
rect 19798 25256 19854 25265
rect 19996 25242 20024 26454
rect 20180 26450 20208 28358
rect 20272 27674 20300 29566
rect 20456 29102 20484 30738
rect 20536 30660 20588 30666
rect 20536 30602 20588 30608
rect 20548 30394 20576 30602
rect 20536 30388 20588 30394
rect 20536 30330 20588 30336
rect 20534 30288 20590 30297
rect 20534 30223 20590 30232
rect 20548 30122 20576 30223
rect 20536 30116 20588 30122
rect 20536 30058 20588 30064
rect 20640 30002 20668 31726
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 20824 30258 20852 31282
rect 20812 30252 20864 30258
rect 20812 30194 20864 30200
rect 20548 29974 20668 30002
rect 20444 29096 20496 29102
rect 20444 29038 20496 29044
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20260 27668 20312 27674
rect 20260 27610 20312 27616
rect 20074 26415 20130 26424
rect 20168 26444 20220 26450
rect 20088 26382 20116 26415
rect 20168 26386 20220 26392
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 20168 25356 20220 25362
rect 20168 25298 20220 25304
rect 19996 25214 20116 25242
rect 19798 25191 19800 25200
rect 19852 25191 19854 25200
rect 19800 25162 19852 25168
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23798 20024 25094
rect 20088 24886 20116 25214
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 20180 24721 20208 25298
rect 20166 24712 20222 24721
rect 20166 24647 20222 24656
rect 20272 24562 20300 27610
rect 20364 26382 20392 28494
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20088 24534 20300 24562
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19260 20942 19288 21422
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19800 21004 19852 21010
rect 19800 20946 19852 20952
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19812 20874 19840 20946
rect 19904 20874 19932 21286
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 19892 20868 19944 20874
rect 19892 20810 19944 20816
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19076 19306 19196 19334
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18800 15706 18828 15846
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18800 14906 18828 14962
rect 19076 14929 19104 19306
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19168 16182 19196 16934
rect 19156 16176 19208 16182
rect 19156 16118 19208 16124
rect 18524 14878 18828 14906
rect 19062 14920 19118 14929
rect 19062 14855 19118 14864
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18432 14006 18460 14758
rect 18708 14346 18736 14758
rect 18696 14340 18748 14346
rect 18696 14282 18748 14288
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18064 13462 18092 13738
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 19076 12918 19104 14855
rect 19260 14550 19288 19450
rect 19444 18970 19472 19722
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19996 18850 20024 23598
rect 20088 22030 20116 24534
rect 20364 24206 20392 26318
rect 20444 26308 20496 26314
rect 20444 26250 20496 26256
rect 20456 25974 20484 26250
rect 20548 25974 20576 29974
rect 20628 29504 20680 29510
rect 20628 29446 20680 29452
rect 20640 29238 20668 29446
rect 20628 29232 20680 29238
rect 20628 29174 20680 29180
rect 20824 28778 20852 30194
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 20916 29306 20944 29582
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 20824 28750 20944 28778
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20444 25968 20496 25974
rect 20444 25910 20496 25916
rect 20536 25968 20588 25974
rect 20536 25910 20588 25916
rect 20442 25256 20498 25265
rect 20442 25191 20444 25200
rect 20496 25191 20498 25200
rect 20444 25162 20496 25168
rect 20444 24744 20496 24750
rect 20444 24686 20496 24692
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20456 23746 20484 24686
rect 20640 24426 20668 28494
rect 20916 28490 20944 28750
rect 20904 28484 20956 28490
rect 20904 28426 20956 28432
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 20180 23718 20484 23746
rect 20548 24398 20668 24426
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20180 21962 20208 23718
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 19996 18822 20116 18850
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19352 17678 19380 18702
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19812 17746 19840 18022
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19444 17338 19472 17614
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19352 16250 19380 16458
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19352 16046 19380 16186
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19168 13870 19196 14282
rect 19260 14006 19288 14486
rect 19352 14278 19380 15846
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 14278 19472 15302
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19892 14000 19944 14006
rect 19892 13942 19944 13948
rect 19904 13870 19932 13942
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 19064 12912 19116 12918
rect 19064 12854 19116 12860
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17868 12708 17920 12714
rect 17868 12650 17920 12656
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17880 12238 17908 12650
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 18156 11830 18184 12310
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11830 18460 12038
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 18420 11824 18472 11830
rect 18420 11766 18472 11772
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18972 11688 19024 11694
rect 19076 11676 19104 12854
rect 19996 12434 20024 18702
rect 20088 16522 20116 18822
rect 20076 16516 20128 16522
rect 20076 16458 20128 16464
rect 20088 15978 20116 16458
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 20180 14822 20208 21898
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20272 19378 20300 19858
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20364 19514 20392 19790
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20272 15502 20300 19314
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19352 12406 20024 12434
rect 19352 12170 19380 12406
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19024 11648 19104 11676
rect 18972 11630 19024 11636
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17236 10810 17264 10950
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17328 10674 17356 10950
rect 18340 10810 18368 11630
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 9994 17448 10406
rect 17880 10266 17908 10542
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17972 10198 18000 10678
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 17052 3058 17080 7142
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16868 2446 16896 2790
rect 17512 2446 17540 7686
rect 18248 2650 18276 10542
rect 19352 10198 19380 12106
rect 19444 11014 19472 12174
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11830 20024 12038
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10266 20024 11154
rect 20088 11082 20116 12582
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 20180 10606 20208 11630
rect 20272 10810 20300 12106
rect 20364 11218 20392 13194
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 20456 10130 20484 23598
rect 20548 23322 20576 24398
rect 20626 24168 20682 24177
rect 20626 24103 20682 24112
rect 20720 24132 20772 24138
rect 20640 24070 20668 24103
rect 20720 24074 20772 24080
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20626 23624 20682 23633
rect 20626 23559 20682 23568
rect 20640 23526 20668 23559
rect 20732 23526 20760 24074
rect 20628 23520 20680 23526
rect 20628 23462 20680 23468
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20718 23352 20774 23361
rect 20536 23316 20588 23322
rect 20718 23287 20774 23296
rect 20536 23258 20588 23264
rect 20548 23186 20576 23258
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20732 23118 20760 23287
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20824 23050 20852 28018
rect 20812 23044 20864 23050
rect 20812 22986 20864 22992
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 19922 20576 20198
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20640 16182 20668 21830
rect 20916 21554 20944 28426
rect 21008 23186 21036 31726
rect 21088 30660 21140 30666
rect 21088 30602 21140 30608
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 20996 23044 21048 23050
rect 20996 22986 21048 22992
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20640 15910 20668 15982
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20640 15638 20668 15846
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20640 11626 20668 14758
rect 20732 14074 20760 20946
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 20824 18358 20852 18770
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20824 17610 20852 17682
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20824 13190 20852 17546
rect 20916 14958 20944 19858
rect 21008 15502 21036 22986
rect 21100 21010 21128 30602
rect 21180 25220 21232 25226
rect 21180 25162 21232 25168
rect 21192 24750 21220 25162
rect 21180 24744 21232 24750
rect 21180 24686 21232 24692
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 21008 14482 21036 14826
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20916 10674 20944 14350
rect 21192 12322 21220 24686
rect 21100 12294 21220 12322
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 20640 9722 20668 10542
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 7886 19380 9318
rect 20456 9042 20484 9454
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 20824 8090 20852 9454
rect 21008 8498 21036 11086
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 21008 7886 21036 8230
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 21100 7410 21128 12294
rect 21284 11694 21312 35566
rect 21456 35080 21508 35086
rect 21456 35022 21508 35028
rect 21468 32434 21496 35022
rect 21560 34542 21588 35702
rect 21548 34536 21600 34542
rect 21548 34478 21600 34484
rect 21548 33040 21600 33046
rect 21548 32982 21600 32988
rect 21456 32428 21508 32434
rect 21456 32370 21508 32376
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 21560 30682 21588 32982
rect 21652 31754 21680 36314
rect 22020 36258 22048 36518
rect 21836 36230 22048 36258
rect 21836 35222 21864 36230
rect 22112 36122 22140 36586
rect 22020 36094 22140 36122
rect 22020 35894 22048 36094
rect 22100 36032 22152 36038
rect 22152 35980 22232 35986
rect 22100 35974 22232 35980
rect 22112 35958 22232 35974
rect 22020 35866 22140 35894
rect 22112 35834 22140 35866
rect 22100 35828 22152 35834
rect 22100 35770 22152 35776
rect 22204 35698 22232 35958
rect 22296 35766 22324 36722
rect 22284 35760 22336 35766
rect 22284 35702 22336 35708
rect 22468 35760 22520 35766
rect 22468 35702 22520 35708
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 22100 35624 22152 35630
rect 22100 35566 22152 35572
rect 21824 35216 21876 35222
rect 21824 35158 21876 35164
rect 21824 35012 21876 35018
rect 21824 34954 21876 34960
rect 21730 34912 21786 34921
rect 21730 34847 21786 34856
rect 21744 32434 21772 34847
rect 21732 32428 21784 32434
rect 21732 32370 21784 32376
rect 21652 31726 21772 31754
rect 21468 29186 21496 30670
rect 21560 30654 21680 30682
rect 21546 29880 21602 29889
rect 21546 29815 21548 29824
rect 21600 29815 21602 29824
rect 21548 29786 21600 29792
rect 21652 29714 21680 30654
rect 21640 29708 21692 29714
rect 21640 29650 21692 29656
rect 21468 29170 21680 29186
rect 21468 29164 21692 29170
rect 21468 29158 21640 29164
rect 21640 29106 21692 29112
rect 21548 27668 21600 27674
rect 21548 27610 21600 27616
rect 21362 27568 21418 27577
rect 21362 27503 21364 27512
rect 21416 27503 21418 27512
rect 21364 27474 21416 27480
rect 21560 27441 21588 27610
rect 21546 27432 21602 27441
rect 21364 27396 21416 27402
rect 21546 27367 21602 27376
rect 21364 27338 21416 27344
rect 21376 26858 21404 27338
rect 21652 26926 21680 29106
rect 21640 26920 21692 26926
rect 21640 26862 21692 26868
rect 21364 26852 21416 26858
rect 21364 26794 21416 26800
rect 21640 26784 21692 26790
rect 21640 26726 21692 26732
rect 21652 25294 21680 26726
rect 21640 25288 21692 25294
rect 21640 25230 21692 25236
rect 21364 25220 21416 25226
rect 21364 25162 21416 25168
rect 21376 22710 21404 25162
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21364 22704 21416 22710
rect 21364 22646 21416 22652
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21376 17746 21404 18022
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21364 15428 21416 15434
rect 21364 15370 21416 15376
rect 21376 15026 21404 15370
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21468 13326 21496 24142
rect 21652 23662 21680 24754
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 21744 22094 21772 31726
rect 21836 31346 21864 34954
rect 22112 34746 22140 35566
rect 22284 35488 22336 35494
rect 22284 35430 22336 35436
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 22296 34474 22324 35430
rect 22388 35086 22416 35634
rect 22480 35562 22508 35702
rect 22468 35556 22520 35562
rect 22468 35498 22520 35504
rect 22376 35080 22428 35086
rect 22376 35022 22428 35028
rect 22388 34610 22416 35022
rect 22468 34672 22520 34678
rect 22466 34640 22468 34649
rect 22520 34640 22522 34649
rect 22376 34604 22428 34610
rect 22466 34575 22522 34584
rect 22376 34546 22428 34552
rect 22284 34468 22336 34474
rect 22284 34410 22336 34416
rect 22388 33998 22416 34546
rect 22572 34524 22600 37198
rect 22652 36916 22704 36922
rect 22652 36858 22704 36864
rect 22664 36378 22692 36858
rect 22744 36780 22796 36786
rect 22744 36722 22796 36728
rect 22652 36372 22704 36378
rect 22652 36314 22704 36320
rect 22480 34496 22600 34524
rect 22376 33992 22428 33998
rect 22098 33960 22154 33969
rect 22376 33934 22428 33940
rect 22098 33895 22154 33904
rect 22112 33561 22140 33895
rect 22098 33552 22154 33561
rect 22098 33487 22154 33496
rect 22006 33008 22062 33017
rect 22006 32943 22062 32952
rect 22020 32774 22048 32943
rect 22112 32842 22140 33487
rect 22282 33416 22338 33425
rect 22282 33351 22338 33360
rect 22190 33008 22246 33017
rect 22190 32943 22246 32952
rect 22100 32836 22152 32842
rect 22100 32778 22152 32784
rect 22204 32774 22232 32943
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 22192 32768 22244 32774
rect 22192 32710 22244 32716
rect 21916 32428 21968 32434
rect 21916 32370 21968 32376
rect 21824 31340 21876 31346
rect 21824 31282 21876 31288
rect 21928 30682 21956 32370
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22112 32026 22140 32166
rect 22100 32020 22152 32026
rect 22100 31962 22152 31968
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 22192 31884 22244 31890
rect 22192 31826 22244 31832
rect 21836 30666 21956 30682
rect 21824 30660 21956 30666
rect 21876 30654 21956 30660
rect 21824 30602 21876 30608
rect 21836 28558 21864 30602
rect 22020 30172 22048 31826
rect 22204 31521 22232 31826
rect 22190 31512 22246 31521
rect 22190 31447 22246 31456
rect 22192 31272 22244 31278
rect 22192 31214 22244 31220
rect 22020 30144 22140 30172
rect 22112 30054 22140 30144
rect 22100 30048 22152 30054
rect 22100 29990 22152 29996
rect 22112 28762 22140 29990
rect 22100 28756 22152 28762
rect 22100 28698 22152 28704
rect 22204 28608 22232 31214
rect 22296 31210 22324 33351
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22388 31686 22416 32846
rect 22480 32745 22508 34496
rect 22560 34400 22612 34406
rect 22560 34342 22612 34348
rect 22572 33318 22600 34342
rect 22756 33522 22784 36722
rect 22836 34944 22888 34950
rect 22836 34886 22888 34892
rect 22928 34944 22980 34950
rect 22928 34886 22980 34892
rect 22848 33930 22876 34886
rect 22836 33924 22888 33930
rect 22836 33866 22888 33872
rect 22744 33516 22796 33522
rect 22744 33458 22796 33464
rect 22940 33454 22968 34886
rect 23124 34626 23152 37198
rect 23216 37182 23428 37198
rect 23216 36786 23244 37182
rect 24504 37126 24532 39200
rect 25044 37460 25096 37466
rect 25044 37402 25096 37408
rect 25056 37262 25084 37402
rect 25044 37256 25096 37262
rect 25044 37198 25096 37204
rect 23388 37120 23440 37126
rect 23388 37062 23440 37068
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 23400 36174 23428 37062
rect 24214 36952 24270 36961
rect 24214 36887 24270 36896
rect 24228 36854 24256 36887
rect 24216 36848 24268 36854
rect 24216 36790 24268 36796
rect 23940 36712 23992 36718
rect 23940 36654 23992 36660
rect 24032 36712 24084 36718
rect 24032 36654 24084 36660
rect 23388 36168 23440 36174
rect 23388 36110 23440 36116
rect 23480 36168 23532 36174
rect 23480 36110 23532 36116
rect 23492 35698 23520 36110
rect 23480 35692 23532 35698
rect 23480 35634 23532 35640
rect 23492 35086 23520 35634
rect 23480 35080 23532 35086
rect 23480 35022 23532 35028
rect 23664 35080 23716 35086
rect 23664 35022 23716 35028
rect 23020 34604 23072 34610
rect 23124 34598 23244 34626
rect 23400 34610 23612 34626
rect 23020 34546 23072 34552
rect 22928 33448 22980 33454
rect 22928 33390 22980 33396
rect 22560 33312 22612 33318
rect 22560 33254 22612 33260
rect 22652 33312 22704 33318
rect 22652 33254 22704 33260
rect 22466 32736 22522 32745
rect 22466 32671 22522 32680
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 22284 31204 22336 31210
rect 22284 31146 22336 31152
rect 22376 30184 22428 30190
rect 22376 30126 22428 30132
rect 22388 30054 22416 30126
rect 22376 30048 22428 30054
rect 22376 29990 22428 29996
rect 22376 29504 22428 29510
rect 22376 29446 22428 29452
rect 22284 29300 22336 29306
rect 22284 29242 22336 29248
rect 21928 28580 22232 28608
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21928 28404 21956 28580
rect 22296 28558 22324 29242
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22008 28484 22060 28490
rect 22008 28426 22060 28432
rect 21836 28376 21956 28404
rect 21836 27606 21864 28376
rect 21914 27976 21970 27985
rect 21914 27911 21916 27920
rect 21968 27911 21970 27920
rect 21916 27882 21968 27888
rect 21824 27600 21876 27606
rect 21824 27542 21876 27548
rect 22020 27554 22048 28426
rect 22296 28150 22324 28494
rect 22284 28144 22336 28150
rect 22284 28086 22336 28092
rect 22020 27526 22140 27554
rect 21822 27432 21878 27441
rect 21822 27367 21878 27376
rect 22008 27396 22060 27402
rect 21836 27334 21864 27367
rect 22008 27338 22060 27344
rect 21824 27328 21876 27334
rect 21824 27270 21876 27276
rect 22020 27130 22048 27338
rect 22112 27130 22140 27526
rect 22008 27124 22060 27130
rect 22008 27066 22060 27072
rect 22100 27124 22152 27130
rect 22100 27066 22152 27072
rect 22284 26240 22336 26246
rect 22284 26182 22336 26188
rect 22296 25906 22324 26182
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 21916 25152 21968 25158
rect 21916 25094 21968 25100
rect 21928 24206 21956 25094
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 22112 24290 22140 24550
rect 22204 24410 22232 24754
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 22112 24262 22232 24290
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21836 23866 21864 24142
rect 22204 24138 22232 24262
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 22296 23254 22324 25230
rect 22100 23248 22152 23254
rect 22100 23190 22152 23196
rect 22284 23248 22336 23254
rect 22284 23190 22336 23196
rect 21916 23180 21968 23186
rect 21916 23122 21968 23128
rect 21652 22066 21772 22094
rect 21652 19990 21680 22066
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 21640 19984 21692 19990
rect 21836 19961 21864 20402
rect 21640 19926 21692 19932
rect 21822 19952 21878 19961
rect 21822 19887 21878 19896
rect 21640 18692 21692 18698
rect 21640 18634 21692 18640
rect 21652 14414 21680 18634
rect 21732 18352 21784 18358
rect 21732 18294 21784 18300
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21744 11762 21772 18294
rect 21928 18290 21956 23122
rect 22112 22030 22140 23190
rect 22388 22094 22416 29446
rect 22480 29170 22508 32370
rect 22560 32360 22612 32366
rect 22560 32302 22612 32308
rect 22572 31754 22600 32302
rect 22560 31748 22612 31754
rect 22560 31690 22612 31696
rect 22664 31278 22692 33254
rect 22928 32904 22980 32910
rect 22928 32846 22980 32852
rect 22744 32496 22796 32502
rect 22744 32438 22796 32444
rect 22756 31793 22784 32438
rect 22940 32434 22968 32846
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 22836 31884 22888 31890
rect 22836 31826 22888 31832
rect 22742 31784 22798 31793
rect 22742 31719 22798 31728
rect 22652 31272 22704 31278
rect 22652 31214 22704 31220
rect 22650 31104 22706 31113
rect 22650 31039 22706 31048
rect 22664 30394 22692 31039
rect 22652 30388 22704 30394
rect 22652 30330 22704 30336
rect 22560 29504 22612 29510
rect 22560 29446 22612 29452
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22480 27062 22508 29106
rect 22572 28218 22600 29446
rect 22560 28212 22612 28218
rect 22560 28154 22612 28160
rect 22468 27056 22520 27062
rect 22468 26998 22520 27004
rect 22480 26382 22508 26998
rect 22664 26382 22692 30330
rect 22848 27554 22876 31826
rect 22928 31680 22980 31686
rect 22928 31622 22980 31628
rect 22940 31414 22968 31622
rect 22928 31408 22980 31414
rect 22928 31350 22980 31356
rect 23032 30648 23060 34546
rect 23112 34536 23164 34542
rect 23112 34478 23164 34484
rect 23124 34105 23152 34478
rect 23216 34474 23244 34598
rect 23388 34604 23612 34610
rect 23440 34598 23612 34604
rect 23388 34546 23440 34552
rect 23480 34536 23532 34542
rect 23294 34504 23350 34513
rect 23204 34468 23256 34474
rect 23480 34478 23532 34484
rect 23294 34439 23350 34448
rect 23204 34410 23256 34416
rect 23110 34096 23166 34105
rect 23110 34031 23166 34040
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 23124 32910 23152 33458
rect 23308 33153 23336 34439
rect 23492 33969 23520 34478
rect 23584 34474 23612 34598
rect 23572 34468 23624 34474
rect 23572 34410 23624 34416
rect 23572 34128 23624 34134
rect 23572 34070 23624 34076
rect 23478 33960 23534 33969
rect 23478 33895 23534 33904
rect 23492 33522 23520 33895
rect 23480 33516 23532 33522
rect 23480 33458 23532 33464
rect 23294 33144 23350 33153
rect 23294 33079 23350 33088
rect 23204 33040 23256 33046
rect 23204 32982 23256 32988
rect 23112 32904 23164 32910
rect 23112 32846 23164 32852
rect 23216 32366 23244 32982
rect 23296 32496 23348 32502
rect 23296 32438 23348 32444
rect 23204 32360 23256 32366
rect 23204 32302 23256 32308
rect 23112 32224 23164 32230
rect 23112 32166 23164 32172
rect 23124 31890 23152 32166
rect 23308 32026 23336 32438
rect 23296 32020 23348 32026
rect 23296 31962 23348 31968
rect 23388 31952 23440 31958
rect 23440 31900 23520 31906
rect 23388 31894 23520 31900
rect 23112 31884 23164 31890
rect 23400 31878 23520 31894
rect 23112 31826 23164 31832
rect 23388 31748 23440 31754
rect 23388 31690 23440 31696
rect 23112 31680 23164 31686
rect 23112 31622 23164 31628
rect 23124 31482 23152 31622
rect 23112 31476 23164 31482
rect 23112 31418 23164 31424
rect 23112 30660 23164 30666
rect 23032 30620 23112 30648
rect 23112 30602 23164 30608
rect 23124 29646 23152 30602
rect 23400 29753 23428 31690
rect 23492 31346 23520 31878
rect 23584 31482 23612 34070
rect 23676 32774 23704 35022
rect 23952 34746 23980 36654
rect 24044 36106 24072 36654
rect 25148 36242 25176 39200
rect 25412 37392 25464 37398
rect 25412 37334 25464 37340
rect 26240 37392 26292 37398
rect 26240 37334 26292 37340
rect 25228 37188 25280 37194
rect 25228 37130 25280 37136
rect 25320 37188 25372 37194
rect 25320 37130 25372 37136
rect 25240 36922 25268 37130
rect 25228 36916 25280 36922
rect 25228 36858 25280 36864
rect 25240 36553 25268 36858
rect 25226 36544 25282 36553
rect 25226 36479 25282 36488
rect 25136 36236 25188 36242
rect 25136 36178 25188 36184
rect 24032 36100 24084 36106
rect 24032 36042 24084 36048
rect 24676 36100 24728 36106
rect 24676 36042 24728 36048
rect 24768 36100 24820 36106
rect 24768 36042 24820 36048
rect 24582 36000 24638 36009
rect 24582 35935 24638 35944
rect 24596 35698 24624 35935
rect 24688 35834 24716 36042
rect 24676 35828 24728 35834
rect 24676 35770 24728 35776
rect 24584 35692 24636 35698
rect 24584 35634 24636 35640
rect 24780 35290 24808 36042
rect 24768 35284 24820 35290
rect 24768 35226 24820 35232
rect 23940 34740 23992 34746
rect 23940 34682 23992 34688
rect 25044 34740 25096 34746
rect 25044 34682 25096 34688
rect 23848 34604 23900 34610
rect 23848 34546 23900 34552
rect 23756 34536 23808 34542
rect 23754 34504 23756 34513
rect 23808 34504 23810 34513
rect 23754 34439 23810 34448
rect 23664 32768 23716 32774
rect 23664 32710 23716 32716
rect 23572 31476 23624 31482
rect 23572 31418 23624 31424
rect 23480 31340 23532 31346
rect 23480 31282 23532 31288
rect 23664 31340 23716 31346
rect 23664 31282 23716 31288
rect 23572 31272 23624 31278
rect 23676 31249 23704 31282
rect 23860 31278 23888 34546
rect 24400 34400 24452 34406
rect 24400 34342 24452 34348
rect 23940 34060 23992 34066
rect 23940 34002 23992 34008
rect 23952 33590 23980 34002
rect 24412 33590 24440 34342
rect 24952 34060 25004 34066
rect 24952 34002 25004 34008
rect 24492 33992 24544 33998
rect 24492 33934 24544 33940
rect 24504 33658 24532 33934
rect 24492 33652 24544 33658
rect 24492 33594 24544 33600
rect 23940 33584 23992 33590
rect 23940 33526 23992 33532
rect 24308 33584 24360 33590
rect 24308 33526 24360 33532
rect 24400 33584 24452 33590
rect 24400 33526 24452 33532
rect 23952 33114 23980 33526
rect 24032 33516 24084 33522
rect 24032 33458 24084 33464
rect 23940 33108 23992 33114
rect 23940 33050 23992 33056
rect 23848 31272 23900 31278
rect 23572 31214 23624 31220
rect 23662 31240 23718 31249
rect 23584 31142 23612 31214
rect 23718 31198 23796 31226
rect 23848 31214 23900 31220
rect 23662 31175 23718 31184
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23768 30734 23796 31198
rect 24044 30870 24072 33458
rect 24124 33040 24176 33046
rect 24124 32982 24176 32988
rect 24136 32298 24164 32982
rect 24320 32978 24348 33526
rect 24860 33312 24912 33318
rect 24860 33254 24912 33260
rect 24308 32972 24360 32978
rect 24308 32914 24360 32920
rect 24492 32768 24544 32774
rect 24492 32710 24544 32716
rect 24124 32292 24176 32298
rect 24124 32234 24176 32240
rect 24400 31476 24452 31482
rect 24400 31418 24452 31424
rect 24032 30864 24084 30870
rect 24032 30806 24084 30812
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23664 30320 23716 30326
rect 23664 30262 23716 30268
rect 24124 30320 24176 30326
rect 24124 30262 24176 30268
rect 23386 29744 23442 29753
rect 23386 29679 23442 29688
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23124 29306 23152 29582
rect 23388 29572 23440 29578
rect 23388 29514 23440 29520
rect 23112 29300 23164 29306
rect 23112 29242 23164 29248
rect 23400 29102 23428 29514
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 23204 28756 23256 28762
rect 23204 28698 23256 28704
rect 23216 28014 23244 28698
rect 23204 28008 23256 28014
rect 23204 27950 23256 27956
rect 22848 27526 23060 27554
rect 22928 27396 22980 27402
rect 22928 27338 22980 27344
rect 22744 26444 22796 26450
rect 22744 26386 22796 26392
rect 22468 26376 22520 26382
rect 22652 26376 22704 26382
rect 22520 26324 22600 26330
rect 22468 26318 22600 26324
rect 22652 26318 22704 26324
rect 22480 26302 22600 26318
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 22480 24750 22508 25774
rect 22572 24818 22600 26302
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 22560 24200 22612 24206
rect 22756 24154 22784 26386
rect 22836 26376 22888 26382
rect 22836 26318 22888 26324
rect 22848 24682 22876 26318
rect 22836 24676 22888 24682
rect 22836 24618 22888 24624
rect 22836 24336 22888 24342
rect 22836 24278 22888 24284
rect 22560 24142 22612 24148
rect 22572 23798 22600 24142
rect 22664 24126 22784 24154
rect 22560 23792 22612 23798
rect 22560 23734 22612 23740
rect 22468 23656 22520 23662
rect 22664 23644 22692 24126
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22468 23598 22520 23604
rect 22572 23616 22692 23644
rect 22296 22066 22416 22094
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 21412 22060 21418
rect 22008 21354 22060 21360
rect 22020 21078 22048 21354
rect 22008 21072 22060 21078
rect 22008 21014 22060 21020
rect 22020 20466 22048 21014
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 22112 18290 22140 20198
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22100 16584 22152 16590
rect 21822 16552 21878 16561
rect 22100 16526 22152 16532
rect 21822 16487 21878 16496
rect 21836 15094 21864 16487
rect 22112 16250 22140 16526
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21928 14958 21956 15914
rect 22020 15706 22048 16050
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 22020 15042 22048 15302
rect 22100 15088 22152 15094
rect 22020 15036 22100 15042
rect 22020 15030 22152 15036
rect 22020 15014 22140 15030
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 12170 22140 12582
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21744 11150 21772 11698
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21180 11008 21232 11014
rect 21180 10950 21232 10956
rect 21192 10674 21220 10950
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21192 9722 21220 10406
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 19996 2446 20024 7210
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20640 2514 20668 2790
rect 22020 2650 22048 9998
rect 22204 6914 22232 20266
rect 22296 13734 22324 22066
rect 22480 19174 22508 23598
rect 22572 20534 22600 23616
rect 22756 23050 22784 24006
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 22664 19990 22692 22986
rect 22652 19984 22704 19990
rect 22652 19926 22704 19932
rect 22848 19786 22876 24278
rect 22940 23662 22968 27338
rect 22928 23656 22980 23662
rect 22926 23624 22928 23633
rect 22980 23624 22982 23633
rect 22926 23559 22982 23568
rect 23032 23050 23060 27526
rect 23216 26926 23244 27950
rect 23296 27940 23348 27946
rect 23296 27882 23348 27888
rect 23204 26920 23256 26926
rect 23204 26862 23256 26868
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23124 24954 23152 25230
rect 23112 24948 23164 24954
rect 23112 24890 23164 24896
rect 23124 24342 23152 24890
rect 23112 24336 23164 24342
rect 23112 24278 23164 24284
rect 23112 24200 23164 24206
rect 23110 24168 23112 24177
rect 23164 24168 23166 24177
rect 23110 24103 23166 24112
rect 23216 23474 23244 26862
rect 23308 25430 23336 27882
rect 23386 27568 23442 27577
rect 23386 27503 23442 27512
rect 23400 27470 23428 27503
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23296 25424 23348 25430
rect 23296 25366 23348 25372
rect 23400 24750 23428 26318
rect 23492 25974 23520 27270
rect 23480 25968 23532 25974
rect 23480 25910 23532 25916
rect 23676 25498 23704 30262
rect 24032 30048 24084 30054
rect 24032 29990 24084 29996
rect 23756 29640 23808 29646
rect 23754 29608 23756 29617
rect 23808 29608 23810 29617
rect 23754 29543 23810 29552
rect 23756 29504 23808 29510
rect 23756 29446 23808 29452
rect 23940 29504 23992 29510
rect 23940 29446 23992 29452
rect 23768 28150 23796 29446
rect 23952 29306 23980 29446
rect 23940 29300 23992 29306
rect 23940 29242 23992 29248
rect 24044 29034 24072 29990
rect 24032 29028 24084 29034
rect 24032 28970 24084 28976
rect 23940 28484 23992 28490
rect 23940 28426 23992 28432
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23848 26920 23900 26926
rect 23848 26862 23900 26868
rect 23860 26353 23888 26862
rect 23952 26586 23980 28426
rect 24044 28014 24072 28970
rect 24136 28490 24164 30262
rect 24124 28484 24176 28490
rect 24124 28426 24176 28432
rect 24032 28008 24084 28014
rect 24032 27950 24084 27956
rect 23940 26580 23992 26586
rect 23940 26522 23992 26528
rect 23846 26344 23902 26353
rect 23846 26279 23902 26288
rect 23664 25492 23716 25498
rect 23664 25434 23716 25440
rect 24044 25378 24072 27950
rect 23676 25350 24072 25378
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23492 24818 23520 25230
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23584 24886 23612 25094
rect 23572 24880 23624 24886
rect 23572 24822 23624 24828
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 23296 24064 23348 24070
rect 23296 24006 23348 24012
rect 23124 23446 23244 23474
rect 23020 23044 23072 23050
rect 23020 22986 23072 22992
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22836 19780 22888 19786
rect 22836 19722 22888 19728
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22376 17060 22428 17066
rect 22376 17002 22428 17008
rect 22388 13818 22416 17002
rect 22480 16538 22508 19110
rect 22756 18970 22784 19722
rect 23124 19446 23152 23446
rect 23308 22094 23336 24006
rect 23400 23526 23428 24686
rect 23388 23520 23440 23526
rect 23388 23462 23440 23468
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23216 22066 23336 22094
rect 23388 22092 23440 22098
rect 23112 19440 23164 19446
rect 23112 19382 23164 19388
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 22756 18426 22784 18906
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22756 17882 22784 18362
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22480 16510 22876 16538
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22480 15502 22508 16118
rect 22572 15706 22600 16186
rect 22664 15706 22692 16390
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22480 13938 22508 14350
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22388 13790 22508 13818
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22296 12434 22324 13670
rect 22296 12406 22416 12434
rect 22388 12170 22416 12406
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22480 11150 22508 13790
rect 22756 12306 22784 16390
rect 22848 14940 22876 16510
rect 22940 16182 22968 18566
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 22928 16176 22980 16182
rect 22928 16118 22980 16124
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22940 15434 22968 15846
rect 23032 15450 23060 17614
rect 23124 17338 23152 18906
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23216 16522 23244 22066
rect 23388 22034 23440 22040
rect 23400 21554 23428 22034
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23492 21434 23520 22918
rect 23676 22094 23704 25350
rect 23848 25220 23900 25226
rect 23848 25162 23900 25168
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23400 21406 23520 21434
rect 23584 22066 23704 22094
rect 23204 16516 23256 16522
rect 23204 16458 23256 16464
rect 23400 16402 23428 21406
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23492 16561 23520 20334
rect 23478 16552 23534 16561
rect 23478 16487 23534 16496
rect 23216 16374 23428 16402
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23124 15570 23152 15846
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 23032 15434 23152 15450
rect 22928 15428 22980 15434
rect 23032 15428 23164 15434
rect 23032 15422 23112 15428
rect 22928 15370 22980 15376
rect 23112 15370 23164 15376
rect 22928 14952 22980 14958
rect 22848 14912 22928 14940
rect 22928 14894 22980 14900
rect 23124 12986 23152 15370
rect 23216 13462 23244 16374
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23584 16130 23612 22066
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23676 20602 23704 20878
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23768 20534 23796 23462
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23860 19378 23888 25162
rect 23940 23044 23992 23050
rect 23940 22986 23992 22992
rect 23848 19372 23900 19378
rect 23848 19314 23900 19320
rect 23204 13456 23256 13462
rect 23204 13398 23256 13404
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 23308 12918 23336 16118
rect 23584 16102 23704 16130
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23492 15366 23520 15914
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23400 13258 23428 14214
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 23308 12306 23336 12718
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 22756 12102 22784 12242
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22848 11558 22876 12174
rect 23020 11688 23072 11694
rect 23020 11630 23072 11636
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22480 10674 22508 11086
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22296 10266 22324 10542
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 23032 10198 23060 11630
rect 23204 11620 23256 11626
rect 23204 11562 23256 11568
rect 23216 11286 23244 11562
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 23492 10810 23520 15302
rect 23584 15094 23612 15982
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23676 14550 23704 16102
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23572 14340 23624 14346
rect 23572 14282 23624 14288
rect 23584 12782 23612 14282
rect 23572 12776 23624 12782
rect 23572 12718 23624 12724
rect 23584 11762 23612 12718
rect 23952 12434 23980 22986
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 24044 19990 24072 20334
rect 24032 19984 24084 19990
rect 24032 19926 24084 19932
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 24044 18426 24072 19314
rect 24032 18420 24084 18426
rect 24032 18362 24084 18368
rect 24030 17640 24086 17649
rect 24030 17575 24032 17584
rect 24084 17575 24086 17584
rect 24032 17546 24084 17552
rect 24136 14618 24164 28426
rect 24216 27328 24268 27334
rect 24216 27270 24268 27276
rect 24228 27062 24256 27270
rect 24216 27056 24268 27062
rect 24216 26998 24268 27004
rect 24216 26852 24268 26858
rect 24216 26794 24268 26800
rect 24228 25838 24256 26794
rect 24216 25832 24268 25838
rect 24216 25774 24268 25780
rect 24308 25832 24360 25838
rect 24308 25774 24360 25780
rect 24228 24954 24256 25774
rect 24216 24948 24268 24954
rect 24216 24890 24268 24896
rect 24320 22574 24348 25774
rect 24412 23118 24440 31418
rect 24504 29322 24532 32710
rect 24872 32502 24900 33254
rect 24964 32881 24992 34002
rect 25056 33454 25084 34682
rect 25332 34542 25360 37130
rect 25424 35698 25452 37334
rect 25872 36780 25924 36786
rect 25872 36722 25924 36728
rect 25884 36689 25912 36722
rect 25870 36680 25926 36689
rect 25870 36615 25872 36624
rect 25924 36615 25926 36624
rect 25872 36586 25924 36592
rect 25884 36555 25912 36586
rect 26252 36106 26280 37334
rect 26332 36780 26384 36786
rect 26332 36722 26384 36728
rect 26344 36417 26372 36722
rect 26436 36666 26464 39200
rect 26608 37256 26660 37262
rect 26608 37198 26660 37204
rect 26620 36922 26648 37198
rect 27724 37126 27752 39200
rect 27804 37256 27856 37262
rect 27804 37198 27856 37204
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 27816 36922 27844 37198
rect 26608 36916 26660 36922
rect 26608 36858 26660 36864
rect 27804 36916 27856 36922
rect 27804 36858 27856 36864
rect 27896 36916 27948 36922
rect 27896 36858 27948 36864
rect 27436 36848 27488 36854
rect 27264 36796 27436 36802
rect 27908 36802 27936 36858
rect 27264 36790 27488 36796
rect 27264 36786 27476 36790
rect 26608 36780 26660 36786
rect 26608 36722 26660 36728
rect 27252 36780 27476 36786
rect 27304 36774 27476 36780
rect 27724 36774 27936 36802
rect 28078 36816 28134 36825
rect 27252 36722 27304 36728
rect 26436 36638 26556 36666
rect 26424 36576 26476 36582
rect 26424 36518 26476 36524
rect 26330 36408 26386 36417
rect 26330 36343 26386 36352
rect 25504 36100 25556 36106
rect 25504 36042 25556 36048
rect 25964 36100 26016 36106
rect 25964 36042 26016 36048
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 25412 35692 25464 35698
rect 25412 35634 25464 35640
rect 25228 34536 25280 34542
rect 25228 34478 25280 34484
rect 25320 34536 25372 34542
rect 25320 34478 25372 34484
rect 25044 33448 25096 33454
rect 25044 33390 25096 33396
rect 24950 32872 25006 32881
rect 24950 32807 25006 32816
rect 24952 32768 25004 32774
rect 24952 32710 25004 32716
rect 24860 32496 24912 32502
rect 24860 32438 24912 32444
rect 24964 32366 24992 32710
rect 24952 32360 25004 32366
rect 24952 32302 25004 32308
rect 24860 32292 24912 32298
rect 24860 32234 24912 32240
rect 24768 31816 24820 31822
rect 24766 31784 24768 31793
rect 24820 31784 24822 31793
rect 24766 31719 24822 31728
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24780 29578 24808 31078
rect 24872 29594 24900 32234
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 24964 30938 24992 31282
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 25056 30190 25084 33390
rect 25136 32972 25188 32978
rect 25136 32914 25188 32920
rect 25044 30184 25096 30190
rect 25044 30126 25096 30132
rect 24872 29578 24992 29594
rect 24768 29572 24820 29578
rect 24872 29572 25004 29578
rect 24872 29566 24952 29572
rect 24768 29514 24820 29520
rect 24952 29514 25004 29520
rect 24504 29294 24808 29322
rect 24676 29232 24728 29238
rect 24676 29174 24728 29180
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24504 27062 24532 28358
rect 24688 27606 24716 29174
rect 24780 27606 24808 29294
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 24858 27976 24914 27985
rect 24858 27911 24860 27920
rect 24912 27911 24914 27920
rect 24860 27882 24912 27888
rect 24676 27600 24728 27606
rect 24676 27542 24728 27548
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24584 27464 24636 27470
rect 24780 27418 24808 27542
rect 24584 27406 24636 27412
rect 24492 27056 24544 27062
rect 24492 26998 24544 27004
rect 24596 26790 24624 27406
rect 24688 27390 24808 27418
rect 24860 27464 24912 27470
rect 24860 27406 24912 27412
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24504 26194 24532 26318
rect 24504 26166 24624 26194
rect 24492 26036 24544 26042
rect 24492 25978 24544 25984
rect 24504 25226 24532 25978
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24400 22976 24452 22982
rect 24400 22918 24452 22924
rect 24412 22710 24440 22918
rect 24400 22704 24452 22710
rect 24400 22646 24452 22652
rect 24308 22568 24360 22574
rect 24308 22510 24360 22516
rect 24320 22094 24348 22510
rect 24228 22066 24348 22094
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 23952 12406 24164 12434
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23768 11150 23796 11834
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23860 10606 23888 11018
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 23112 10464 23164 10470
rect 23112 10406 23164 10412
rect 23020 10192 23072 10198
rect 23020 10134 23072 10140
rect 23124 10062 23152 10406
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23860 8974 23888 10542
rect 24136 9586 24164 12406
rect 24228 11286 24256 22066
rect 24492 18284 24544 18290
rect 24492 18226 24544 18232
rect 24308 14884 24360 14890
rect 24308 14826 24360 14832
rect 24320 12374 24348 14826
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24412 14074 24440 14350
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 24308 12368 24360 12374
rect 24308 12310 24360 12316
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 22204 6886 22324 6914
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22296 2582 22324 6886
rect 24504 6254 24532 18226
rect 24596 16250 24624 26166
rect 24688 23730 24716 27390
rect 24768 27328 24820 27334
rect 24872 27316 24900 27406
rect 24820 27288 24900 27316
rect 24768 27270 24820 27276
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 24768 26308 24820 26314
rect 24768 26250 24820 26256
rect 24780 25226 24808 26250
rect 24964 26246 24992 26862
rect 25056 26382 25084 28018
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 24952 26240 25004 26246
rect 24952 26182 25004 26188
rect 24768 25220 24820 25226
rect 24768 25162 24820 25168
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24872 24138 24900 25094
rect 24964 24886 24992 26182
rect 24952 24880 25004 24886
rect 24952 24822 25004 24828
rect 24950 24712 25006 24721
rect 24950 24647 25006 24656
rect 24964 24274 24992 24647
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24780 23050 24808 23258
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24964 22710 24992 24210
rect 25148 23254 25176 32914
rect 25240 31385 25268 34478
rect 25516 34134 25544 36042
rect 25976 35834 26004 36042
rect 25964 35828 26016 35834
rect 25964 35770 26016 35776
rect 26436 35766 26464 36518
rect 26424 35760 26476 35766
rect 25778 35728 25834 35737
rect 25688 35692 25740 35698
rect 26424 35702 26476 35708
rect 25778 35663 25834 35672
rect 25688 35634 25740 35640
rect 25596 35080 25648 35086
rect 25596 35022 25648 35028
rect 25608 34610 25636 35022
rect 25596 34604 25648 34610
rect 25596 34546 25648 34552
rect 25504 34128 25556 34134
rect 25504 34070 25556 34076
rect 25412 34060 25464 34066
rect 25412 34002 25464 34008
rect 25424 33862 25452 34002
rect 25412 33856 25464 33862
rect 25412 33798 25464 33804
rect 25412 32836 25464 32842
rect 25412 32778 25464 32784
rect 25320 31816 25372 31822
rect 25320 31758 25372 31764
rect 25226 31376 25282 31385
rect 25226 31311 25282 31320
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 25240 27878 25268 29514
rect 25332 29238 25360 31758
rect 25320 29232 25372 29238
rect 25320 29174 25372 29180
rect 25228 27872 25280 27878
rect 25228 27814 25280 27820
rect 25320 27464 25372 27470
rect 25318 27432 25320 27441
rect 25372 27432 25374 27441
rect 25318 27367 25374 27376
rect 25320 26240 25372 26246
rect 25320 26182 25372 26188
rect 25332 25770 25360 26182
rect 25320 25764 25372 25770
rect 25320 25706 25372 25712
rect 25320 25492 25372 25498
rect 25320 25434 25372 25440
rect 25332 25294 25360 25434
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25136 23248 25188 23254
rect 25136 23190 25188 23196
rect 24952 22704 25004 22710
rect 24952 22646 25004 22652
rect 25148 22094 25176 23190
rect 25148 22066 25268 22094
rect 25136 21616 25188 21622
rect 25136 21558 25188 21564
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24584 15088 24636 15094
rect 24584 15030 24636 15036
rect 24596 14618 24624 15030
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24596 10062 24624 13874
rect 24780 11898 24808 19382
rect 24872 17814 24900 20402
rect 24950 19952 25006 19961
rect 24950 19887 25006 19896
rect 24964 19854 24992 19887
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24860 17808 24912 17814
rect 24860 17750 24912 17756
rect 24860 15904 24912 15910
rect 24860 15846 24912 15852
rect 24872 14958 24900 15846
rect 25056 15434 25084 19654
rect 25148 18630 25176 21558
rect 25240 20874 25268 22066
rect 25424 21690 25452 32778
rect 25516 32774 25544 34070
rect 25596 33992 25648 33998
rect 25594 33960 25596 33969
rect 25648 33960 25650 33969
rect 25594 33895 25650 33904
rect 25504 32768 25556 32774
rect 25504 32710 25556 32716
rect 25504 32224 25556 32230
rect 25504 32166 25556 32172
rect 25516 31793 25544 32166
rect 25502 31784 25558 31793
rect 25502 31719 25558 31728
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25516 31249 25544 31282
rect 25502 31240 25558 31249
rect 25502 31175 25558 31184
rect 25596 31204 25648 31210
rect 25516 30938 25544 31175
rect 25596 31146 25648 31152
rect 25504 30932 25556 30938
rect 25504 30874 25556 30880
rect 25608 30666 25636 31146
rect 25700 30682 25728 35634
rect 25792 31822 25820 35663
rect 26422 35456 26478 35465
rect 26422 35391 26478 35400
rect 26240 35148 26292 35154
rect 26240 35090 26292 35096
rect 26252 35057 26280 35090
rect 26238 35048 26294 35057
rect 26238 34983 26294 34992
rect 26436 34610 26464 35391
rect 26528 35290 26556 36638
rect 26516 35284 26568 35290
rect 26516 35226 26568 35232
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 25872 33856 25924 33862
rect 25872 33798 25924 33804
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 25792 31278 25820 31758
rect 25884 31686 25912 33798
rect 25964 33448 26016 33454
rect 25964 33390 26016 33396
rect 25976 33289 26004 33390
rect 25962 33280 26018 33289
rect 25962 33215 26018 33224
rect 26330 32600 26386 32609
rect 26330 32535 26332 32544
rect 26384 32535 26386 32544
rect 26332 32506 26384 32512
rect 25872 31680 25924 31686
rect 25872 31622 25924 31628
rect 26056 31408 26108 31414
rect 26056 31350 26108 31356
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25504 30660 25556 30666
rect 25504 30602 25556 30608
rect 25596 30660 25648 30666
rect 25700 30654 25820 30682
rect 25596 30602 25648 30608
rect 25516 30190 25544 30602
rect 25688 30592 25740 30598
rect 25688 30534 25740 30540
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25504 30184 25556 30190
rect 25504 30126 25556 30132
rect 25608 28490 25636 30194
rect 25596 28484 25648 28490
rect 25596 28426 25648 28432
rect 25700 28150 25728 30534
rect 25688 28144 25740 28150
rect 25688 28086 25740 28092
rect 25596 28008 25648 28014
rect 25596 27950 25648 27956
rect 25502 25392 25558 25401
rect 25502 25327 25558 25336
rect 25516 25294 25544 25327
rect 25504 25288 25556 25294
rect 25504 25230 25556 25236
rect 25608 24818 25636 27950
rect 25792 26489 25820 30654
rect 26068 30326 26096 31350
rect 26516 31136 26568 31142
rect 26516 31078 26568 31084
rect 26056 30320 26108 30326
rect 26056 30262 26108 30268
rect 26424 29232 26476 29238
rect 26424 29174 26476 29180
rect 26056 29096 26108 29102
rect 26056 29038 26108 29044
rect 25778 26480 25834 26489
rect 25778 26415 25834 26424
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 25504 24608 25556 24614
rect 25504 24550 25556 24556
rect 25516 24070 25544 24550
rect 25608 24410 25636 24754
rect 25596 24404 25648 24410
rect 25596 24346 25648 24352
rect 25688 24132 25740 24138
rect 25688 24074 25740 24080
rect 25504 24064 25556 24070
rect 25504 24006 25556 24012
rect 25596 24064 25648 24070
rect 25596 24006 25648 24012
rect 25516 23866 25544 24006
rect 25504 23860 25556 23866
rect 25504 23802 25556 23808
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25608 21622 25636 24006
rect 25700 23254 25728 24074
rect 25792 23730 25820 26415
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 25964 23520 26016 23526
rect 25964 23462 26016 23468
rect 25688 23248 25740 23254
rect 25688 23190 25740 23196
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25228 20868 25280 20874
rect 25228 20810 25280 20816
rect 25240 18902 25268 20810
rect 25700 19922 25728 23190
rect 25976 21962 26004 23462
rect 25964 21956 26016 21962
rect 25964 21898 26016 21904
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 25792 20534 25820 20742
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25228 18896 25280 18902
rect 25228 18838 25280 18844
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25136 16788 25188 16794
rect 25136 16730 25188 16736
rect 25044 15428 25096 15434
rect 25044 15370 25096 15376
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 24860 12708 24912 12714
rect 24860 12650 24912 12656
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24688 11218 24716 11630
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 24872 10674 24900 12650
rect 25148 11762 25176 16730
rect 26068 15434 26096 29038
rect 26436 28694 26464 29174
rect 26424 28688 26476 28694
rect 26424 28630 26476 28636
rect 26436 28218 26464 28630
rect 26424 28212 26476 28218
rect 26424 28154 26476 28160
rect 26528 28150 26556 31078
rect 26516 28144 26568 28150
rect 26516 28086 26568 28092
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 26436 26450 26464 27270
rect 26528 26926 26556 28086
rect 26516 26920 26568 26926
rect 26516 26862 26568 26868
rect 26424 26444 26476 26450
rect 26424 26386 26476 26392
rect 26516 26376 26568 26382
rect 26516 26318 26568 26324
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 26160 23866 26188 24142
rect 26148 23860 26200 23866
rect 26148 23802 26200 23808
rect 26424 22976 26476 22982
rect 26424 22918 26476 22924
rect 26436 22098 26464 22918
rect 26424 22092 26476 22098
rect 26424 22034 26476 22040
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26148 20392 26200 20398
rect 26148 20334 26200 20340
rect 26160 19922 26188 20334
rect 26148 19916 26200 19922
rect 26148 19858 26200 19864
rect 26252 19786 26280 21830
rect 26424 21412 26476 21418
rect 26424 21354 26476 21360
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26240 19780 26292 19786
rect 26240 19722 26292 19728
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26160 15570 26188 15982
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 25320 13252 25372 13258
rect 25320 13194 25372 13200
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 25240 11898 25268 12174
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24964 11354 24992 11494
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 25332 11082 25360 13194
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25700 11898 25728 12038
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 25044 11076 25096 11082
rect 25044 11018 25096 11024
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24492 6248 24544 6254
rect 24492 6190 24544 6196
rect 24688 2650 24716 10610
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24780 7886 24808 8774
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 24780 5234 24808 5510
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24676 2644 24728 2650
rect 24676 2586 24728 2592
rect 22284 2576 22336 2582
rect 22284 2518 22336 2524
rect 24872 2514 24900 10406
rect 25056 10266 25084 11018
rect 25332 10742 25360 11018
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 25792 3058 25820 12786
rect 26068 12442 26096 15370
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 26160 13258 26188 13806
rect 26344 13462 26372 21286
rect 26436 20874 26464 21354
rect 26424 20868 26476 20874
rect 26424 20810 26476 20816
rect 26424 20324 26476 20330
rect 26424 20266 26476 20272
rect 26436 15978 26464 20266
rect 26528 16590 26556 26318
rect 26620 25974 26648 36722
rect 27724 36718 27752 36774
rect 28078 36751 28134 36760
rect 28092 36718 28120 36751
rect 27712 36712 27764 36718
rect 27712 36654 27764 36660
rect 27804 36712 27856 36718
rect 27804 36654 27856 36660
rect 28080 36712 28132 36718
rect 28080 36654 28132 36660
rect 26700 36644 26752 36650
rect 26700 36586 26752 36592
rect 26712 36310 26740 36586
rect 27344 36576 27396 36582
rect 27344 36518 27396 36524
rect 26700 36304 26752 36310
rect 26700 36246 26752 36252
rect 26804 36242 27292 36258
rect 26804 36236 27304 36242
rect 26804 36230 27252 36236
rect 26700 34400 26752 34406
rect 26700 34342 26752 34348
rect 26712 33930 26740 34342
rect 26700 33924 26752 33930
rect 26700 33866 26752 33872
rect 26804 33810 26832 36230
rect 27252 36178 27304 36184
rect 27068 36100 27120 36106
rect 27068 36042 27120 36048
rect 26884 35624 26936 35630
rect 26884 35566 26936 35572
rect 26896 35018 26924 35566
rect 26884 35012 26936 35018
rect 26884 34954 26936 34960
rect 26896 34626 26924 34954
rect 26896 34598 27016 34626
rect 26884 34536 26936 34542
rect 26884 34478 26936 34484
rect 26712 33782 26832 33810
rect 26712 31142 26740 33782
rect 26792 33516 26844 33522
rect 26792 33458 26844 33464
rect 26804 33425 26832 33458
rect 26790 33416 26846 33425
rect 26790 33351 26846 33360
rect 26790 32736 26846 32745
rect 26790 32671 26846 32680
rect 26700 31136 26752 31142
rect 26700 31078 26752 31084
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 26712 29170 26740 30534
rect 26700 29164 26752 29170
rect 26700 29106 26752 29112
rect 26804 26908 26832 32671
rect 26896 31754 26924 34478
rect 26988 32978 27016 34598
rect 26976 32972 27028 32978
rect 26976 32914 27028 32920
rect 26976 32428 27028 32434
rect 26976 32370 27028 32376
rect 26988 31754 27016 32370
rect 26884 31748 26936 31754
rect 26884 31690 26936 31696
rect 26976 31748 27028 31754
rect 26976 31690 27028 31696
rect 27080 31634 27108 36042
rect 27160 35692 27212 35698
rect 27160 35634 27212 35640
rect 27172 35494 27200 35634
rect 27160 35488 27212 35494
rect 27160 35430 27212 35436
rect 27160 35012 27212 35018
rect 27160 34954 27212 34960
rect 26712 26880 26832 26908
rect 26896 31606 27108 31634
rect 26608 25968 26660 25974
rect 26608 25910 26660 25916
rect 26608 22568 26660 22574
rect 26608 22510 26660 22516
rect 26620 19922 26648 22510
rect 26712 21554 26740 26880
rect 26792 25424 26844 25430
rect 26792 25366 26844 25372
rect 26700 21548 26752 21554
rect 26700 21490 26752 21496
rect 26608 19916 26660 19922
rect 26608 19858 26660 19864
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26424 15972 26476 15978
rect 26424 15914 26476 15920
rect 26332 13456 26384 13462
rect 26332 13398 26384 13404
rect 26148 13252 26200 13258
rect 26148 13194 26200 13200
rect 26620 13190 26648 19858
rect 26608 13184 26660 13190
rect 26608 13126 26660 13132
rect 26056 12436 26108 12442
rect 26804 12434 26832 25366
rect 26896 24274 26924 31606
rect 27172 31498 27200 34954
rect 27252 34196 27304 34202
rect 27252 34138 27304 34144
rect 27264 33522 27292 34138
rect 27252 33516 27304 33522
rect 27252 33458 27304 33464
rect 27252 31748 27304 31754
rect 27252 31690 27304 31696
rect 26988 31470 27200 31498
rect 26884 24268 26936 24274
rect 26884 24210 26936 24216
rect 26884 24064 26936 24070
rect 26884 24006 26936 24012
rect 26896 23798 26924 24006
rect 26884 23792 26936 23798
rect 26884 23734 26936 23740
rect 26988 23594 27016 31470
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 27172 30938 27200 31282
rect 27160 30932 27212 30938
rect 27160 30874 27212 30880
rect 27172 29646 27200 30874
rect 27160 29640 27212 29646
rect 27160 29582 27212 29588
rect 27264 29492 27292 31690
rect 27356 29510 27384 36518
rect 27436 36304 27488 36310
rect 27436 36246 27488 36252
rect 27448 36009 27476 36246
rect 27434 36000 27490 36009
rect 27434 35935 27490 35944
rect 27618 35864 27674 35873
rect 27618 35799 27620 35808
rect 27672 35799 27674 35808
rect 27620 35770 27672 35776
rect 27712 35760 27764 35766
rect 27710 35728 27712 35737
rect 27764 35728 27766 35737
rect 27710 35663 27766 35672
rect 27436 35556 27488 35562
rect 27436 35498 27488 35504
rect 27448 35154 27476 35498
rect 27816 35442 27844 36654
rect 28078 36136 28134 36145
rect 28078 36071 28080 36080
rect 28132 36071 28134 36080
rect 28080 36042 28132 36048
rect 27988 35760 28040 35766
rect 27988 35702 28040 35708
rect 27724 35414 27844 35442
rect 27896 35488 27948 35494
rect 27896 35430 27948 35436
rect 27436 35148 27488 35154
rect 27436 35090 27488 35096
rect 27526 35048 27582 35057
rect 27526 34983 27528 34992
rect 27580 34983 27582 34992
rect 27528 34954 27580 34960
rect 27436 34536 27488 34542
rect 27436 34478 27488 34484
rect 27448 34066 27476 34478
rect 27528 34400 27580 34406
rect 27528 34342 27580 34348
rect 27540 34241 27568 34342
rect 27526 34232 27582 34241
rect 27526 34167 27582 34176
rect 27436 34060 27488 34066
rect 27436 34002 27488 34008
rect 27436 33108 27488 33114
rect 27436 33050 27488 33056
rect 27172 29464 27292 29492
rect 27344 29504 27396 29510
rect 27172 27826 27200 29464
rect 27344 29446 27396 29452
rect 27252 28484 27304 28490
rect 27252 28426 27304 28432
rect 27264 28014 27292 28426
rect 27344 28144 27396 28150
rect 27344 28086 27396 28092
rect 27252 28008 27304 28014
rect 27252 27950 27304 27956
rect 27172 27798 27292 27826
rect 27264 27033 27292 27798
rect 27356 27606 27384 28086
rect 27344 27600 27396 27606
rect 27344 27542 27396 27548
rect 27448 27470 27476 33050
rect 27540 32366 27568 34167
rect 27724 33561 27752 35414
rect 27802 35320 27858 35329
rect 27802 35255 27858 35264
rect 27816 34610 27844 35255
rect 27908 35018 27936 35430
rect 28000 35193 28028 35702
rect 28172 35624 28224 35630
rect 28170 35592 28172 35601
rect 28264 35624 28316 35630
rect 28224 35592 28226 35601
rect 28264 35566 28316 35572
rect 28170 35527 28226 35536
rect 28276 35476 28304 35566
rect 28184 35448 28304 35476
rect 28080 35216 28132 35222
rect 27986 35184 28042 35193
rect 28080 35158 28132 35164
rect 27986 35119 28042 35128
rect 27986 35048 28042 35057
rect 27896 35012 27948 35018
rect 27986 34983 27988 34992
rect 27896 34954 27948 34960
rect 28040 34983 28042 34992
rect 27988 34954 28040 34960
rect 28092 34678 28120 35158
rect 28184 35154 28212 35448
rect 28368 35222 28396 39200
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 28552 36281 28580 37198
rect 28908 37188 28960 37194
rect 28908 37130 28960 37136
rect 28632 37120 28684 37126
rect 28632 37062 28684 37068
rect 28644 36582 28672 37062
rect 28632 36576 28684 36582
rect 28632 36518 28684 36524
rect 28538 36272 28594 36281
rect 28538 36207 28594 36216
rect 28356 35216 28408 35222
rect 28356 35158 28408 35164
rect 28172 35148 28224 35154
rect 28172 35090 28224 35096
rect 28080 34672 28132 34678
rect 28080 34614 28132 34620
rect 27804 34604 27856 34610
rect 27804 34546 27856 34552
rect 28184 34134 28212 35090
rect 28920 35086 28948 37130
rect 29000 36712 29052 36718
rect 28998 36680 29000 36689
rect 29092 36712 29144 36718
rect 29052 36680 29054 36689
rect 29092 36654 29144 36660
rect 28998 36615 29054 36624
rect 29000 36100 29052 36106
rect 29000 36042 29052 36048
rect 28908 35080 28960 35086
rect 28908 35022 28960 35028
rect 29012 35034 29040 36042
rect 29104 35494 29132 36654
rect 29092 35488 29144 35494
rect 29656 35476 29684 39200
rect 30944 37330 30972 39200
rect 30380 37324 30432 37330
rect 30380 37266 30432 37272
rect 30932 37324 30984 37330
rect 30932 37266 30984 37272
rect 30288 36848 30340 36854
rect 30288 36790 30340 36796
rect 30300 36700 30328 36790
rect 30392 36718 30420 37266
rect 30472 37188 30524 37194
rect 30472 37130 30524 37136
rect 30380 36712 30432 36718
rect 30300 36672 30380 36700
rect 30380 36654 30432 36660
rect 30380 36032 30432 36038
rect 30380 35974 30432 35980
rect 29828 35760 29880 35766
rect 29828 35702 29880 35708
rect 29736 35488 29788 35494
rect 29656 35448 29736 35476
rect 29092 35430 29144 35436
rect 29736 35430 29788 35436
rect 29012 35006 29132 35034
rect 28540 34944 28592 34950
rect 28540 34886 28592 34892
rect 29000 34944 29052 34950
rect 29000 34886 29052 34892
rect 28552 34746 28580 34886
rect 28540 34740 28592 34746
rect 28540 34682 28592 34688
rect 28448 34604 28500 34610
rect 28448 34546 28500 34552
rect 28172 34128 28224 34134
rect 28172 34070 28224 34076
rect 27804 33924 27856 33930
rect 27804 33866 27856 33872
rect 27710 33552 27766 33561
rect 27710 33487 27766 33496
rect 27620 33312 27672 33318
rect 27620 33254 27672 33260
rect 27632 32774 27660 33254
rect 27620 32768 27672 32774
rect 27620 32710 27672 32716
rect 27816 32570 27844 33866
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 27896 33448 27948 33454
rect 27896 33390 27948 33396
rect 27804 32564 27856 32570
rect 27804 32506 27856 32512
rect 27620 32428 27672 32434
rect 27620 32370 27672 32376
rect 27528 32360 27580 32366
rect 27528 32302 27580 32308
rect 27632 32042 27660 32370
rect 27540 32014 27660 32042
rect 27540 30394 27568 32014
rect 27620 31952 27672 31958
rect 27620 31894 27672 31900
rect 27632 31414 27660 31894
rect 27908 31482 27936 33390
rect 27896 31476 27948 31482
rect 27896 31418 27948 31424
rect 27620 31408 27672 31414
rect 27620 31350 27672 31356
rect 27804 31204 27856 31210
rect 27804 31146 27856 31152
rect 27712 30592 27764 30598
rect 27712 30534 27764 30540
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27724 29578 27752 30534
rect 27816 30190 27844 31146
rect 27896 30592 27948 30598
rect 27896 30534 27948 30540
rect 27804 30184 27856 30190
rect 27804 30126 27856 30132
rect 27712 29572 27764 29578
rect 27712 29514 27764 29520
rect 27804 29504 27856 29510
rect 27724 29452 27804 29458
rect 27724 29446 27856 29452
rect 27724 29430 27844 29446
rect 27724 28642 27752 29430
rect 27804 28960 27856 28966
rect 27804 28902 27856 28908
rect 27816 28694 27844 28902
rect 27632 28626 27752 28642
rect 27804 28688 27856 28694
rect 27804 28630 27856 28636
rect 27620 28620 27752 28626
rect 27672 28614 27752 28620
rect 27620 28562 27672 28568
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27344 27328 27396 27334
rect 27344 27270 27396 27276
rect 27356 27062 27384 27270
rect 27344 27056 27396 27062
rect 27250 27024 27306 27033
rect 27344 26998 27396 27004
rect 27250 26959 27306 26968
rect 27068 25288 27120 25294
rect 27068 25230 27120 25236
rect 26976 23588 27028 23594
rect 26976 23530 27028 23536
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 26884 22160 26936 22166
rect 26884 22102 26936 22108
rect 26896 21962 26924 22102
rect 26988 21962 27016 23258
rect 26884 21956 26936 21962
rect 26884 21898 26936 21904
rect 26976 21956 27028 21962
rect 26976 21898 27028 21904
rect 27080 21078 27108 25230
rect 27160 25152 27212 25158
rect 27160 25094 27212 25100
rect 27172 24818 27200 25094
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27172 24342 27200 24550
rect 27160 24336 27212 24342
rect 27160 24278 27212 24284
rect 27264 23322 27292 26959
rect 27252 23316 27304 23322
rect 27252 23258 27304 23264
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27068 21072 27120 21078
rect 27068 21014 27120 21020
rect 26976 21004 27028 21010
rect 26976 20946 27028 20952
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26896 14006 26924 14826
rect 26884 14000 26936 14006
rect 26884 13942 26936 13948
rect 26056 12378 26108 12384
rect 26252 12406 26832 12434
rect 26988 12434 27016 20946
rect 27356 20466 27384 22578
rect 27448 22094 27476 27406
rect 27528 26784 27580 26790
rect 27528 26726 27580 26732
rect 27540 25974 27568 26726
rect 27528 25968 27580 25974
rect 27528 25910 27580 25916
rect 27448 22066 27568 22094
rect 27436 22024 27488 22030
rect 27436 21966 27488 21972
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27356 19718 27384 20402
rect 27448 19854 27476 21966
rect 27436 19848 27488 19854
rect 27436 19790 27488 19796
rect 27344 19712 27396 19718
rect 27344 19654 27396 19660
rect 27448 19514 27476 19790
rect 27436 19508 27488 19514
rect 27436 19450 27488 19456
rect 26988 12406 27108 12434
rect 26252 11830 26280 12406
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 25872 11756 25924 11762
rect 25872 11698 25924 11704
rect 25884 11626 25912 11698
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26976 11688 27028 11694
rect 26976 11630 27028 11636
rect 25872 11620 25924 11626
rect 25872 11562 25924 11568
rect 26068 11354 26096 11630
rect 26056 11348 26108 11354
rect 26056 11290 26108 11296
rect 26344 9178 26372 11630
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26528 11150 26556 11494
rect 26988 11218 27016 11630
rect 26976 11212 27028 11218
rect 26976 11154 27028 11160
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 20628 2508 20680 2514
rect 20628 2450 20680 2456
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 25240 2446 25268 2790
rect 25976 2446 26004 7686
rect 26344 2650 26372 8910
rect 27080 8498 27108 12406
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27356 11354 27384 11630
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 27540 6914 27568 22066
rect 27724 14958 27752 28614
rect 27908 28422 27936 30534
rect 28000 30138 28028 33798
rect 28080 33380 28132 33386
rect 28080 33322 28132 33328
rect 28092 31754 28120 33322
rect 28356 32836 28408 32842
rect 28356 32778 28408 32784
rect 28368 31890 28396 32778
rect 28356 31884 28408 31890
rect 28356 31826 28408 31832
rect 28460 31770 28488 34546
rect 29012 34066 29040 34886
rect 29104 34202 29132 35006
rect 29276 34944 29328 34950
rect 29276 34886 29328 34892
rect 29092 34196 29144 34202
rect 29092 34138 29144 34144
rect 29184 34128 29236 34134
rect 29184 34070 29236 34076
rect 29000 34060 29052 34066
rect 29000 34002 29052 34008
rect 28540 33992 28592 33998
rect 28540 33934 28592 33940
rect 28552 32230 28580 33934
rect 29000 33584 29052 33590
rect 29000 33526 29052 33532
rect 28906 33144 28962 33153
rect 28906 33079 28962 33088
rect 28540 32224 28592 32230
rect 28540 32166 28592 32172
rect 28920 31890 28948 33079
rect 29012 32570 29040 33526
rect 29196 33454 29224 34070
rect 29184 33448 29236 33454
rect 29184 33390 29236 33396
rect 29000 32564 29052 32570
rect 29000 32506 29052 32512
rect 28908 31884 28960 31890
rect 28908 31826 28960 31832
rect 28080 31748 28132 31754
rect 28080 31690 28132 31696
rect 28368 31742 28488 31770
rect 28262 31512 28318 31521
rect 28262 31447 28318 31456
rect 28000 30110 28120 30138
rect 27988 30048 28040 30054
rect 27988 29990 28040 29996
rect 28000 29306 28028 29990
rect 27988 29300 28040 29306
rect 27988 29242 28040 29248
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 27896 28416 27948 28422
rect 27896 28358 27948 28364
rect 28000 27334 28028 29106
rect 28092 27878 28120 30110
rect 28172 28960 28224 28966
rect 28172 28902 28224 28908
rect 28184 28762 28212 28902
rect 28172 28756 28224 28762
rect 28172 28698 28224 28704
rect 28276 28150 28304 31447
rect 28368 28694 28396 31742
rect 29092 31340 29144 31346
rect 29092 31282 29144 31288
rect 28448 31272 28500 31278
rect 28448 31214 28500 31220
rect 28460 30258 28488 31214
rect 28632 30592 28684 30598
rect 28632 30534 28684 30540
rect 28448 30252 28500 30258
rect 28448 30194 28500 30200
rect 28644 29714 28672 30534
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 28736 29889 28764 30194
rect 29104 30054 29132 31282
rect 29184 31136 29236 31142
rect 29184 31078 29236 31084
rect 29196 30802 29224 31078
rect 29184 30796 29236 30802
rect 29184 30738 29236 30744
rect 29092 30048 29144 30054
rect 29092 29990 29144 29996
rect 28722 29880 28778 29889
rect 28722 29815 28778 29824
rect 28632 29708 28684 29714
rect 28632 29650 28684 29656
rect 28538 29200 28594 29209
rect 28538 29135 28594 29144
rect 28356 28688 28408 28694
rect 28356 28630 28408 28636
rect 28264 28144 28316 28150
rect 28264 28086 28316 28092
rect 28080 27872 28132 27878
rect 28080 27814 28132 27820
rect 27988 27328 28040 27334
rect 27908 27288 27988 27316
rect 27908 26926 27936 27288
rect 27988 27270 28040 27276
rect 27896 26920 27948 26926
rect 27896 26862 27948 26868
rect 28172 26920 28224 26926
rect 28172 26862 28224 26868
rect 27804 25492 27856 25498
rect 27804 25434 27856 25440
rect 27816 21418 27844 25434
rect 27896 24948 27948 24954
rect 27896 24890 27948 24896
rect 27804 21412 27856 21418
rect 27804 21354 27856 21360
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27712 14952 27764 14958
rect 27712 14894 27764 14900
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27632 14006 27660 14214
rect 27724 14006 27752 14758
rect 27620 14000 27672 14006
rect 27620 13942 27672 13948
rect 27712 14000 27764 14006
rect 27712 13942 27764 13948
rect 27712 13864 27764 13870
rect 27712 13806 27764 13812
rect 27724 11762 27752 13806
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27448 6886 27568 6914
rect 27448 2650 27476 6886
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 27436 2644 27488 2650
rect 27436 2586 27488 2592
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 15016 2032 15068 2038
rect 15016 1974 15068 1980
rect 16132 800 16160 2246
rect 17420 800 17448 2246
rect 18064 800 18092 2382
rect 19352 800 19380 2382
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20640 800 20668 2246
rect 21928 800 21956 2382
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22572 800 22600 2246
rect 23860 800 23888 2382
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 25148 800 25176 2246
rect 25792 800 25820 2246
rect 27080 800 27108 2382
rect 27816 2378 27844 19654
rect 27908 15570 27936 24890
rect 28184 22098 28212 26862
rect 28276 25498 28304 28086
rect 28368 27538 28396 28630
rect 28552 28558 28580 29135
rect 29000 29096 29052 29102
rect 29000 29038 29052 29044
rect 28540 28552 28592 28558
rect 28540 28494 28592 28500
rect 28448 27872 28500 27878
rect 28448 27814 28500 27820
rect 28356 27532 28408 27538
rect 28356 27474 28408 27480
rect 28356 27396 28408 27402
rect 28356 27338 28408 27344
rect 28264 25492 28316 25498
rect 28264 25434 28316 25440
rect 28368 25294 28396 27338
rect 28356 25288 28408 25294
rect 28276 25248 28356 25276
rect 28172 22092 28224 22098
rect 28172 22034 28224 22040
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 28000 21622 28028 21830
rect 27988 21616 28040 21622
rect 27988 21558 28040 21564
rect 28080 21480 28132 21486
rect 28080 21422 28132 21428
rect 28092 19378 28120 21422
rect 28276 20058 28304 25248
rect 28356 25230 28408 25236
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 28368 20874 28396 24550
rect 28460 22778 28488 27814
rect 28552 27470 28580 28494
rect 29012 28218 29040 29038
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 29288 28150 29316 34886
rect 29840 34746 29868 35702
rect 30012 35556 30064 35562
rect 30012 35498 30064 35504
rect 29920 35284 29972 35290
rect 29920 35226 29972 35232
rect 29932 35086 29960 35226
rect 30024 35222 30052 35498
rect 30012 35216 30064 35222
rect 30012 35158 30064 35164
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 30012 35080 30064 35086
rect 30012 35022 30064 35028
rect 29828 34740 29880 34746
rect 29828 34682 29880 34688
rect 30024 34542 30052 35022
rect 30392 34746 30420 35974
rect 30484 35290 30512 37130
rect 32232 36922 32260 39200
rect 32588 37256 32640 37262
rect 32588 37198 32640 37204
rect 32220 36916 32272 36922
rect 32220 36858 32272 36864
rect 32496 36576 32548 36582
rect 32496 36518 32548 36524
rect 31852 36168 31904 36174
rect 31852 36110 31904 36116
rect 32312 36168 32364 36174
rect 32312 36110 32364 36116
rect 30840 36100 30892 36106
rect 30840 36042 30892 36048
rect 31024 36100 31076 36106
rect 31024 36042 31076 36048
rect 30852 35834 30880 36042
rect 30840 35828 30892 35834
rect 30840 35770 30892 35776
rect 30562 35728 30618 35737
rect 30562 35663 30564 35672
rect 30616 35663 30618 35672
rect 30564 35634 30616 35640
rect 30472 35284 30524 35290
rect 30472 35226 30524 35232
rect 31036 35018 31064 36042
rect 31864 35562 31892 36110
rect 31852 35556 31904 35562
rect 31852 35498 31904 35504
rect 32036 35488 32088 35494
rect 32036 35430 32088 35436
rect 31024 35012 31076 35018
rect 31024 34954 31076 34960
rect 30380 34740 30432 34746
rect 30380 34682 30432 34688
rect 30012 34536 30064 34542
rect 30012 34478 30064 34484
rect 29736 33856 29788 33862
rect 29736 33798 29788 33804
rect 29828 33856 29880 33862
rect 29828 33798 29880 33804
rect 29748 33658 29776 33798
rect 29736 33652 29788 33658
rect 29736 33594 29788 33600
rect 29840 32842 29868 33798
rect 29828 32836 29880 32842
rect 29828 32778 29880 32784
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 30104 31136 30156 31142
rect 30104 31078 30156 31084
rect 30116 30870 30144 31078
rect 30392 30870 30420 31758
rect 31760 31340 31812 31346
rect 31760 31282 31812 31288
rect 30104 30864 30156 30870
rect 30104 30806 30156 30812
rect 30380 30864 30432 30870
rect 30380 30806 30432 30812
rect 29828 30660 29880 30666
rect 29828 30602 29880 30608
rect 29920 30660 29972 30666
rect 29920 30602 29972 30608
rect 29644 28552 29696 28558
rect 29644 28494 29696 28500
rect 29276 28144 29328 28150
rect 29276 28086 29328 28092
rect 29184 28076 29236 28082
rect 29184 28018 29236 28024
rect 29196 27606 29224 28018
rect 29184 27600 29236 27606
rect 29184 27542 29236 27548
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 29184 26988 29236 26994
rect 29184 26930 29236 26936
rect 29196 26586 29224 26930
rect 29184 26580 29236 26586
rect 29184 26522 29236 26528
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 28724 26376 28776 26382
rect 28724 26318 28776 26324
rect 29092 26376 29144 26382
rect 29092 26318 29144 26324
rect 28552 26042 28580 26318
rect 28540 26036 28592 26042
rect 28540 25978 28592 25984
rect 28736 25498 28764 26318
rect 28724 25492 28776 25498
rect 28724 25434 28776 25440
rect 29104 25362 29132 26318
rect 29092 25356 29144 25362
rect 29092 25298 29144 25304
rect 29288 24750 29316 28086
rect 29276 24744 29328 24750
rect 29276 24686 29328 24692
rect 29092 24608 29144 24614
rect 29092 24550 29144 24556
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 28356 20868 28408 20874
rect 28356 20810 28408 20816
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 28460 19854 28488 21966
rect 28908 20868 28960 20874
rect 28908 20810 28960 20816
rect 28920 19990 28948 20810
rect 29012 20466 29040 23802
rect 29104 23662 29132 24550
rect 29092 23656 29144 23662
rect 29092 23598 29144 23604
rect 29552 21004 29604 21010
rect 29552 20946 29604 20952
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29564 20398 29592 20946
rect 29552 20392 29604 20398
rect 29552 20334 29604 20340
rect 28908 19984 28960 19990
rect 28828 19944 28908 19972
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28080 19372 28132 19378
rect 28080 19314 28132 19320
rect 28828 19242 28856 19944
rect 28908 19926 28960 19932
rect 29656 19786 29684 28494
rect 29840 23322 29868 30602
rect 29932 30326 29960 30602
rect 29920 30320 29972 30326
rect 29920 30262 29972 30268
rect 31484 28960 31536 28966
rect 31484 28902 31536 28908
rect 31496 28558 31524 28902
rect 31484 28552 31536 28558
rect 31484 28494 31536 28500
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 31576 27464 31628 27470
rect 31576 27406 31628 27412
rect 30392 26586 30420 27406
rect 30472 27328 30524 27334
rect 30472 27270 30524 27276
rect 30484 26858 30512 27270
rect 31588 27130 31616 27406
rect 31576 27124 31628 27130
rect 31576 27066 31628 27072
rect 30472 26852 30524 26858
rect 30472 26794 30524 26800
rect 30380 26580 30432 26586
rect 30380 26522 30432 26528
rect 29920 25832 29972 25838
rect 29920 25774 29972 25780
rect 30840 25832 30892 25838
rect 30840 25774 30892 25780
rect 29932 25362 29960 25774
rect 30288 25696 30340 25702
rect 30288 25638 30340 25644
rect 29920 25356 29972 25362
rect 29920 25298 29972 25304
rect 29828 23316 29880 23322
rect 29828 23258 29880 23264
rect 30300 23050 30328 25638
rect 30852 23254 30880 25774
rect 31772 25294 31800 31282
rect 32048 30598 32076 35430
rect 32324 35290 32352 36110
rect 32312 35284 32364 35290
rect 32312 35226 32364 35232
rect 32128 31884 32180 31890
rect 32128 31826 32180 31832
rect 32036 30592 32088 30598
rect 32036 30534 32088 30540
rect 31760 25288 31812 25294
rect 31760 25230 31812 25236
rect 31576 25152 31628 25158
rect 31576 25094 31628 25100
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 30840 23248 30892 23254
rect 30840 23190 30892 23196
rect 30288 23044 30340 23050
rect 30288 22986 30340 22992
rect 30852 22642 30880 23190
rect 31128 23186 31156 23598
rect 31116 23180 31168 23186
rect 31116 23122 31168 23128
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 29828 21888 29880 21894
rect 29828 21830 29880 21836
rect 29840 21690 29868 21830
rect 29828 21684 29880 21690
rect 29828 21626 29880 21632
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29748 20942 29776 21286
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 30472 20800 30524 20806
rect 30472 20742 30524 20748
rect 30484 20602 30512 20742
rect 30472 20596 30524 20602
rect 30472 20538 30524 20544
rect 30380 20392 30432 20398
rect 30380 20334 30432 20340
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29644 19780 29696 19786
rect 29644 19722 29696 19728
rect 29000 19712 29052 19718
rect 29000 19654 29052 19660
rect 29012 19446 29040 19654
rect 29000 19440 29052 19446
rect 29000 19382 29052 19388
rect 28908 19304 28960 19310
rect 28908 19246 28960 19252
rect 28816 19236 28868 19242
rect 28816 19178 28868 19184
rect 28920 17338 28948 19246
rect 28908 17332 28960 17338
rect 28908 17274 28960 17280
rect 27896 15564 27948 15570
rect 27896 15506 27948 15512
rect 27908 12434 27936 15506
rect 27988 14952 28040 14958
rect 27988 14894 28040 14900
rect 28000 13870 28028 14894
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 27908 12406 28120 12434
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 28000 3398 28028 11086
rect 28092 11082 28120 12406
rect 28448 12232 28500 12238
rect 28448 12174 28500 12180
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 28460 2990 28488 12174
rect 28908 8356 28960 8362
rect 28908 8298 28960 8304
rect 28920 7886 28948 8298
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 28448 2984 28500 2990
rect 28448 2926 28500 2932
rect 29748 2446 29776 20198
rect 30392 19514 30420 20334
rect 30564 19712 30616 19718
rect 30564 19654 30616 19660
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30104 19168 30156 19174
rect 30104 19110 30156 19116
rect 30116 18970 30144 19110
rect 30104 18964 30156 18970
rect 30104 18906 30156 18912
rect 29828 15428 29880 15434
rect 29828 15370 29880 15376
rect 29840 14482 29868 15370
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 30392 13530 30420 19450
rect 30576 19446 30604 19654
rect 30564 19440 30616 19446
rect 30564 19382 30616 19388
rect 30472 19304 30524 19310
rect 30472 19246 30524 19252
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30484 13394 30512 19246
rect 30564 13524 30616 13530
rect 30564 13466 30616 13472
rect 30576 13394 30604 13466
rect 30472 13388 30524 13394
rect 30472 13330 30524 13336
rect 30564 13388 30616 13394
rect 30564 13330 30616 13336
rect 30484 12434 30512 13330
rect 30392 12406 30512 12434
rect 30392 9654 30420 12406
rect 30380 9648 30432 9654
rect 30380 9590 30432 9596
rect 30472 5024 30524 5030
rect 30472 4966 30524 4972
rect 30484 2446 30512 4966
rect 31588 2582 31616 25094
rect 32140 23050 32168 31826
rect 32508 24410 32536 36518
rect 32600 31346 32628 37198
rect 32876 37108 32904 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 33140 37120 33192 37126
rect 32876 37080 33140 37108
rect 33140 37062 33192 37068
rect 33048 36780 33100 36786
rect 33048 36722 33100 36728
rect 32680 36644 32732 36650
rect 32680 36586 32732 36592
rect 32588 31340 32640 31346
rect 32588 31282 32640 31288
rect 32692 31142 32720 36586
rect 33060 36378 33088 36722
rect 33048 36372 33100 36378
rect 33048 36314 33100 36320
rect 33048 33992 33100 33998
rect 33048 33934 33100 33940
rect 33060 32570 33088 33934
rect 33048 32564 33100 32570
rect 33048 32506 33100 32512
rect 32680 31136 32732 31142
rect 32680 31078 32732 31084
rect 33048 28416 33100 28422
rect 33048 28358 33100 28364
rect 33060 27470 33088 28358
rect 33048 27464 33100 27470
rect 33048 27406 33100 27412
rect 32496 24404 32548 24410
rect 32496 24346 32548 24352
rect 32128 23044 32180 23050
rect 32128 22986 32180 22992
rect 31852 11620 31904 11626
rect 31852 11562 31904 11568
rect 31864 11150 31892 11562
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 31668 7744 31720 7750
rect 31668 7686 31720 7692
rect 31576 2576 31628 2582
rect 31576 2518 31628 2524
rect 31680 2446 31708 7686
rect 32140 4622 32168 22986
rect 33324 15904 33376 15910
rect 33324 15846 33376 15852
rect 32588 11076 32640 11082
rect 32588 11018 32640 11024
rect 32600 8974 32628 11018
rect 33140 11008 33192 11014
rect 33140 10950 33192 10956
rect 32588 8968 32640 8974
rect 32588 8910 32640 8916
rect 33152 7886 33180 10950
rect 33140 7880 33192 7886
rect 33140 7822 33192 7828
rect 32128 4616 32180 4622
rect 32128 4558 32180 4564
rect 33336 2446 33364 15846
rect 33612 14890 33640 37198
rect 34440 37108 34468 39222
rect 35438 39200 35494 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 34520 37120 34572 37126
rect 34440 37080 34520 37108
rect 34520 37062 34572 37068
rect 34520 36032 34572 36038
rect 34520 35974 34572 35980
rect 34532 30258 34560 35974
rect 34520 30252 34572 30258
rect 34520 30194 34572 30200
rect 34808 15638 34836 37198
rect 35452 36786 35480 39200
rect 36096 37262 36124 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 36084 37256 36136 37262
rect 36084 37198 36136 37204
rect 36360 37120 36412 37126
rect 36360 37062 36412 37068
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 36372 26450 36400 37062
rect 36728 36576 36780 36582
rect 36728 36518 36780 36524
rect 36740 34610 36768 36518
rect 37200 36378 37228 38791
rect 37384 37262 37412 39200
rect 38106 37496 38162 37505
rect 38106 37431 38162 37440
rect 37372 37256 37424 37262
rect 37372 37198 37424 37204
rect 37648 37120 37700 37126
rect 37648 37062 37700 37068
rect 37280 36576 37332 36582
rect 37280 36518 37332 36524
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 36728 34604 36780 34610
rect 36728 34546 36780 34552
rect 36636 29640 36688 29646
rect 36636 29582 36688 29588
rect 36648 27606 36676 29582
rect 37292 28626 37320 36518
rect 37372 36168 37424 36174
rect 37372 36110 37424 36116
rect 37384 30870 37412 36110
rect 37464 35624 37516 35630
rect 37464 35566 37516 35572
rect 37476 35465 37504 35566
rect 37462 35456 37518 35465
rect 37462 35391 37518 35400
rect 37372 30864 37424 30870
rect 37372 30806 37424 30812
rect 37464 30728 37516 30734
rect 37462 30696 37464 30705
rect 37516 30696 37518 30705
rect 37462 30631 37518 30640
rect 37280 28620 37332 28626
rect 37280 28562 37332 28568
rect 36636 27600 36688 27606
rect 36636 27542 36688 27548
rect 37464 27396 37516 27402
rect 37464 27338 37516 27344
rect 36360 26444 36412 26450
rect 36360 26386 36412 26392
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 36084 23112 36136 23118
rect 36084 23054 36136 23060
rect 36096 22778 36124 23054
rect 36084 22772 36136 22778
rect 36084 22714 36136 22720
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 36636 22024 36688 22030
rect 36636 21966 36688 21972
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 36648 18426 36676 21966
rect 36636 18420 36688 18426
rect 36636 18362 36688 18368
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 37280 17604 37332 17610
rect 37280 17546 37332 17552
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 36544 16040 36596 16046
rect 36544 15982 36596 15988
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 15632 34848 15638
rect 34796 15574 34848 15580
rect 33600 14884 33652 14890
rect 33600 14826 33652 14832
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 36556 14618 36584 15982
rect 36544 14612 36596 14618
rect 36544 14554 36596 14560
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 37292 13326 37320 17546
rect 37280 13320 37332 13326
rect 37280 13262 37332 13268
rect 37372 13184 37424 13190
rect 37372 13126 37424 13132
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 37384 12238 37412 13126
rect 37372 12232 37424 12238
rect 37372 12174 37424 12180
rect 34428 11552 34480 11558
rect 34428 11494 34480 11500
rect 34244 9580 34296 9586
rect 34244 9522 34296 9528
rect 34152 8832 34204 8838
rect 34152 8774 34204 8780
rect 34164 7886 34192 8774
rect 34152 7880 34204 7886
rect 34152 7822 34204 7828
rect 34256 3194 34284 9522
rect 34336 9512 34388 9518
rect 34334 9480 34336 9489
rect 34388 9480 34390 9489
rect 34334 9415 34390 9424
rect 34440 7410 34468 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 37476 11286 37504 27338
rect 37660 26234 37688 37062
rect 38120 36854 38148 37431
rect 38108 36848 38160 36854
rect 38108 36790 38160 36796
rect 38672 36242 38700 39200
rect 39316 36786 39344 39200
rect 39304 36780 39356 36786
rect 39304 36722 39356 36728
rect 38660 36236 38712 36242
rect 38660 36178 38712 36184
rect 38198 36136 38254 36145
rect 38198 36071 38254 36080
rect 38384 36100 38436 36106
rect 38212 36038 38240 36071
rect 38384 36042 38436 36048
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 37740 35624 37792 35630
rect 37740 35566 37792 35572
rect 37568 26206 37688 26234
rect 37568 20942 37596 26206
rect 37648 22976 37700 22982
rect 37648 22918 37700 22924
rect 37556 20936 37608 20942
rect 37556 20878 37608 20884
rect 37568 17270 37596 20878
rect 37660 19514 37688 22918
rect 37648 19508 37700 19514
rect 37648 19450 37700 19456
rect 37752 19122 37780 35566
rect 38016 34944 38068 34950
rect 38016 34886 38068 34892
rect 37832 34604 37884 34610
rect 37832 34546 37884 34552
rect 37844 34202 37872 34546
rect 37832 34196 37884 34202
rect 37832 34138 37884 34144
rect 38028 33998 38056 34886
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 38212 34105 38240 34342
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38016 33992 38068 33998
rect 38016 33934 38068 33940
rect 38108 32836 38160 32842
rect 38108 32778 38160 32784
rect 37832 32768 37884 32774
rect 38120 32745 38148 32778
rect 37832 32710 37884 32716
rect 38106 32736 38162 32745
rect 37844 26234 37872 32710
rect 38106 32671 38162 32680
rect 38292 32428 38344 32434
rect 38292 32370 38344 32376
rect 38304 32065 38332 32370
rect 38290 32056 38346 32065
rect 38290 31991 38346 32000
rect 38200 29504 38252 29510
rect 38200 29446 38252 29452
rect 38212 29345 38240 29446
rect 38198 29336 38254 29345
rect 38198 29271 38254 29280
rect 38016 28076 38068 28082
rect 38016 28018 38068 28024
rect 37924 27396 37976 27402
rect 37924 27338 37976 27344
rect 37936 26994 37964 27338
rect 37924 26988 37976 26994
rect 37924 26930 37976 26936
rect 38028 26518 38056 28018
rect 38198 27976 38254 27985
rect 38198 27911 38200 27920
rect 38252 27911 38254 27920
rect 38200 27882 38252 27888
rect 38200 27328 38252 27334
rect 38198 27296 38200 27305
rect 38252 27296 38254 27305
rect 38198 27231 38254 27240
rect 38396 27130 38424 36042
rect 38384 27124 38436 27130
rect 38384 27066 38436 27072
rect 38016 26512 38068 26518
rect 38016 26454 38068 26460
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 37844 26206 37964 26234
rect 37832 24812 37884 24818
rect 37832 24754 37884 24760
rect 37844 24410 37872 24754
rect 37832 24404 37884 24410
rect 37832 24346 37884 24352
rect 37660 19094 37780 19122
rect 37556 17264 37608 17270
rect 37556 17206 37608 17212
rect 37660 16114 37688 19094
rect 37936 18766 37964 26206
rect 38304 25945 38332 26318
rect 38290 25936 38346 25945
rect 38290 25871 38346 25880
rect 38016 24812 38068 24818
rect 38016 24754 38068 24760
rect 38028 24342 38056 24754
rect 38200 24608 38252 24614
rect 38198 24576 38200 24585
rect 38252 24576 38254 24585
rect 38198 24511 38254 24520
rect 38016 24336 38068 24342
rect 38016 24278 38068 24284
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 38304 23905 38332 24142
rect 38290 23896 38346 23905
rect 38290 23831 38346 23840
rect 38016 22976 38068 22982
rect 38016 22918 38068 22924
rect 38028 22642 38056 22918
rect 38016 22636 38068 22642
rect 38016 22578 38068 22584
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38292 21548 38344 21554
rect 38292 21490 38344 21496
rect 38304 21185 38332 21490
rect 38290 21176 38346 21185
rect 38290 21111 38346 21120
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 38304 20505 38332 20878
rect 38290 20496 38346 20505
rect 38290 20431 38346 20440
rect 38292 19372 38344 19378
rect 38292 19314 38344 19320
rect 38304 19145 38332 19314
rect 38290 19136 38346 19145
rect 38290 19071 38346 19080
rect 37924 18760 37976 18766
rect 37924 18702 37976 18708
rect 37740 17196 37792 17202
rect 37740 17138 37792 17144
rect 37752 16250 37780 17138
rect 37832 16992 37884 16998
rect 37832 16934 37884 16940
rect 37740 16244 37792 16250
rect 37740 16186 37792 16192
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 37464 11280 37516 11286
rect 37464 11222 37516 11228
rect 37188 11144 37240 11150
rect 37188 11086 37240 11092
rect 37200 10985 37228 11086
rect 37186 10976 37242 10985
rect 37186 10911 37242 10920
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 36452 10056 36504 10062
rect 36452 9998 36504 10004
rect 36464 9450 36492 9998
rect 36452 9444 36504 9450
rect 36452 9386 36504 9392
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34796 7744 34848 7750
rect 34796 7686 34848 7692
rect 34428 7404 34480 7410
rect 34428 7346 34480 7352
rect 34808 6798 34836 7686
rect 37740 7200 37792 7206
rect 37740 7142 37792 7148
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34796 6792 34848 6798
rect 34796 6734 34848 6740
rect 37464 6248 37516 6254
rect 37462 6216 37464 6225
rect 37516 6216 37518 6225
rect 37462 6151 37518 6160
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 37752 4622 37780 7142
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 35348 4480 35400 4486
rect 35348 4422 35400 4428
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34244 3188 34296 3194
rect 34244 3130 34296 3136
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 2446 35388 4422
rect 37844 3602 37872 16934
rect 37936 16590 37964 18702
rect 38292 18284 38344 18290
rect 38292 18226 38344 18232
rect 38304 17785 38332 18226
rect 38290 17776 38346 17785
rect 38290 17711 38346 17720
rect 37924 16584 37976 16590
rect 37924 16526 37976 16532
rect 38108 16516 38160 16522
rect 38108 16458 38160 16464
rect 37924 16448 37976 16454
rect 38120 16425 38148 16458
rect 38200 16448 38252 16454
rect 37924 16390 37976 16396
rect 38106 16416 38162 16425
rect 37936 4146 37964 16390
rect 38200 16390 38252 16396
rect 38106 16351 38162 16360
rect 38212 13734 38240 16390
rect 38292 16108 38344 16114
rect 38292 16050 38344 16056
rect 38304 15745 38332 16050
rect 38290 15736 38346 15745
rect 38290 15671 38346 15680
rect 38292 14408 38344 14414
rect 38290 14376 38292 14385
rect 38344 14376 38346 14385
rect 38290 14311 38346 14320
rect 38200 13728 38252 13734
rect 38200 13670 38252 13676
rect 38200 13184 38252 13190
rect 38200 13126 38252 13132
rect 38212 13025 38240 13126
rect 38198 13016 38254 13025
rect 38198 12951 38254 12960
rect 38016 12844 38068 12850
rect 38016 12786 38068 12792
rect 38028 12442 38056 12786
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38016 12436 38068 12442
rect 38016 12378 38068 12384
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38200 9920 38252 9926
rect 38200 9862 38252 9868
rect 38212 9625 38240 9862
rect 38198 9616 38254 9625
rect 38198 9551 38254 9560
rect 38108 8492 38160 8498
rect 38108 8434 38160 8440
rect 38120 8265 38148 8434
rect 38106 8256 38162 8265
rect 38106 8191 38162 8200
rect 38200 7744 38252 7750
rect 38200 7686 38252 7692
rect 38212 7585 38240 7686
rect 38198 7576 38254 7585
rect 38198 7511 38254 7520
rect 38016 6656 38068 6662
rect 38016 6598 38068 6604
rect 38028 5234 38056 6598
rect 38016 5228 38068 5234
rect 38016 5170 38068 5176
rect 38200 5024 38252 5030
rect 38200 4966 38252 4972
rect 38212 4865 38240 4966
rect 38198 4856 38254 4865
rect 38198 4791 38254 4800
rect 38200 4480 38252 4486
rect 38200 4422 38252 4428
rect 38212 4185 38240 4422
rect 38198 4176 38254 4185
rect 37924 4140 37976 4146
rect 38198 4111 38254 4120
rect 37924 4082 37976 4088
rect 39304 3936 39356 3942
rect 39304 3878 39356 3884
rect 37832 3596 37884 3602
rect 37832 3538 37884 3544
rect 37924 3528 37976 3534
rect 37924 3470 37976 3476
rect 37280 3120 37332 3126
rect 37280 3062 37332 3068
rect 36728 3052 36780 3058
rect 36728 2994 36780 3000
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 30472 2440 30524 2446
rect 30472 2382 30524 2388
rect 31668 2440 31720 2446
rect 31668 2382 31720 2388
rect 33324 2440 33376 2446
rect 33324 2382 33376 2388
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 27804 2372 27856 2378
rect 27804 2314 27856 2320
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 28368 800 28396 2314
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 29656 800 29684 2246
rect 30300 800 30328 2246
rect 31588 800 31616 2246
rect 32876 800 32904 2246
rect 33520 800 33548 2246
rect 34808 800 34836 2246
rect 36096 800 36124 2246
rect 36740 800 36768 2994
rect 37292 2514 37320 3062
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 37476 2825 37504 2926
rect 37462 2816 37518 2825
rect 37462 2751 37518 2760
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 37476 1465 37504 2382
rect 37936 1986 37964 3470
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 37936 1958 38056 1986
rect 37462 1456 37518 1465
rect 37462 1391 37518 1400
rect 38028 800 38056 1958
rect 1674 776 1730 785
rect 1674 711 1730 720
rect 1950 200 2006 800
rect 3238 200 3294 800
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 10966 200 11022 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 14186 200 14242 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 17406 200 17462 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 20626 200 20682 800
rect 21914 200 21970 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 32862 200 32918 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 36726 200 36782 800
rect 38014 200 38070 800
rect 38212 785 38240 3334
rect 39316 800 39344 3878
rect 38198 776 38254 785
rect 38198 711 38254 720
rect 39302 200 39358 800
<< via2 >>
rect 1766 38800 1822 38856
rect 2870 38120 2926 38176
rect 1398 23160 1454 23216
rect 1398 19080 1454 19136
rect 1674 35400 1730 35456
rect 1766 34720 1822 34776
rect 1766 33380 1822 33416
rect 1766 33360 1768 33380
rect 1768 33360 1820 33380
rect 1820 33360 1822 33380
rect 1766 32000 1822 32056
rect 1766 31340 1822 31376
rect 1766 31320 1768 31340
rect 1768 31320 1820 31340
rect 1820 31320 1822 31340
rect 1766 29960 1822 30016
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 3514 36760 3570 36816
rect 1766 28600 1822 28656
rect 1766 27240 1822 27296
rect 1674 26560 1730 26616
rect 1858 26424 1914 26480
rect 1766 25200 1822 25256
rect 1582 24928 1638 24984
rect 1766 23840 1822 23896
rect 2226 27648 2282 27704
rect 1766 21836 1768 21856
rect 1768 21836 1820 21856
rect 1820 21836 1822 21856
rect 1766 21800 1822 21836
rect 1766 20440 1822 20496
rect 1766 18400 1822 18456
rect 1674 17040 1730 17096
rect 1766 15680 1822 15736
rect 1766 15000 1822 15056
rect 1766 13676 1768 13696
rect 1768 13676 1820 13696
rect 1820 13676 1822 13696
rect 1766 13640 1822 13676
rect 1766 12280 1822 12336
rect 1582 7520 1638 7576
rect 2594 16632 2650 16688
rect 2226 9560 2282 9616
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 7746 36524 7748 36544
rect 7748 36524 7800 36544
rect 7800 36524 7802 36544
rect 7746 36488 7802 36524
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4066 34584 4122 34640
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 3422 26308 3478 26344
rect 3422 26288 3424 26308
rect 3424 26288 3476 26308
rect 3476 26288 3478 26308
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 2870 11600 2926 11656
rect 2778 10240 2834 10296
rect 2594 9580 2650 9616
rect 2594 9560 2596 9580
rect 2596 9560 2648 9580
rect 2648 9560 2650 9580
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 3790 21936 3846 21992
rect 2778 8880 2834 8936
rect 1674 6840 1730 6896
rect 1766 5516 1768 5536
rect 1768 5516 1820 5536
rect 1820 5516 1822 5536
rect 1766 5480 1822 5516
rect 1674 4120 1730 4176
rect 3422 14184 3478 14240
rect 3514 10920 3570 10976
rect 1766 3476 1768 3496
rect 1768 3476 1820 3496
rect 1820 3476 1822 3496
rect 1766 3440 1822 3476
rect 2502 2080 2558 2136
rect 5354 31340 5410 31376
rect 5354 31320 5356 31340
rect 5356 31320 5408 31340
rect 5408 31320 5410 31340
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4250 21428 4252 21448
rect 4252 21428 4304 21448
rect 4304 21428 4306 21448
rect 4250 21392 4306 21428
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4158 18164 4160 18184
rect 4160 18164 4212 18184
rect 4212 18164 4214 18184
rect 4158 18128 4214 18164
rect 4526 18128 4582 18184
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 3974 16088 4030 16144
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4894 12824 4950 12880
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 5262 21392 5318 21448
rect 6458 34040 6514 34096
rect 6182 32852 6184 32872
rect 6184 32852 6236 32872
rect 6236 32852 6238 32872
rect 6182 32816 6238 32852
rect 6366 25064 6422 25120
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 6826 25064 6882 25120
rect 7286 14184 7342 14240
rect 7654 15272 7710 15328
rect 9310 36760 9366 36816
rect 9494 34992 9550 35048
rect 10322 36216 10378 36272
rect 10230 35536 10286 35592
rect 11058 33904 11114 33960
rect 11334 33904 11390 33960
rect 8390 21972 8392 21992
rect 8392 21972 8444 21992
rect 8444 21972 8446 21992
rect 8390 21936 8446 21972
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8758 16108 8814 16144
rect 8758 16088 8760 16108
rect 8760 16088 8812 16108
rect 8812 16088 8814 16108
rect 9586 17176 9642 17232
rect 9678 16108 9734 16144
rect 9678 16088 9680 16108
rect 9680 16088 9732 16108
rect 9732 16088 9734 16108
rect 9862 14884 9918 14920
rect 9862 14864 9864 14884
rect 9864 14864 9916 14884
rect 9916 14864 9918 14884
rect 10046 12552 10102 12608
rect 13542 35944 13598 36000
rect 11426 32680 11482 32736
rect 10782 26152 10838 26208
rect 10414 15136 10470 15192
rect 10966 17196 11022 17232
rect 10966 17176 10968 17196
rect 10968 17176 11020 17196
rect 11020 17176 11022 17196
rect 10506 12552 10562 12608
rect 11610 26152 11666 26208
rect 13358 35148 13414 35184
rect 13358 35128 13360 35148
rect 13360 35128 13412 35148
rect 13412 35128 13414 35148
rect 13726 32000 13782 32056
rect 14646 36100 14702 36136
rect 14646 36080 14648 36100
rect 14648 36080 14700 36100
rect 14700 36080 14702 36100
rect 14186 34176 14242 34232
rect 14830 34584 14886 34640
rect 16578 35264 16634 35320
rect 16026 34312 16082 34368
rect 13726 27004 13728 27024
rect 13728 27004 13780 27024
rect 13780 27004 13782 27024
rect 13726 26968 13782 27004
rect 17406 36624 17462 36680
rect 16946 36352 17002 36408
rect 16946 35400 17002 35456
rect 16946 34892 16948 34912
rect 16948 34892 17000 34912
rect 17000 34892 17002 34912
rect 16946 34856 17002 34892
rect 16302 29824 16358 29880
rect 15842 28328 15898 28384
rect 15750 28056 15806 28112
rect 15382 26696 15438 26752
rect 14646 13368 14702 13424
rect 13358 12144 13414 12200
rect 16762 30252 16818 30288
rect 18326 36352 18382 36408
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 20534 36896 20590 36952
rect 19246 36352 19302 36408
rect 18694 35980 18696 36000
rect 18696 35980 18748 36000
rect 18748 35980 18750 36000
rect 18694 35944 18750 35980
rect 18510 35672 18566 35728
rect 17958 34856 18014 34912
rect 18142 34312 18198 34368
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 20074 35808 20130 35864
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19246 33088 19302 33144
rect 17682 31184 17738 31240
rect 16762 30232 16764 30252
rect 16764 30232 16816 30252
rect 16816 30232 16818 30252
rect 16946 30116 17002 30152
rect 16946 30096 16948 30116
rect 16948 30096 17000 30116
rect 17000 30096 17002 30116
rect 16486 27532 16542 27568
rect 16486 27512 16488 27532
rect 16488 27512 16540 27532
rect 16540 27512 16542 27532
rect 16946 26308 17002 26344
rect 16946 26288 16948 26308
rect 16948 26288 17000 26308
rect 17000 26288 17002 26308
rect 17406 26288 17462 26344
rect 17774 29844 17830 29880
rect 17774 29824 17776 29844
rect 17776 29824 17828 29844
rect 17828 29824 17830 29844
rect 18142 29688 18198 29744
rect 18326 30116 18382 30152
rect 18326 30096 18328 30116
rect 18328 30096 18380 30116
rect 18380 30096 18382 30116
rect 17866 28364 17868 28384
rect 17868 28364 17920 28384
rect 17920 28364 17922 28384
rect 17866 28328 17922 28364
rect 17866 28056 17922 28112
rect 17958 27668 18014 27704
rect 17958 27648 17960 27668
rect 17960 27648 18012 27668
rect 18012 27648 18014 27668
rect 17774 27376 17830 27432
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19430 31048 19486 31104
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19706 30096 19762 30152
rect 19338 29552 19394 29608
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19430 29144 19486 29200
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 18786 27668 18842 27704
rect 18786 27648 18788 27668
rect 18788 27648 18840 27668
rect 18840 27648 18842 27668
rect 18326 25608 18382 25664
rect 18786 26732 18788 26752
rect 18788 26732 18840 26752
rect 18840 26732 18842 26752
rect 18786 26696 18842 26732
rect 18786 26152 18842 26208
rect 16670 15020 16726 15056
rect 16670 15000 16672 15020
rect 16672 15000 16724 15020
rect 16724 15000 16726 15020
rect 15658 13504 15714 13560
rect 18050 15000 18106 15056
rect 18418 15136 18474 15192
rect 19154 25608 19210 25664
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 20350 34856 20406 34912
rect 20718 36624 20774 36680
rect 21638 36624 21694 36680
rect 22190 36644 22246 36680
rect 22190 36624 22192 36644
rect 22192 36624 22244 36644
rect 22244 36624 22246 36644
rect 20810 35400 20866 35456
rect 20994 35436 20996 35456
rect 20996 35436 21048 35456
rect 21048 35436 21050 35456
rect 20994 35400 21050 35436
rect 20994 32680 21050 32736
rect 21178 32544 21234 32600
rect 21086 32000 21142 32056
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19890 25372 19892 25392
rect 19892 25372 19944 25392
rect 19944 25372 19946 25392
rect 19890 25336 19946 25372
rect 19798 25220 19854 25256
rect 19798 25200 19800 25220
rect 19800 25200 19852 25220
rect 19852 25200 19854 25220
rect 20074 26424 20130 26480
rect 20534 30232 20590 30288
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 20166 24656 20222 24712
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19062 14864 19118 14920
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20442 25220 20498 25256
rect 20442 25200 20444 25220
rect 20444 25200 20496 25220
rect 20496 25200 20498 25220
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 20626 24112 20682 24168
rect 20626 23568 20682 23624
rect 20718 23296 20774 23352
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 21730 34856 21786 34912
rect 21546 29844 21602 29880
rect 21546 29824 21548 29844
rect 21548 29824 21600 29844
rect 21600 29824 21602 29844
rect 21362 27532 21418 27568
rect 21362 27512 21364 27532
rect 21364 27512 21416 27532
rect 21416 27512 21418 27532
rect 21546 27376 21602 27432
rect 22466 34620 22468 34640
rect 22468 34620 22520 34640
rect 22520 34620 22522 34640
rect 22466 34584 22522 34620
rect 22098 33904 22154 33960
rect 22098 33496 22154 33552
rect 22006 32952 22062 33008
rect 22282 33360 22338 33416
rect 22190 32952 22246 33008
rect 22190 31456 22246 31512
rect 24214 36896 24270 36952
rect 22466 32680 22522 32736
rect 21914 27940 21970 27976
rect 21914 27920 21916 27940
rect 21916 27920 21968 27940
rect 21968 27920 21970 27940
rect 21822 27376 21878 27432
rect 21822 19896 21878 19952
rect 22742 31728 22798 31784
rect 22650 31048 22706 31104
rect 23294 34448 23350 34504
rect 23110 34040 23166 34096
rect 23478 33904 23534 33960
rect 23294 33088 23350 33144
rect 25226 36488 25282 36544
rect 24582 35944 24638 36000
rect 23754 34484 23756 34504
rect 23756 34484 23808 34504
rect 23808 34484 23810 34504
rect 23754 34448 23810 34484
rect 23662 31184 23718 31240
rect 23386 29688 23442 29744
rect 21822 16496 21878 16552
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 22926 23604 22928 23624
rect 22928 23604 22980 23624
rect 22980 23604 22982 23624
rect 22926 23568 22982 23604
rect 23110 24148 23112 24168
rect 23112 24148 23164 24168
rect 23164 24148 23166 24168
rect 23110 24112 23166 24148
rect 23386 27512 23442 27568
rect 23754 29588 23756 29608
rect 23756 29588 23808 29608
rect 23808 29588 23810 29608
rect 23754 29552 23810 29588
rect 23846 26288 23902 26344
rect 23478 16496 23534 16552
rect 24030 17604 24086 17640
rect 24030 17584 24032 17604
rect 24032 17584 24084 17604
rect 24084 17584 24086 17604
rect 25870 36644 25926 36680
rect 25870 36624 25872 36644
rect 25872 36624 25924 36644
rect 25924 36624 25926 36644
rect 26330 36352 26386 36408
rect 24950 32816 25006 32872
rect 24766 31764 24768 31784
rect 24768 31764 24820 31784
rect 24820 31764 24822 31784
rect 24766 31728 24822 31764
rect 24858 27940 24914 27976
rect 24858 27920 24860 27940
rect 24860 27920 24912 27940
rect 24912 27920 24914 27940
rect 24950 24656 25006 24712
rect 25778 35672 25834 35728
rect 25226 31320 25282 31376
rect 25318 27412 25320 27432
rect 25320 27412 25372 27432
rect 25372 27412 25374 27432
rect 25318 27376 25374 27412
rect 24950 19896 25006 19952
rect 25594 33940 25596 33960
rect 25596 33940 25648 33960
rect 25648 33940 25650 33960
rect 25594 33904 25650 33940
rect 25502 31728 25558 31784
rect 25502 31184 25558 31240
rect 26422 35400 26478 35456
rect 26238 34992 26294 35048
rect 25962 33224 26018 33280
rect 26330 32564 26386 32600
rect 26330 32544 26332 32564
rect 26332 32544 26384 32564
rect 26384 32544 26386 32564
rect 25502 25336 25558 25392
rect 25778 26424 25834 26480
rect 28078 36760 28134 36816
rect 26790 33360 26846 33416
rect 26790 32680 26846 32736
rect 27434 35944 27490 36000
rect 27618 35828 27674 35864
rect 27618 35808 27620 35828
rect 27620 35808 27672 35828
rect 27672 35808 27674 35828
rect 27710 35708 27712 35728
rect 27712 35708 27764 35728
rect 27764 35708 27766 35728
rect 27710 35672 27766 35708
rect 28078 36100 28134 36136
rect 28078 36080 28080 36100
rect 28080 36080 28132 36100
rect 28132 36080 28134 36100
rect 27526 35012 27582 35048
rect 27526 34992 27528 35012
rect 27528 34992 27580 35012
rect 27580 34992 27582 35012
rect 27526 34176 27582 34232
rect 27802 35264 27858 35320
rect 28170 35572 28172 35592
rect 28172 35572 28224 35592
rect 28224 35572 28226 35592
rect 28170 35536 28226 35572
rect 27986 35128 28042 35184
rect 27986 35012 28042 35048
rect 27986 34992 27988 35012
rect 27988 34992 28040 35012
rect 28040 34992 28042 35012
rect 28538 36216 28594 36272
rect 28998 36660 29000 36680
rect 29000 36660 29052 36680
rect 29052 36660 29054 36680
rect 28998 36624 29054 36660
rect 27710 33496 27766 33552
rect 27250 26968 27306 27024
rect 28906 33088 28962 33144
rect 28262 31456 28318 31512
rect 28722 29824 28778 29880
rect 28538 29144 28594 29200
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 30562 35692 30618 35728
rect 30562 35672 30564 35692
rect 30564 35672 30616 35692
rect 30616 35672 30618 35692
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37186 38800 37242 38856
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 38106 37440 38162 37496
rect 37462 35400 37518 35456
rect 37462 30676 37464 30696
rect 37464 30676 37516 30696
rect 37516 30676 37518 30696
rect 37462 30640 37518 30676
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34334 9460 34336 9480
rect 34336 9460 34388 9480
rect 34388 9460 34390 9480
rect 34334 9424 34390 9460
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 38198 36080 38254 36136
rect 38198 34040 38254 34096
rect 38106 32680 38162 32736
rect 38290 32000 38346 32056
rect 38198 29280 38254 29336
rect 38198 27940 38254 27976
rect 38198 27920 38200 27940
rect 38200 27920 38252 27940
rect 38252 27920 38254 27940
rect 38198 27276 38200 27296
rect 38200 27276 38252 27296
rect 38252 27276 38254 27296
rect 38198 27240 38254 27276
rect 38290 25880 38346 25936
rect 38198 24556 38200 24576
rect 38200 24556 38252 24576
rect 38252 24556 38254 24576
rect 38198 24520 38254 24556
rect 38290 23840 38346 23896
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38290 21120 38346 21176
rect 38290 20440 38346 20496
rect 38290 19080 38346 19136
rect 37186 10920 37242 10976
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 37462 6196 37464 6216
rect 37464 6196 37516 6216
rect 37516 6196 37518 6216
rect 37462 6160 37518 6196
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38290 17720 38346 17776
rect 38106 16360 38162 16416
rect 38290 15680 38346 15736
rect 38290 14356 38292 14376
rect 38292 14356 38344 14376
rect 38344 14356 38346 14376
rect 38290 14320 38346 14356
rect 38198 12960 38254 13016
rect 38198 12280 38254 12336
rect 38198 9560 38254 9616
rect 38106 8200 38162 8256
rect 38198 7520 38254 7576
rect 38198 4800 38254 4856
rect 38198 4120 38254 4176
rect 37462 2760 37518 2816
rect 37462 1400 37518 1456
rect 1674 720 1730 776
rect 38198 720 38254 776
<< metal3 >>
rect 200 38858 800 38888
rect 1761 38858 1827 38861
rect 200 38856 1827 38858
rect 200 38800 1766 38856
rect 1822 38800 1827 38856
rect 200 38798 1827 38800
rect 200 38768 800 38798
rect 1761 38795 1827 38798
rect 37181 38858 37247 38861
rect 39200 38858 39800 38888
rect 37181 38856 39800 38858
rect 37181 38800 37186 38856
rect 37242 38800 39800 38856
rect 37181 38798 39800 38800
rect 37181 38795 37247 38798
rect 39200 38768 39800 38798
rect 200 38178 800 38208
rect 2865 38178 2931 38181
rect 200 38176 2931 38178
rect 200 38120 2870 38176
rect 2926 38120 2931 38176
rect 200 38118 2931 38120
rect 200 38088 800 38118
rect 2865 38115 2931 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 38101 37498 38167 37501
rect 39200 37498 39800 37528
rect 38101 37496 39800 37498
rect 38101 37440 38106 37496
rect 38162 37440 39800 37496
rect 38101 37438 39800 37440
rect 38101 37435 38167 37438
rect 39200 37408 39800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 20529 36954 20595 36957
rect 24209 36954 24275 36957
rect 20529 36952 24275 36954
rect 20529 36896 20534 36952
rect 20590 36896 24214 36952
rect 24270 36896 24275 36952
rect 20529 36894 24275 36896
rect 20529 36891 20595 36894
rect 24209 36891 24275 36894
rect 200 36818 800 36848
rect 3509 36818 3575 36821
rect 200 36816 3575 36818
rect 200 36760 3514 36816
rect 3570 36760 3575 36816
rect 200 36758 3575 36760
rect 200 36728 800 36758
rect 3509 36755 3575 36758
rect 9305 36818 9371 36821
rect 28073 36818 28139 36821
rect 9305 36816 28139 36818
rect 9305 36760 9310 36816
rect 9366 36760 28078 36816
rect 28134 36760 28139 36816
rect 9305 36758 28139 36760
rect 9305 36755 9371 36758
rect 28073 36755 28139 36758
rect 17401 36682 17467 36685
rect 20713 36682 20779 36685
rect 17401 36680 20779 36682
rect 17401 36624 17406 36680
rect 17462 36624 20718 36680
rect 20774 36624 20779 36680
rect 17401 36622 20779 36624
rect 17401 36619 17467 36622
rect 20713 36619 20779 36622
rect 21633 36682 21699 36685
rect 22185 36682 22251 36685
rect 21633 36680 22251 36682
rect 21633 36624 21638 36680
rect 21694 36624 22190 36680
rect 22246 36624 22251 36680
rect 21633 36622 22251 36624
rect 21633 36619 21699 36622
rect 22185 36619 22251 36622
rect 25865 36682 25931 36685
rect 28993 36682 29059 36685
rect 25865 36680 29059 36682
rect 25865 36624 25870 36680
rect 25926 36624 28998 36680
rect 29054 36624 29059 36680
rect 25865 36622 29059 36624
rect 25865 36619 25931 36622
rect 28993 36619 29059 36622
rect 7741 36546 7807 36549
rect 25221 36546 25287 36549
rect 7741 36544 25287 36546
rect 7741 36488 7746 36544
rect 7802 36488 25226 36544
rect 25282 36488 25287 36544
rect 7741 36486 25287 36488
rect 7741 36483 7807 36486
rect 25221 36483 25287 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 16941 36410 17007 36413
rect 18321 36410 18387 36413
rect 16941 36408 18387 36410
rect 16941 36352 16946 36408
rect 17002 36352 18326 36408
rect 18382 36352 18387 36408
rect 16941 36350 18387 36352
rect 16941 36347 17007 36350
rect 18321 36347 18387 36350
rect 19241 36410 19307 36413
rect 26325 36410 26391 36413
rect 19241 36408 26391 36410
rect 19241 36352 19246 36408
rect 19302 36352 26330 36408
rect 26386 36352 26391 36408
rect 19241 36350 26391 36352
rect 19241 36347 19307 36350
rect 26325 36347 26391 36350
rect 10317 36274 10383 36277
rect 28533 36274 28599 36277
rect 10317 36272 28599 36274
rect 10317 36216 10322 36272
rect 10378 36216 28538 36272
rect 28594 36216 28599 36272
rect 10317 36214 28599 36216
rect 10317 36211 10383 36214
rect 28533 36211 28599 36214
rect 14641 36138 14707 36141
rect 28073 36138 28139 36141
rect 14641 36136 28139 36138
rect 14641 36080 14646 36136
rect 14702 36080 28078 36136
rect 28134 36080 28139 36136
rect 14641 36078 28139 36080
rect 14641 36075 14707 36078
rect 28073 36075 28139 36078
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 13537 36002 13603 36005
rect 18689 36002 18755 36005
rect 13537 36000 18755 36002
rect 13537 35944 13542 36000
rect 13598 35944 18694 36000
rect 18750 35944 18755 36000
rect 13537 35942 18755 35944
rect 13537 35939 13603 35942
rect 18689 35939 18755 35942
rect 24577 36002 24643 36005
rect 27429 36002 27495 36005
rect 24577 36000 27495 36002
rect 24577 35944 24582 36000
rect 24638 35944 27434 36000
rect 27490 35944 27495 36000
rect 24577 35942 27495 35944
rect 24577 35939 24643 35942
rect 27429 35939 27495 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 20069 35866 20135 35869
rect 27613 35866 27679 35869
rect 20069 35864 27679 35866
rect 20069 35808 20074 35864
rect 20130 35808 27618 35864
rect 27674 35808 27679 35864
rect 20069 35806 27679 35808
rect 20069 35803 20135 35806
rect 27613 35803 27679 35806
rect 18505 35730 18571 35733
rect 25773 35730 25839 35733
rect 18505 35728 25839 35730
rect 18505 35672 18510 35728
rect 18566 35672 25778 35728
rect 25834 35672 25839 35728
rect 18505 35670 25839 35672
rect 18505 35667 18571 35670
rect 25773 35667 25839 35670
rect 27705 35730 27771 35733
rect 30557 35730 30623 35733
rect 27705 35728 30623 35730
rect 27705 35672 27710 35728
rect 27766 35672 30562 35728
rect 30618 35672 30623 35728
rect 27705 35670 30623 35672
rect 27705 35667 27771 35670
rect 30557 35667 30623 35670
rect 10225 35594 10291 35597
rect 28165 35594 28231 35597
rect 10225 35592 28231 35594
rect 10225 35536 10230 35592
rect 10286 35536 28170 35592
rect 28226 35536 28231 35592
rect 10225 35534 28231 35536
rect 10225 35531 10291 35534
rect 28165 35531 28231 35534
rect 200 35458 800 35488
rect 1669 35458 1735 35461
rect 200 35456 1735 35458
rect 200 35400 1674 35456
rect 1730 35400 1735 35456
rect 200 35398 1735 35400
rect 200 35368 800 35398
rect 1669 35395 1735 35398
rect 16941 35458 17007 35461
rect 20805 35458 20871 35461
rect 16941 35456 20871 35458
rect 16941 35400 16946 35456
rect 17002 35400 20810 35456
rect 20866 35400 20871 35456
rect 16941 35398 20871 35400
rect 16941 35395 17007 35398
rect 20805 35395 20871 35398
rect 20989 35458 21055 35461
rect 26417 35458 26483 35461
rect 20989 35456 26483 35458
rect 20989 35400 20994 35456
rect 21050 35400 26422 35456
rect 26478 35400 26483 35456
rect 20989 35398 26483 35400
rect 20989 35395 21055 35398
rect 26417 35395 26483 35398
rect 37457 35458 37523 35461
rect 39200 35458 39800 35488
rect 37457 35456 39800 35458
rect 37457 35400 37462 35456
rect 37518 35400 39800 35456
rect 37457 35398 39800 35400
rect 37457 35395 37523 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 16573 35322 16639 35325
rect 27797 35322 27863 35325
rect 16573 35320 27863 35322
rect 16573 35264 16578 35320
rect 16634 35264 27802 35320
rect 27858 35264 27863 35320
rect 16573 35262 27863 35264
rect 16573 35259 16639 35262
rect 27797 35259 27863 35262
rect 13353 35186 13419 35189
rect 27981 35186 28047 35189
rect 13353 35184 28047 35186
rect 13353 35128 13358 35184
rect 13414 35128 27986 35184
rect 28042 35128 28047 35184
rect 13353 35126 28047 35128
rect 13353 35123 13419 35126
rect 27981 35123 28047 35126
rect 9489 35050 9555 35053
rect 26233 35050 26299 35053
rect 9489 35048 26299 35050
rect 9489 34992 9494 35048
rect 9550 34992 26238 35048
rect 26294 34992 26299 35048
rect 9489 34990 26299 34992
rect 9489 34987 9555 34990
rect 26233 34987 26299 34990
rect 27521 35050 27587 35053
rect 27981 35050 28047 35053
rect 27521 35048 28047 35050
rect 27521 34992 27526 35048
rect 27582 34992 27986 35048
rect 28042 34992 28047 35048
rect 27521 34990 28047 34992
rect 27521 34987 27587 34990
rect 27981 34987 28047 34990
rect 16941 34914 17007 34917
rect 17953 34914 18019 34917
rect 16941 34912 18019 34914
rect 16941 34856 16946 34912
rect 17002 34856 17958 34912
rect 18014 34856 18019 34912
rect 16941 34854 18019 34856
rect 16941 34851 17007 34854
rect 17953 34851 18019 34854
rect 20345 34914 20411 34917
rect 21725 34914 21791 34917
rect 20345 34912 21791 34914
rect 20345 34856 20350 34912
rect 20406 34856 21730 34912
rect 21786 34856 21791 34912
rect 20345 34854 21791 34856
rect 20345 34851 20411 34854
rect 21725 34851 21791 34854
rect 19570 34848 19886 34849
rect 200 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 1761 34778 1827 34781
rect 200 34776 1827 34778
rect 200 34720 1766 34776
rect 1822 34720 1827 34776
rect 200 34718 1827 34720
rect 200 34688 800 34718
rect 1761 34715 1827 34718
rect 3918 34580 3924 34644
rect 3988 34642 3994 34644
rect 4061 34642 4127 34645
rect 3988 34640 4127 34642
rect 3988 34584 4066 34640
rect 4122 34584 4127 34640
rect 3988 34582 4127 34584
rect 3988 34580 3994 34582
rect 4061 34579 4127 34582
rect 14825 34642 14891 34645
rect 22461 34642 22527 34645
rect 14825 34640 22527 34642
rect 14825 34584 14830 34640
rect 14886 34584 22466 34640
rect 22522 34584 22527 34640
rect 14825 34582 22527 34584
rect 14825 34579 14891 34582
rect 22461 34579 22527 34582
rect 23289 34506 23355 34509
rect 23749 34506 23815 34509
rect 23289 34504 23815 34506
rect 23289 34448 23294 34504
rect 23350 34448 23754 34504
rect 23810 34448 23815 34504
rect 23289 34446 23815 34448
rect 23289 34443 23355 34446
rect 23749 34443 23815 34446
rect 16021 34370 16087 34373
rect 18137 34370 18203 34373
rect 16021 34368 18203 34370
rect 16021 34312 16026 34368
rect 16082 34312 18142 34368
rect 18198 34312 18203 34368
rect 16021 34310 18203 34312
rect 16021 34307 16087 34310
rect 18137 34307 18203 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 14181 34234 14247 34237
rect 27521 34234 27587 34237
rect 14181 34232 27587 34234
rect 14181 34176 14186 34232
rect 14242 34176 27526 34232
rect 27582 34176 27587 34232
rect 14181 34174 27587 34176
rect 14181 34171 14247 34174
rect 27521 34171 27587 34174
rect 6453 34098 6519 34101
rect 23105 34098 23171 34101
rect 6453 34096 23171 34098
rect 6453 34040 6458 34096
rect 6514 34040 23110 34096
rect 23166 34040 23171 34096
rect 6453 34038 23171 34040
rect 6453 34035 6519 34038
rect 23105 34035 23171 34038
rect 38193 34098 38259 34101
rect 39200 34098 39800 34128
rect 38193 34096 39800 34098
rect 38193 34040 38198 34096
rect 38254 34040 39800 34096
rect 38193 34038 39800 34040
rect 38193 34035 38259 34038
rect 39200 34008 39800 34038
rect 11053 33962 11119 33965
rect 11329 33962 11395 33965
rect 22093 33962 22159 33965
rect 11053 33960 22159 33962
rect 11053 33904 11058 33960
rect 11114 33904 11334 33960
rect 11390 33904 22098 33960
rect 22154 33904 22159 33960
rect 11053 33902 22159 33904
rect 11053 33899 11119 33902
rect 11329 33899 11395 33902
rect 22093 33899 22159 33902
rect 23473 33962 23539 33965
rect 25589 33962 25655 33965
rect 23473 33960 25655 33962
rect 23473 33904 23478 33960
rect 23534 33904 25594 33960
rect 25650 33904 25655 33960
rect 23473 33902 25655 33904
rect 23473 33899 23539 33902
rect 25589 33899 25655 33902
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 22093 33554 22159 33557
rect 27705 33554 27771 33557
rect 22093 33552 27771 33554
rect 22093 33496 22098 33552
rect 22154 33496 27710 33552
rect 27766 33496 27771 33552
rect 22093 33494 27771 33496
rect 22093 33491 22159 33494
rect 27705 33491 27771 33494
rect 200 33418 800 33448
rect 1761 33418 1827 33421
rect 200 33416 1827 33418
rect 200 33360 1766 33416
rect 1822 33360 1827 33416
rect 200 33358 1827 33360
rect 200 33328 800 33358
rect 1761 33355 1827 33358
rect 22277 33418 22343 33421
rect 26785 33418 26851 33421
rect 22277 33416 26851 33418
rect 22277 33360 22282 33416
rect 22338 33360 26790 33416
rect 26846 33360 26851 33416
rect 22277 33358 26851 33360
rect 22277 33355 22343 33358
rect 26785 33355 26851 33358
rect 25957 33282 26023 33285
rect 25957 33280 28642 33282
rect 25957 33224 25962 33280
rect 26018 33224 28642 33280
rect 25957 33222 28642 33224
rect 25957 33219 26023 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 19241 33146 19307 33149
rect 23289 33146 23355 33149
rect 19241 33144 23355 33146
rect 19241 33088 19246 33144
rect 19302 33088 23294 33144
rect 23350 33088 23355 33144
rect 19241 33086 23355 33088
rect 28582 33146 28642 33222
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 28901 33146 28967 33149
rect 28582 33144 28967 33146
rect 28582 33088 28906 33144
rect 28962 33088 28967 33144
rect 28582 33086 28967 33088
rect 19241 33083 19307 33086
rect 23289 33083 23355 33086
rect 28901 33083 28967 33086
rect 22001 33010 22067 33013
rect 22185 33010 22251 33013
rect 22001 33008 22251 33010
rect 22001 32952 22006 33008
rect 22062 32952 22190 33008
rect 22246 32952 22251 33008
rect 22001 32950 22251 32952
rect 22001 32947 22067 32950
rect 22185 32947 22251 32950
rect 6177 32874 6243 32877
rect 24945 32874 25011 32877
rect 6177 32872 25011 32874
rect 6177 32816 6182 32872
rect 6238 32816 24950 32872
rect 25006 32816 25011 32872
rect 6177 32814 25011 32816
rect 6177 32811 6243 32814
rect 24945 32811 25011 32814
rect 11421 32738 11487 32741
rect 11830 32738 11836 32740
rect 11421 32736 11836 32738
rect 11421 32680 11426 32736
rect 11482 32680 11836 32736
rect 11421 32678 11836 32680
rect 11421 32675 11487 32678
rect 11830 32676 11836 32678
rect 11900 32676 11906 32740
rect 20989 32738 21055 32741
rect 22461 32738 22527 32741
rect 26785 32738 26851 32741
rect 20989 32736 26851 32738
rect 20989 32680 20994 32736
rect 21050 32680 22466 32736
rect 22522 32680 26790 32736
rect 26846 32680 26851 32736
rect 20989 32678 26851 32680
rect 20989 32675 21055 32678
rect 22461 32675 22527 32678
rect 26785 32675 26851 32678
rect 38101 32738 38167 32741
rect 39200 32738 39800 32768
rect 38101 32736 39800 32738
rect 38101 32680 38106 32736
rect 38162 32680 39800 32736
rect 38101 32678 39800 32680
rect 38101 32675 38167 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 21173 32602 21239 32605
rect 26325 32602 26391 32605
rect 21173 32600 26391 32602
rect 21173 32544 21178 32600
rect 21234 32544 26330 32600
rect 26386 32544 26391 32600
rect 21173 32542 26391 32544
rect 21173 32539 21239 32542
rect 26325 32539 26391 32542
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 13721 32058 13787 32061
rect 21081 32058 21147 32061
rect 13721 32056 21147 32058
rect 13721 32000 13726 32056
rect 13782 32000 21086 32056
rect 21142 32000 21147 32056
rect 13721 31998 21147 32000
rect 13721 31995 13787 31998
rect 21081 31995 21147 31998
rect 38285 32058 38351 32061
rect 39200 32058 39800 32088
rect 38285 32056 39800 32058
rect 38285 32000 38290 32056
rect 38346 32000 39800 32056
rect 38285 31998 39800 32000
rect 38285 31995 38351 31998
rect 39200 31968 39800 31998
rect 22737 31786 22803 31789
rect 24761 31786 24827 31789
rect 25497 31786 25563 31789
rect 22737 31784 25563 31786
rect 22737 31728 22742 31784
rect 22798 31728 24766 31784
rect 24822 31728 25502 31784
rect 25558 31728 25563 31784
rect 22737 31726 25563 31728
rect 22737 31723 22803 31726
rect 24761 31723 24827 31726
rect 25497 31723 25563 31726
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 22185 31514 22251 31517
rect 28257 31514 28323 31517
rect 22185 31512 28323 31514
rect 22185 31456 22190 31512
rect 22246 31456 28262 31512
rect 28318 31456 28323 31512
rect 22185 31454 28323 31456
rect 22185 31451 22251 31454
rect 28257 31451 28323 31454
rect 200 31378 800 31408
rect 1761 31378 1827 31381
rect 200 31376 1827 31378
rect 200 31320 1766 31376
rect 1822 31320 1827 31376
rect 200 31318 1827 31320
rect 200 31288 800 31318
rect 1761 31315 1827 31318
rect 5349 31378 5415 31381
rect 25221 31378 25287 31381
rect 5349 31376 25287 31378
rect 5349 31320 5354 31376
rect 5410 31320 25226 31376
rect 25282 31320 25287 31376
rect 5349 31318 25287 31320
rect 5349 31315 5415 31318
rect 25221 31315 25287 31318
rect 17677 31242 17743 31245
rect 23657 31242 23723 31245
rect 17677 31240 23723 31242
rect 17677 31184 17682 31240
rect 17738 31184 23662 31240
rect 23718 31184 23723 31240
rect 17677 31182 23723 31184
rect 17677 31179 17743 31182
rect 23657 31179 23723 31182
rect 25078 31180 25084 31244
rect 25148 31242 25154 31244
rect 25497 31242 25563 31245
rect 25148 31240 25563 31242
rect 25148 31184 25502 31240
rect 25558 31184 25563 31240
rect 25148 31182 25563 31184
rect 25148 31180 25154 31182
rect 25497 31179 25563 31182
rect 19425 31106 19491 31109
rect 22645 31106 22711 31109
rect 19425 31104 22711 31106
rect 19425 31048 19430 31104
rect 19486 31048 22650 31104
rect 22706 31048 22711 31104
rect 19425 31046 22711 31048
rect 19425 31043 19491 31046
rect 22645 31043 22711 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 37457 30698 37523 30701
rect 39200 30698 39800 30728
rect 37457 30696 39800 30698
rect 37457 30640 37462 30696
rect 37518 30640 39800 30696
rect 37457 30638 39800 30640
rect 37457 30635 37523 30638
rect 39200 30608 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 16757 30290 16823 30293
rect 20529 30290 20595 30293
rect 16757 30288 20595 30290
rect 16757 30232 16762 30288
rect 16818 30232 20534 30288
rect 20590 30232 20595 30288
rect 16757 30230 20595 30232
rect 16757 30227 16823 30230
rect 20529 30227 20595 30230
rect 16941 30154 17007 30157
rect 18321 30154 18387 30157
rect 16941 30152 18387 30154
rect 16941 30096 16946 30152
rect 17002 30096 18326 30152
rect 18382 30096 18387 30152
rect 16941 30094 18387 30096
rect 16941 30091 17007 30094
rect 18321 30091 18387 30094
rect 19701 30154 19767 30157
rect 20110 30154 20116 30156
rect 19701 30152 20116 30154
rect 19701 30096 19706 30152
rect 19762 30096 20116 30152
rect 19701 30094 20116 30096
rect 19701 30091 19767 30094
rect 20110 30092 20116 30094
rect 20180 30092 20186 30156
rect 200 30018 800 30048
rect 1761 30018 1827 30021
rect 200 30016 1827 30018
rect 200 29960 1766 30016
rect 1822 29960 1827 30016
rect 200 29958 1827 29960
rect 200 29928 800 29958
rect 1761 29955 1827 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 16297 29882 16363 29885
rect 17769 29882 17835 29885
rect 16297 29880 17835 29882
rect 16297 29824 16302 29880
rect 16358 29824 17774 29880
rect 17830 29824 17835 29880
rect 16297 29822 17835 29824
rect 16297 29819 16363 29822
rect 17769 29819 17835 29822
rect 21541 29882 21607 29885
rect 28717 29882 28783 29885
rect 21541 29880 28783 29882
rect 21541 29824 21546 29880
rect 21602 29824 28722 29880
rect 28778 29824 28783 29880
rect 21541 29822 28783 29824
rect 21541 29819 21607 29822
rect 28717 29819 28783 29822
rect 18137 29746 18203 29749
rect 23381 29746 23447 29749
rect 18137 29744 23447 29746
rect 18137 29688 18142 29744
rect 18198 29688 23386 29744
rect 23442 29688 23447 29744
rect 18137 29686 23447 29688
rect 18137 29683 18203 29686
rect 23381 29683 23447 29686
rect 19333 29610 19399 29613
rect 23749 29610 23815 29613
rect 19333 29608 23815 29610
rect 19333 29552 19338 29608
rect 19394 29552 23754 29608
rect 23810 29552 23815 29608
rect 19333 29550 23815 29552
rect 19333 29547 19399 29550
rect 23749 29547 23815 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 38193 29338 38259 29341
rect 39200 29338 39800 29368
rect 38193 29336 39800 29338
rect 38193 29280 38198 29336
rect 38254 29280 39800 29336
rect 38193 29278 39800 29280
rect 38193 29275 38259 29278
rect 39200 29248 39800 29278
rect 19425 29202 19491 29205
rect 28533 29202 28599 29205
rect 19425 29200 28599 29202
rect 19425 29144 19430 29200
rect 19486 29144 28538 29200
rect 28594 29144 28599 29200
rect 19425 29142 28599 29144
rect 19425 29139 19491 29142
rect 28533 29139 28599 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 15837 28386 15903 28389
rect 17861 28386 17927 28389
rect 15837 28384 17927 28386
rect 15837 28328 15842 28384
rect 15898 28328 17866 28384
rect 17922 28328 17927 28384
rect 15837 28326 17927 28328
rect 15837 28323 15903 28326
rect 17861 28323 17927 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 15745 28114 15811 28117
rect 17861 28114 17927 28117
rect 15745 28112 17927 28114
rect 15745 28056 15750 28112
rect 15806 28056 17866 28112
rect 17922 28056 17927 28112
rect 15745 28054 17927 28056
rect 15745 28051 15811 28054
rect 17861 28051 17927 28054
rect 21909 27978 21975 27981
rect 24853 27978 24919 27981
rect 21909 27976 24919 27978
rect 21909 27920 21914 27976
rect 21970 27920 24858 27976
rect 24914 27920 24919 27976
rect 21909 27918 24919 27920
rect 21909 27915 21975 27918
rect 24853 27915 24919 27918
rect 38193 27978 38259 27981
rect 39200 27978 39800 28008
rect 38193 27976 39800 27978
rect 38193 27920 38198 27976
rect 38254 27920 39800 27976
rect 38193 27918 39800 27920
rect 38193 27915 38259 27918
rect 39200 27888 39800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 2221 27708 2287 27709
rect 2221 27704 2268 27708
rect 2332 27706 2338 27708
rect 17953 27706 18019 27709
rect 18781 27706 18847 27709
rect 2221 27648 2226 27704
rect 2221 27644 2268 27648
rect 2332 27646 2378 27706
rect 17953 27704 18847 27706
rect 17953 27648 17958 27704
rect 18014 27648 18786 27704
rect 18842 27648 18847 27704
rect 17953 27646 18847 27648
rect 2332 27644 2338 27646
rect 2221 27643 2287 27644
rect 17953 27643 18019 27646
rect 18781 27643 18847 27646
rect 11830 27508 11836 27572
rect 11900 27570 11906 27572
rect 16481 27570 16547 27573
rect 11900 27568 16547 27570
rect 11900 27512 16486 27568
rect 16542 27512 16547 27568
rect 11900 27510 16547 27512
rect 11900 27508 11906 27510
rect 16481 27507 16547 27510
rect 21357 27570 21423 27573
rect 23381 27570 23447 27573
rect 21357 27568 23447 27570
rect 21357 27512 21362 27568
rect 21418 27512 23386 27568
rect 23442 27512 23447 27568
rect 21357 27510 23447 27512
rect 21357 27507 21423 27510
rect 23381 27507 23447 27510
rect 17769 27434 17835 27437
rect 21541 27434 21607 27437
rect 17769 27432 21607 27434
rect 17769 27376 17774 27432
rect 17830 27376 21546 27432
rect 21602 27376 21607 27432
rect 17769 27374 21607 27376
rect 17769 27371 17835 27374
rect 21541 27371 21607 27374
rect 21817 27434 21883 27437
rect 25313 27434 25379 27437
rect 21817 27432 25379 27434
rect 21817 27376 21822 27432
rect 21878 27376 25318 27432
rect 25374 27376 25379 27432
rect 21817 27374 25379 27376
rect 21817 27371 21883 27374
rect 25313 27371 25379 27374
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 38193 27298 38259 27301
rect 39200 27298 39800 27328
rect 38193 27296 39800 27298
rect 38193 27240 38198 27296
rect 38254 27240 39800 27296
rect 38193 27238 39800 27240
rect 38193 27235 38259 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 13721 27026 13787 27029
rect 27245 27026 27311 27029
rect 13721 27024 27311 27026
rect 13721 26968 13726 27024
rect 13782 26968 27250 27024
rect 27306 26968 27311 27024
rect 13721 26966 27311 26968
rect 13721 26963 13787 26966
rect 27245 26963 27311 26966
rect 15377 26754 15443 26757
rect 18781 26754 18847 26757
rect 15377 26752 18847 26754
rect 15377 26696 15382 26752
rect 15438 26696 18786 26752
rect 18842 26696 18847 26752
rect 15377 26694 18847 26696
rect 15377 26691 15443 26694
rect 18781 26691 18847 26694
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1669 26618 1735 26621
rect 200 26616 1735 26618
rect 200 26560 1674 26616
rect 1730 26560 1735 26616
rect 200 26558 1735 26560
rect 200 26528 800 26558
rect 1669 26555 1735 26558
rect 1853 26484 1919 26485
rect 1853 26480 1900 26484
rect 1964 26482 1970 26484
rect 20069 26482 20135 26485
rect 25773 26482 25839 26485
rect 1853 26424 1858 26480
rect 1853 26420 1900 26424
rect 1964 26422 2010 26482
rect 20069 26480 25839 26482
rect 20069 26424 20074 26480
rect 20130 26424 25778 26480
rect 25834 26424 25839 26480
rect 20069 26422 25839 26424
rect 1964 26420 1970 26422
rect 1853 26419 1919 26420
rect 20069 26419 20135 26422
rect 25773 26419 25839 26422
rect 3417 26346 3483 26349
rect 3550 26346 3556 26348
rect 3417 26344 3556 26346
rect 3417 26288 3422 26344
rect 3478 26288 3556 26344
rect 3417 26286 3556 26288
rect 3417 26283 3483 26286
rect 3550 26284 3556 26286
rect 3620 26284 3626 26348
rect 16941 26346 17007 26349
rect 17401 26346 17467 26349
rect 16941 26344 17467 26346
rect 16941 26288 16946 26344
rect 17002 26288 17406 26344
rect 17462 26288 17467 26344
rect 16941 26286 17467 26288
rect 16941 26283 17007 26286
rect 17401 26283 17467 26286
rect 23841 26346 23907 26349
rect 23974 26346 23980 26348
rect 23841 26344 23980 26346
rect 23841 26288 23846 26344
rect 23902 26288 23980 26344
rect 23841 26286 23980 26288
rect 23841 26283 23907 26286
rect 23974 26284 23980 26286
rect 24044 26284 24050 26348
rect 10777 26210 10843 26213
rect 11605 26210 11671 26213
rect 18781 26210 18847 26213
rect 10777 26208 18847 26210
rect 10777 26152 10782 26208
rect 10838 26152 11610 26208
rect 11666 26152 18786 26208
rect 18842 26152 18847 26208
rect 10777 26150 18847 26152
rect 10777 26147 10843 26150
rect 11605 26147 11671 26150
rect 18781 26147 18847 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 38285 25938 38351 25941
rect 39200 25938 39800 25968
rect 38285 25936 39800 25938
rect 38285 25880 38290 25936
rect 38346 25880 39800 25936
rect 38285 25878 39800 25880
rect 38285 25875 38351 25878
rect 39200 25848 39800 25878
rect 18321 25666 18387 25669
rect 19149 25666 19215 25669
rect 18321 25664 19215 25666
rect 18321 25608 18326 25664
rect 18382 25608 19154 25664
rect 19210 25608 19215 25664
rect 18321 25606 19215 25608
rect 18321 25603 18387 25606
rect 19149 25603 19215 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19885 25394 19951 25397
rect 25497 25394 25563 25397
rect 19885 25392 25563 25394
rect 19885 25336 19890 25392
rect 19946 25336 25502 25392
rect 25558 25336 25563 25392
rect 19885 25334 25563 25336
rect 19885 25331 19951 25334
rect 25497 25331 25563 25334
rect 200 25258 800 25288
rect 1761 25258 1827 25261
rect 200 25256 1827 25258
rect 200 25200 1766 25256
rect 1822 25200 1827 25256
rect 200 25198 1827 25200
rect 200 25168 800 25198
rect 1761 25195 1827 25198
rect 19793 25258 19859 25261
rect 20437 25258 20503 25261
rect 19793 25256 20503 25258
rect 19793 25200 19798 25256
rect 19854 25200 20442 25256
rect 20498 25200 20503 25256
rect 19793 25198 20503 25200
rect 19793 25195 19859 25198
rect 20437 25195 20503 25198
rect 6361 25122 6427 25125
rect 6494 25122 6500 25124
rect 6361 25120 6500 25122
rect 6361 25064 6366 25120
rect 6422 25064 6500 25120
rect 6361 25062 6500 25064
rect 6361 25059 6427 25062
rect 6494 25060 6500 25062
rect 6564 25122 6570 25124
rect 6821 25122 6887 25125
rect 6564 25120 6887 25122
rect 6564 25064 6826 25120
rect 6882 25064 6887 25120
rect 6564 25062 6887 25064
rect 6564 25060 6570 25062
rect 6821 25059 6887 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 1577 24986 1643 24989
rect 1710 24986 1716 24988
rect 1577 24984 1716 24986
rect 1577 24928 1582 24984
rect 1638 24928 1716 24984
rect 1577 24926 1716 24928
rect 1577 24923 1643 24926
rect 1710 24924 1716 24926
rect 1780 24924 1786 24988
rect 20161 24714 20227 24717
rect 24945 24714 25011 24717
rect 20161 24712 25011 24714
rect 20161 24656 20166 24712
rect 20222 24656 24950 24712
rect 25006 24656 25011 24712
rect 20161 24654 25011 24656
rect 20161 24651 20227 24654
rect 24945 24651 25011 24654
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 20621 24170 20687 24173
rect 23105 24170 23171 24173
rect 20621 24168 23171 24170
rect 20621 24112 20626 24168
rect 20682 24112 23110 24168
rect 23166 24112 23171 24168
rect 20621 24110 23171 24112
rect 20621 24107 20687 24110
rect 23105 24107 23171 24110
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 38285 23898 38351 23901
rect 39200 23898 39800 23928
rect 38285 23896 39800 23898
rect 38285 23840 38290 23896
rect 38346 23840 39800 23896
rect 38285 23838 39800 23840
rect 38285 23835 38351 23838
rect 39200 23808 39800 23838
rect 20621 23626 20687 23629
rect 22921 23626 22987 23629
rect 20621 23624 22987 23626
rect 20621 23568 20626 23624
rect 20682 23568 22926 23624
rect 22982 23568 22987 23624
rect 20621 23566 22987 23568
rect 20621 23563 20687 23566
rect 22921 23563 22987 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 20110 23292 20116 23356
rect 20180 23354 20186 23356
rect 20713 23354 20779 23357
rect 20180 23352 20779 23354
rect 20180 23296 20718 23352
rect 20774 23296 20779 23352
rect 20180 23294 20779 23296
rect 20180 23292 20186 23294
rect 20713 23291 20779 23294
rect 200 23218 800 23248
rect 1393 23218 1459 23221
rect 200 23216 1459 23218
rect 200 23160 1398 23216
rect 1454 23160 1459 23216
rect 200 23158 1459 23160
rect 200 23128 800 23158
rect 1393 23155 1459 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 3785 21994 3851 21997
rect 8385 21994 8451 21997
rect 3785 21992 8451 21994
rect 3785 21936 3790 21992
rect 3846 21936 8390 21992
rect 8446 21936 8451 21992
rect 3785 21934 8451 21936
rect 3785 21931 3851 21934
rect 8385 21931 8451 21934
rect 200 21858 800 21888
rect 1761 21858 1827 21861
rect 200 21856 1827 21858
rect 200 21800 1766 21856
rect 1822 21800 1827 21856
rect 200 21798 1827 21800
rect 200 21768 800 21798
rect 1761 21795 1827 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4245 21450 4311 21453
rect 4838 21450 4844 21452
rect 4245 21448 4844 21450
rect 4245 21392 4250 21448
rect 4306 21392 4844 21448
rect 4245 21390 4844 21392
rect 4245 21387 4311 21390
rect 4838 21388 4844 21390
rect 4908 21450 4914 21452
rect 5257 21450 5323 21453
rect 4908 21448 5323 21450
rect 4908 21392 5262 21448
rect 5318 21392 5323 21448
rect 4908 21390 5323 21392
rect 4908 21388 4914 21390
rect 5257 21387 5323 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 38285 21178 38351 21181
rect 39200 21178 39800 21208
rect 38285 21176 39800 21178
rect 38285 21120 38290 21176
rect 38346 21120 39800 21176
rect 38285 21118 39800 21120
rect 38285 21115 38351 21118
rect 39200 21088 39800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 38285 20498 38351 20501
rect 39200 20498 39800 20528
rect 38285 20496 39800 20498
rect 38285 20440 38290 20496
rect 38346 20440 39800 20496
rect 38285 20438 39800 20440
rect 38285 20435 38351 20438
rect 39200 20408 39800 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 21817 19954 21883 19957
rect 24945 19954 25011 19957
rect 25078 19954 25084 19956
rect 21817 19952 25084 19954
rect 21817 19896 21822 19952
rect 21878 19896 24950 19952
rect 25006 19896 25084 19952
rect 21817 19894 25084 19896
rect 21817 19891 21883 19894
rect 24945 19891 25011 19894
rect 25078 19892 25084 19894
rect 25148 19892 25154 19956
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 19138 800 19168
rect 1393 19138 1459 19141
rect 200 19136 1459 19138
rect 200 19080 1398 19136
rect 1454 19080 1459 19136
rect 200 19078 1459 19080
rect 200 19048 800 19078
rect 1393 19075 1459 19078
rect 38285 19138 38351 19141
rect 39200 19138 39800 19168
rect 38285 19136 39800 19138
rect 38285 19080 38290 19136
rect 38346 19080 39800 19136
rect 38285 19078 39800 19080
rect 38285 19075 38351 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 200 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 1761 18458 1827 18461
rect 200 18456 1827 18458
rect 200 18400 1766 18456
rect 1822 18400 1827 18456
rect 200 18398 1827 18400
rect 200 18368 800 18398
rect 1761 18395 1827 18398
rect 4153 18186 4219 18189
rect 4521 18186 4587 18189
rect 4654 18186 4660 18188
rect 4153 18184 4660 18186
rect 4153 18128 4158 18184
rect 4214 18128 4526 18184
rect 4582 18128 4660 18184
rect 4153 18126 4660 18128
rect 4153 18123 4219 18126
rect 4521 18123 4587 18126
rect 4654 18124 4660 18126
rect 4724 18124 4730 18188
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 38285 17778 38351 17781
rect 39200 17778 39800 17808
rect 38285 17776 39800 17778
rect 38285 17720 38290 17776
rect 38346 17720 39800 17776
rect 38285 17718 39800 17720
rect 38285 17715 38351 17718
rect 39200 17688 39800 17718
rect 24025 17644 24091 17645
rect 23974 17642 23980 17644
rect 23934 17582 23980 17642
rect 24044 17640 24091 17644
rect 24086 17584 24091 17640
rect 23974 17580 23980 17582
rect 24044 17580 24091 17584
rect 24025 17579 24091 17580
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 9581 17234 9647 17237
rect 10961 17234 11027 17237
rect 9581 17232 11027 17234
rect 9581 17176 9586 17232
rect 9642 17176 10966 17232
rect 11022 17176 11027 17232
rect 9581 17174 11027 17176
rect 9581 17171 9647 17174
rect 10961 17171 11027 17174
rect 200 17098 800 17128
rect 1669 17098 1735 17101
rect 200 17096 1735 17098
rect 200 17040 1674 17096
rect 1730 17040 1735 17096
rect 200 17038 1735 17040
rect 200 17008 800 17038
rect 1669 17035 1735 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 2589 16692 2655 16693
rect 2589 16688 2636 16692
rect 2700 16690 2706 16692
rect 2589 16632 2594 16688
rect 2589 16628 2636 16632
rect 2700 16630 2746 16690
rect 2700 16628 2706 16630
rect 2589 16627 2655 16628
rect 21817 16554 21883 16557
rect 23473 16554 23539 16557
rect 21817 16552 23539 16554
rect 21817 16496 21822 16552
rect 21878 16496 23478 16552
rect 23534 16496 23539 16552
rect 21817 16494 23539 16496
rect 21817 16491 21883 16494
rect 23473 16491 23539 16494
rect 38101 16418 38167 16421
rect 39200 16418 39800 16448
rect 38101 16416 39800 16418
rect 38101 16360 38106 16416
rect 38162 16360 39800 16416
rect 38101 16358 39800 16360
rect 38101 16355 38167 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 39200 16328 39800 16358
rect 19570 16287 19886 16288
rect 3969 16146 4035 16149
rect 8753 16146 8819 16149
rect 3969 16144 8819 16146
rect 3969 16088 3974 16144
rect 4030 16088 8758 16144
rect 8814 16088 8819 16144
rect 3969 16086 8819 16088
rect 3969 16083 4035 16086
rect 8753 16083 8819 16086
rect 9673 16146 9739 16149
rect 11830 16146 11836 16148
rect 9673 16144 11836 16146
rect 9673 16088 9678 16144
rect 9734 16088 11836 16144
rect 9673 16086 11836 16088
rect 9673 16083 9739 16086
rect 11830 16084 11836 16086
rect 11900 16084 11906 16148
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 38285 15738 38351 15741
rect 39200 15738 39800 15768
rect 38285 15736 39800 15738
rect 38285 15680 38290 15736
rect 38346 15680 39800 15736
rect 38285 15678 39800 15680
rect 38285 15675 38351 15678
rect 39200 15648 39800 15678
rect 3918 15268 3924 15332
rect 3988 15330 3994 15332
rect 7649 15330 7715 15333
rect 3988 15328 7715 15330
rect 3988 15272 7654 15328
rect 7710 15272 7715 15328
rect 3988 15270 7715 15272
rect 3988 15268 3994 15270
rect 7649 15267 7715 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 10409 15194 10475 15197
rect 18413 15194 18479 15197
rect 10409 15192 18479 15194
rect 10409 15136 10414 15192
rect 10470 15136 18418 15192
rect 18474 15136 18479 15192
rect 10409 15134 18479 15136
rect 10409 15131 10475 15134
rect 18413 15131 18479 15134
rect 200 15058 800 15088
rect 1761 15058 1827 15061
rect 200 15056 1827 15058
rect 200 15000 1766 15056
rect 1822 15000 1827 15056
rect 200 14998 1827 15000
rect 200 14968 800 14998
rect 1761 14995 1827 14998
rect 16665 15058 16731 15061
rect 18045 15058 18111 15061
rect 16665 15056 18111 15058
rect 16665 15000 16670 15056
rect 16726 15000 18050 15056
rect 18106 15000 18111 15056
rect 16665 14998 18111 15000
rect 16665 14995 16731 14998
rect 18045 14995 18111 14998
rect 9857 14922 9923 14925
rect 19057 14922 19123 14925
rect 9857 14920 19123 14922
rect 9857 14864 9862 14920
rect 9918 14864 19062 14920
rect 19118 14864 19123 14920
rect 9857 14862 19123 14864
rect 9857 14859 9923 14862
rect 19057 14859 19123 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 38285 14378 38351 14381
rect 39200 14378 39800 14408
rect 38285 14376 39800 14378
rect 38285 14320 38290 14376
rect 38346 14320 39800 14376
rect 38285 14318 39800 14320
rect 38285 14315 38351 14318
rect 39200 14288 39800 14318
rect 3417 14242 3483 14245
rect 7281 14242 7347 14245
rect 3417 14240 7347 14242
rect 3417 14184 3422 14240
rect 3478 14184 7286 14240
rect 7342 14184 7347 14240
rect 3417 14182 7347 14184
rect 3417 14179 3483 14182
rect 7281 14179 7347 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13698 800 13728
rect 1761 13698 1827 13701
rect 200 13696 1827 13698
rect 200 13640 1766 13696
rect 1822 13640 1827 13696
rect 200 13638 1827 13640
rect 200 13608 800 13638
rect 1761 13635 1827 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 6494 13500 6500 13564
rect 6564 13562 6570 13564
rect 15653 13562 15719 13565
rect 6564 13560 15719 13562
rect 6564 13504 15658 13560
rect 15714 13504 15719 13560
rect 6564 13502 15719 13504
rect 6564 13500 6570 13502
rect 15653 13499 15719 13502
rect 2630 13364 2636 13428
rect 2700 13426 2706 13428
rect 14641 13426 14707 13429
rect 2700 13424 14707 13426
rect 2700 13368 14646 13424
rect 14702 13368 14707 13424
rect 2700 13366 14707 13368
rect 2700 13364 2706 13366
rect 14641 13363 14707 13366
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 38193 13018 38259 13021
rect 39200 13018 39800 13048
rect 38193 13016 39800 13018
rect 38193 12960 38198 13016
rect 38254 12960 39800 13016
rect 38193 12958 39800 12960
rect 38193 12955 38259 12958
rect 39200 12928 39800 12958
rect 4654 12820 4660 12884
rect 4724 12882 4730 12884
rect 4889 12882 4955 12885
rect 4724 12880 4955 12882
rect 4724 12824 4894 12880
rect 4950 12824 4955 12880
rect 4724 12822 4955 12824
rect 4724 12820 4730 12822
rect 4889 12819 4955 12822
rect 10041 12610 10107 12613
rect 10501 12610 10567 12613
rect 10041 12608 10567 12610
rect 10041 12552 10046 12608
rect 10102 12552 10506 12608
rect 10562 12552 10567 12608
rect 10041 12550 10567 12552
rect 10041 12547 10107 12550
rect 10501 12547 10567 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 1710 12140 1716 12204
rect 1780 12202 1786 12204
rect 13353 12202 13419 12205
rect 1780 12200 13419 12202
rect 1780 12144 13358 12200
rect 13414 12144 13419 12200
rect 1780 12142 13419 12144
rect 1780 12140 1786 12142
rect 13353 12139 13419 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 200 11658 800 11688
rect 2865 11658 2931 11661
rect 200 11656 2931 11658
rect 200 11600 2870 11656
rect 2926 11600 2931 11656
rect 200 11598 2931 11600
rect 200 11568 800 11598
rect 2865 11595 2931 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 3509 10980 3575 10981
rect 3509 10976 3556 10980
rect 3620 10978 3626 10980
rect 37181 10978 37247 10981
rect 39200 10978 39800 11008
rect 3509 10920 3514 10976
rect 3509 10916 3556 10920
rect 3620 10918 3666 10978
rect 37181 10976 39800 10978
rect 37181 10920 37186 10976
rect 37242 10920 39800 10976
rect 37181 10918 39800 10920
rect 3620 10916 3626 10918
rect 3509 10915 3575 10916
rect 37181 10915 37247 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 2773 10298 2839 10301
rect 200 10296 2839 10298
rect 200 10240 2778 10296
rect 2834 10240 2839 10296
rect 200 10238 2839 10240
rect 200 10208 800 10238
rect 2773 10235 2839 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 2221 9620 2287 9621
rect 2221 9616 2268 9620
rect 2332 9618 2338 9620
rect 2589 9618 2655 9621
rect 4838 9618 4844 9620
rect 2221 9560 2226 9616
rect 2221 9556 2268 9560
rect 2332 9558 2378 9618
rect 2589 9616 4844 9618
rect 2589 9560 2594 9616
rect 2650 9560 4844 9616
rect 2589 9558 4844 9560
rect 2332 9556 2338 9558
rect 2221 9555 2287 9556
rect 2589 9555 2655 9558
rect 4838 9556 4844 9558
rect 4908 9556 4914 9620
rect 38193 9618 38259 9621
rect 39200 9618 39800 9648
rect 38193 9616 39800 9618
rect 38193 9560 38198 9616
rect 38254 9560 39800 9616
rect 38193 9558 39800 9560
rect 38193 9555 38259 9558
rect 39200 9528 39800 9558
rect 1894 9420 1900 9484
rect 1964 9482 1970 9484
rect 34329 9482 34395 9485
rect 1964 9480 34395 9482
rect 1964 9424 34334 9480
rect 34390 9424 34395 9480
rect 1964 9422 34395 9424
rect 1964 9420 1970 9422
rect 34329 9419 34395 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 200 8938 800 8968
rect 2773 8938 2839 8941
rect 200 8936 2839 8938
rect 200 8880 2778 8936
rect 2834 8880 2839 8936
rect 200 8878 2839 8880
rect 200 8848 800 8878
rect 2773 8875 2839 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 38101 8258 38167 8261
rect 39200 8258 39800 8288
rect 38101 8256 39800 8258
rect 38101 8200 38106 8256
rect 38162 8200 39800 8256
rect 38101 8198 39800 8200
rect 38101 8195 38167 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 39800 8198
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1577 7578 1643 7581
rect 200 7576 1643 7578
rect 200 7520 1582 7576
rect 1638 7520 1643 7576
rect 200 7518 1643 7520
rect 200 7488 800 7518
rect 1577 7515 1643 7518
rect 38193 7578 38259 7581
rect 39200 7578 39800 7608
rect 38193 7576 39800 7578
rect 38193 7520 38198 7576
rect 38254 7520 39800 7576
rect 38193 7518 39800 7520
rect 38193 7515 38259 7518
rect 39200 7488 39800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1669 6898 1735 6901
rect 200 6896 1735 6898
rect 200 6840 1674 6896
rect 1730 6840 1735 6896
rect 200 6838 1735 6840
rect 200 6808 800 6838
rect 1669 6835 1735 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 37457 6218 37523 6221
rect 39200 6218 39800 6248
rect 37457 6216 39800 6218
rect 37457 6160 37462 6216
rect 37518 6160 39800 6216
rect 37457 6158 39800 6160
rect 37457 6155 37523 6158
rect 39200 6128 39800 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5538 800 5568
rect 1761 5538 1827 5541
rect 200 5536 1827 5538
rect 200 5480 1766 5536
rect 1822 5480 1827 5536
rect 200 5478 1827 5480
rect 200 5448 800 5478
rect 1761 5475 1827 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 38193 4858 38259 4861
rect 39200 4858 39800 4888
rect 38193 4856 39800 4858
rect 38193 4800 38198 4856
rect 38254 4800 39800 4856
rect 38193 4798 39800 4800
rect 38193 4795 38259 4798
rect 39200 4768 39800 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 200 4178 800 4208
rect 1669 4178 1735 4181
rect 200 4176 1735 4178
rect 200 4120 1674 4176
rect 1730 4120 1735 4176
rect 200 4118 1735 4120
rect 200 4088 800 4118
rect 1669 4115 1735 4118
rect 38193 4178 38259 4181
rect 39200 4178 39800 4208
rect 38193 4176 39800 4178
rect 38193 4120 38198 4176
rect 38254 4120 39800 4176
rect 38193 4118 39800 4120
rect 38193 4115 38259 4118
rect 39200 4088 39800 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3528
rect 1761 3498 1827 3501
rect 200 3496 1827 3498
rect 200 3440 1766 3496
rect 1822 3440 1827 3496
rect 200 3438 1827 3440
rect 200 3408 800 3438
rect 1761 3435 1827 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 37457 2818 37523 2821
rect 39200 2818 39800 2848
rect 37457 2816 39800 2818
rect 37457 2760 37462 2816
rect 37518 2760 39800 2816
rect 37457 2758 39800 2760
rect 37457 2755 37523 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 200 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 2497 2138 2563 2141
rect 200 2136 2563 2138
rect 200 2080 2502 2136
rect 2558 2080 2563 2136
rect 200 2078 2563 2080
rect 200 2048 800 2078
rect 2497 2075 2563 2078
rect 37457 1458 37523 1461
rect 39200 1458 39800 1488
rect 37457 1456 39800 1458
rect 37457 1400 37462 1456
rect 37518 1400 39800 1456
rect 37457 1398 39800 1400
rect 37457 1395 37523 1398
rect 39200 1368 39800 1398
rect 200 778 800 808
rect 1669 778 1735 781
rect 200 776 1735 778
rect 200 720 1674 776
rect 1730 720 1735 776
rect 200 718 1735 720
rect 200 688 800 718
rect 1669 715 1735 718
rect 38193 778 38259 781
rect 39200 778 39800 808
rect 38193 776 39800 778
rect 38193 720 38198 776
rect 38254 720 39800 776
rect 38193 718 39800 720
rect 38193 715 38259 718
rect 39200 688 39800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 3924 34580 3988 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 11836 32676 11900 32740
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 25084 31180 25148 31244
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 20116 30092 20180 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 2268 27704 2332 27708
rect 2268 27648 2282 27704
rect 2282 27648 2332 27704
rect 2268 27644 2332 27648
rect 11836 27508 11900 27572
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 1900 26480 1964 26484
rect 1900 26424 1914 26480
rect 1914 26424 1964 26480
rect 1900 26420 1964 26424
rect 3556 26284 3620 26348
rect 23980 26284 24044 26348
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 6500 25060 6564 25124
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 1716 24924 1780 24988
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 20116 23292 20180 23356
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4844 21388 4908 21452
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 25084 19892 25148 19956
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4660 18124 4724 18188
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 23980 17640 24044 17644
rect 23980 17584 24030 17640
rect 24030 17584 24044 17640
rect 23980 17580 24044 17584
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 2636 16688 2700 16692
rect 2636 16632 2650 16688
rect 2650 16632 2700 16688
rect 2636 16628 2700 16632
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 11836 16084 11900 16148
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 3924 15268 3988 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 6500 13500 6564 13564
rect 2636 13364 2700 13428
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4660 12820 4724 12884
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 1716 12140 1780 12204
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 3556 10976 3620 10980
rect 3556 10920 3570 10976
rect 3570 10920 3620 10976
rect 3556 10916 3620 10920
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 2268 9616 2332 9620
rect 2268 9560 2282 9616
rect 2282 9560 2332 9616
rect 2268 9556 2332 9560
rect 4844 9556 4908 9620
rect 1900 9420 1964 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 3923 34644 3989 34645
rect 3923 34580 3924 34644
rect 3988 34580 3989 34644
rect 3923 34579 3989 34580
rect 2267 27708 2333 27709
rect 2267 27644 2268 27708
rect 2332 27644 2333 27708
rect 2267 27643 2333 27644
rect 1899 26484 1965 26485
rect 1899 26420 1900 26484
rect 1964 26420 1965 26484
rect 1899 26419 1965 26420
rect 1715 24988 1781 24989
rect 1715 24924 1716 24988
rect 1780 24924 1781 24988
rect 1715 24923 1781 24924
rect 1718 12205 1778 24923
rect 1715 12204 1781 12205
rect 1715 12140 1716 12204
rect 1780 12140 1781 12204
rect 1715 12139 1781 12140
rect 1902 9485 1962 26419
rect 2270 9621 2330 27643
rect 3555 26348 3621 26349
rect 3555 26284 3556 26348
rect 3620 26284 3621 26348
rect 3555 26283 3621 26284
rect 2635 16692 2701 16693
rect 2635 16628 2636 16692
rect 2700 16628 2701 16692
rect 2635 16627 2701 16628
rect 2638 13429 2698 16627
rect 2635 13428 2701 13429
rect 2635 13364 2636 13428
rect 2700 13364 2701 13428
rect 2635 13363 2701 13364
rect 3558 10981 3618 26283
rect 3926 15333 3986 34579
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 11835 32740 11901 32741
rect 11835 32676 11836 32740
rect 11900 32676 11901 32740
rect 11835 32675 11901 32676
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 11838 27573 11898 32675
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 25083 31244 25149 31245
rect 25083 31180 25084 31244
rect 25148 31180 25149 31244
rect 25083 31179 25149 31180
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 20115 30156 20181 30157
rect 20115 30092 20116 30156
rect 20180 30092 20181 30156
rect 20115 30091 20181 30092
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 11835 27572 11901 27573
rect 11835 27508 11836 27572
rect 11900 27508 11901 27572
rect 11835 27507 11901 27508
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 6499 25124 6565 25125
rect 6499 25060 6500 25124
rect 6564 25060 6565 25124
rect 6499 25059 6565 25060
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4843 21452 4909 21453
rect 4843 21388 4844 21452
rect 4908 21388 4909 21452
rect 4843 21387 4909 21388
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4659 18188 4725 18189
rect 4659 18124 4660 18188
rect 4724 18124 4725 18188
rect 4659 18123 4725 18124
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 3923 15332 3989 15333
rect 3923 15268 3924 15332
rect 3988 15268 3989 15332
rect 3923 15267 3989 15268
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4662 12885 4722 18123
rect 4659 12884 4725 12885
rect 4659 12820 4660 12884
rect 4724 12820 4725 12884
rect 4659 12819 4725 12820
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 3555 10980 3621 10981
rect 3555 10916 3556 10980
rect 3620 10916 3621 10980
rect 3555 10915 3621 10916
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 2267 9620 2333 9621
rect 2267 9556 2268 9620
rect 2332 9556 2333 9620
rect 2267 9555 2333 9556
rect 1899 9484 1965 9485
rect 1899 9420 1900 9484
rect 1964 9420 1965 9484
rect 1899 9419 1965 9420
rect 4208 9280 4528 10304
rect 4846 9621 4906 21387
rect 6502 13565 6562 25059
rect 11838 16149 11898 27507
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 20118 23357 20178 30091
rect 23979 26348 24045 26349
rect 23979 26284 23980 26348
rect 24044 26284 24045 26348
rect 23979 26283 24045 26284
rect 20115 23356 20181 23357
rect 20115 23292 20116 23356
rect 20180 23292 20181 23356
rect 20115 23291 20181 23292
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 23982 17645 24042 26283
rect 25086 19957 25146 31179
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 25083 19956 25149 19957
rect 25083 19892 25084 19956
rect 25148 19892 25149 19956
rect 25083 19891 25149 19892
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 23979 17644 24045 17645
rect 23979 17580 23980 17644
rect 24044 17580 24045 17644
rect 23979 17579 24045 17580
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 11835 16148 11901 16149
rect 11835 16084 11836 16148
rect 11900 16084 11901 16148
rect 11835 16083 11901 16084
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 6499 13564 6565 13565
rect 6499 13500 6500 13564
rect 6564 13500 6565 13564
rect 6499 13499 6565 13500
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 4843 9620 4909 9621
rect 4843 9556 4844 9620
rect 4908 9556 4909 9620
rect 4843 9555 4909 9556
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 2116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 7636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1667941163
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1667941163
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1667941163
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127
timestamp 1667941163
transform 1 0 12788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_154
timestamp 1667941163
transform 1 0 15272 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1667941163
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1667941163
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1667941163
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_238
timestamp 1667941163
transform 1 0 23000 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_266
timestamp 1667941163
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1667941163
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_294
timestamp 1667941163
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_323
timestamp 1667941163
transform 1 0 30820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_351
timestamp 1667941163
transform 1 0 33396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1667941163
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_379
timestamp 1667941163
transform 1 0 35972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1667941163
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_16
timestamp 1667941163
transform 1 0 2576 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1667941163
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_174
timestamp 1667941163
transform 1 0 17112 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_186
timestamp 1667941163
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_190
timestamp 1667941163
transform 1 0 18584 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_194
timestamp 1667941163
transform 1 0 18952 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_206
timestamp 1667941163
transform 1 0 20056 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1667941163
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_265
timestamp 1667941163
transform 1 0 25484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1667941163
transform 1 0 25852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1667941163
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1667941163
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1667941163
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_393
timestamp 1667941163
transform 1 0 37260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_9
timestamp 1667941163
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1667941163
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_351
timestamp 1667941163
transform 1 0 33396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_371
timestamp 1667941163
transform 1 0 35236 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_375
timestamp 1667941163
transform 1 0 35604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_387
timestamp 1667941163
transform 1 0 36708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_399
timestamp 1667941163
transform 1 0 37812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_35
timestamp 1667941163
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_40
timestamp 1667941163
transform 1 0 4784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1667941163
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_92
timestamp 1667941163
transform 1 0 9568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1667941163
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_258
timestamp 1667941163
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_270
timestamp 1667941163
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1667941163
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_9
timestamp 1667941163
transform 1 0 1932 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_17
timestamp 1667941163
transform 1 0 2668 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1667941163
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1667941163
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_39
timestamp 1667941163
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_51
timestamp 1667941163
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_63
timestamp 1667941163
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1667941163
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_149
timestamp 1667941163
transform 1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_161
timestamp 1667941163
transform 1 0 15916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_173
timestamp 1667941163
transform 1 0 17020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_185
timestamp 1667941163
transform 1 0 18124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1667941163
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1667941163
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_156
timestamp 1667941163
transform 1 0 15456 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1667941163
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_370
timestamp 1667941163
transform 1 0 35144 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_382
timestamp 1667941163
transform 1 0 36248 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_394
timestamp 1667941163
transform 1 0 37352 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1667941163
transform 1 0 38456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_22
timestamp 1667941163
transform 1 0 3128 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_34
timestamp 1667941163
transform 1 0 4232 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1667941163
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_143
timestamp 1667941163
transform 1 0 14260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_155
timestamp 1667941163
transform 1 0 15364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_174
timestamp 1667941163
transform 1 0 17112 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_186
timestamp 1667941163
transform 1 0 18216 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_198
timestamp 1667941163
transform 1 0 19320 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_210
timestamp 1667941163
transform 1 0 20424 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_370
timestamp 1667941163
transform 1 0 35144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_382
timestamp 1667941163
transform 1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1667941163
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_21
timestamp 1667941163
transform 1 0 3036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1667941163
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_46
timestamp 1667941163
transform 1 0 5336 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_58
timestamp 1667941163
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_70
timestamp 1667941163
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_147
timestamp 1667941163
transform 1 0 14628 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_151
timestamp 1667941163
transform 1 0 14996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_163
timestamp 1667941163
transform 1 0 16100 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_175
timestamp 1667941163
transform 1 0 17204 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1667941163
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1667941163
transform 1 0 20700 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_217
timestamp 1667941163
transform 1 0 21068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_229
timestamp 1667941163
transform 1 0 22172 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_241
timestamp 1667941163
transform 1 0 23276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 1667941163
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_270
timestamp 1667941163
transform 1 0 25944 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_282
timestamp 1667941163
transform 1 0 27048 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_294
timestamp 1667941163
transform 1 0 28152 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_302
timestamp 1667941163
transform 1 0 28888 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1667941163
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_353
timestamp 1667941163
transform 1 0 33580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_358
timestamp 1667941163
transform 1 0 34040 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1667941163
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_18
timestamp 1667941163
transform 1 0 2760 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_145
timestamp 1667941163
transform 1 0 14444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_213
timestamp 1667941163
transform 1 0 20700 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_286
timestamp 1667941163
transform 1 0 27416 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_298
timestamp 1667941163
transform 1 0 28520 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_310
timestamp 1667941163
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_322
timestamp 1667941163
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1667941163
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_8
timestamp 1667941163
transform 1 0 1840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1667941163
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 1667941163
transform 1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_50
timestamp 1667941163
transform 1 0 5704 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_62
timestamp 1667941163
transform 1 0 6808 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_74
timestamp 1667941163
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_90
timestamp 1667941163
transform 1 0 9384 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_102
timestamp 1667941163
transform 1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_110
timestamp 1667941163
transform 1 0 11224 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1667941163
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_213
timestamp 1667941163
transform 1 0 20700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_225
timestamp 1667941163
transform 1 0 21804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_237
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1667941163
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_270
timestamp 1667941163
transform 1 0 25944 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_276
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_288
timestamp 1667941163
transform 1 0 27600 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_300
timestamp 1667941163
transform 1 0 28704 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_339
timestamp 1667941163
transform 1 0 32292 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_343
timestamp 1667941163
transform 1 0 32660 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_355
timestamp 1667941163
transform 1 0 33764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_12
timestamp 1667941163
transform 1 0 2208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_19
timestamp 1667941163
transform 1 0 2852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_32
timestamp 1667941163
transform 1 0 4048 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1667941163
transform 1 0 6808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_75
timestamp 1667941163
transform 1 0 8004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_79
timestamp 1667941163
transform 1 0 8372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_85
timestamp 1667941163
transform 1 0 8924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_95
timestamp 1667941163
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1667941163
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_124
timestamp 1667941163
transform 1 0 12512 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_136
timestamp 1667941163
transform 1 0 13616 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_148
timestamp 1667941163
transform 1 0 14720 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1667941163
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1667941163
transform 1 0 19596 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_342
timestamp 1667941163
transform 1 0 32568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_354
timestamp 1667941163
transform 1 0 33672 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_360
timestamp 1667941163
transform 1 0 34224 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_363
timestamp 1667941163
transform 1 0 34500 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_368
timestamp 1667941163
transform 1 0 34960 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_380
timestamp 1667941163
transform 1 0 36064 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_8
timestamp 1667941163
transform 1 0 1840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1667941163
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_45
timestamp 1667941163
transform 1 0 5244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_57
timestamp 1667941163
transform 1 0 6348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_61
timestamp 1667941163
transform 1 0 6716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_74
timestamp 1667941163
transform 1 0 7912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_78
timestamp 1667941163
transform 1 0 8280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1667941163
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_95
timestamp 1667941163
transform 1 0 9844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_107
timestamp 1667941163
transform 1 0 10948 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_111
timestamp 1667941163
transform 1 0 11316 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_119
timestamp 1667941163
transform 1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_125
timestamp 1667941163
transform 1 0 12604 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_131
timestamp 1667941163
transform 1 0 13156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1667941163
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_173
timestamp 1667941163
transform 1 0 17020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1667941163
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_206
timestamp 1667941163
transform 1 0 20056 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_218
timestamp 1667941163
transform 1 0 21160 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1667941163
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_10
timestamp 1667941163
transform 1 0 2024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_31
timestamp 1667941163
transform 1 0 3956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_40
timestamp 1667941163
transform 1 0 4784 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1667941163
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_67
timestamp 1667941163
transform 1 0 7268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_74
timestamp 1667941163
transform 1 0 7912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_87
timestamp 1667941163
transform 1 0 9108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_100
timestamp 1667941163
transform 1 0 10304 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1667941163
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_124
timestamp 1667941163
transform 1 0 12512 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_131
timestamp 1667941163
transform 1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_138
timestamp 1667941163
transform 1 0 13800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1667941163
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1667941163
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1667941163
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_177
timestamp 1667941163
transform 1 0 17388 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_190
timestamp 1667941163
transform 1 0 18584 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_197
timestamp 1667941163
transform 1 0 19228 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_206
timestamp 1667941163
transform 1 0 20056 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_235
timestamp 1667941163
transform 1 0 22724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_242
timestamp 1667941163
transform 1 0 23368 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_257
timestamp 1667941163
transform 1 0 24748 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_10
timestamp 1667941163
transform 1 0 2024 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_17
timestamp 1667941163
transform 1 0 2668 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1667941163
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_34
timestamp 1667941163
transform 1 0 4232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1667941163
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_95
timestamp 1667941163
transform 1 0 9844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_99
timestamp 1667941163
transform 1 0 10212 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_103
timestamp 1667941163
transform 1 0 10580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1667941163
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1667941163
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_152
timestamp 1667941163
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_212
timestamp 1667941163
transform 1 0 20608 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_216
timestamp 1667941163
transform 1 0 20976 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_220
timestamp 1667941163
transform 1 0 21344 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_232
timestamp 1667941163
transform 1 0 22448 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1667941163
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1667941163
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_264
timestamp 1667941163
transform 1 0 25392 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_272
timestamp 1667941163
transform 1 0 26128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_284
timestamp 1667941163
transform 1 0 27232 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_295
timestamp 1667941163
transform 1 0 28244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_337
timestamp 1667941163
transform 1 0 32108 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_349
timestamp 1667941163
transform 1 0 33212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1667941163
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1667941163
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1667941163
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_20
timestamp 1667941163
transform 1 0 2944 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_34
timestamp 1667941163
transform 1 0 4232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp 1667941163
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_64
timestamp 1667941163
transform 1 0 6992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_73
timestamp 1667941163
transform 1 0 7820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_83
timestamp 1667941163
transform 1 0 8740 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1667941163
transform 1 0 9476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_96
timestamp 1667941163
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1667941163
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_128
timestamp 1667941163
transform 1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_141
timestamp 1667941163
transform 1 0 14076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1667941163
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1667941163
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1667941163
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_199
timestamp 1667941163
transform 1 0 19412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1667941163
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_231
timestamp 1667941163
transform 1 0 22356 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_235
timestamp 1667941163
transform 1 0 22724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_247
timestamp 1667941163
transform 1 0 23828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_251
timestamp 1667941163
transform 1 0 24196 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_255
timestamp 1667941163
transform 1 0 24564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_262
timestamp 1667941163
transform 1 0 25208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1667941163
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1667941163
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_291
timestamp 1667941163
transform 1 0 27876 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_298
timestamp 1667941163
transform 1 0 28520 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_310
timestamp 1667941163
transform 1 0 29624 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_322
timestamp 1667941163
transform 1 0 30728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1667941163
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_12
timestamp 1667941163
transform 1 0 2208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1667941163
transform 1 0 2944 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1667941163
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_34
timestamp 1667941163
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_38
timestamp 1667941163
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_42
timestamp 1667941163
transform 1 0 4968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_49
timestamp 1667941163
transform 1 0 5612 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_56
timestamp 1667941163
transform 1 0 6256 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_68
timestamp 1667941163
transform 1 0 7360 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_100
timestamp 1667941163
transform 1 0 10304 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_125
timestamp 1667941163
transform 1 0 12604 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1667941163
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_146
timestamp 1667941163
transform 1 0 14536 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1667941163
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_159
timestamp 1667941163
transform 1 0 15732 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_173
timestamp 1667941163
transform 1 0 17020 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_184
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1667941163
transform 1 0 20884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_223
timestamp 1667941163
transform 1 0 21620 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_238
timestamp 1667941163
transform 1 0 23000 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1667941163
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_268
timestamp 1667941163
transform 1 0 25760 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_280
timestamp 1667941163
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_292
timestamp 1667941163
transform 1 0 27968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_296
timestamp 1667941163
transform 1 0 28336 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 1667941163
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_397
timestamp 1667941163
transform 1 0 37628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1667941163
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1667941163
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_16
timestamp 1667941163
transform 1 0 2576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_20
timestamp 1667941163
transform 1 0 2944 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_24
timestamp 1667941163
transform 1 0 3312 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_31
timestamp 1667941163
transform 1 0 3956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1667941163
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_64
timestamp 1667941163
transform 1 0 6992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_89
timestamp 1667941163
transform 1 0 9292 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1667941163
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1667941163
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_133
timestamp 1667941163
transform 1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_140
timestamp 1667941163
transform 1 0 13984 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_152
timestamp 1667941163
transform 1 0 15088 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1667941163
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_177
timestamp 1667941163
transform 1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_201
timestamp 1667941163
transform 1 0 19596 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_207
timestamp 1667941163
transform 1 0 20148 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1667941163
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_230
timestamp 1667941163
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_238
timestamp 1667941163
transform 1 0 23000 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_253
timestamp 1667941163
transform 1 0 24380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_265
timestamp 1667941163
transform 1 0 25484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_271
timestamp 1667941163
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1667941163
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1667941163
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1667941163
transform 1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_45
timestamp 1667941163
transform 1 0 5244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_49
timestamp 1667941163
transform 1 0 5612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_56
timestamp 1667941163
transform 1 0 6256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_69
timestamp 1667941163
transform 1 0 7452 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1667941163
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_105
timestamp 1667941163
transform 1 0 10764 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_111
timestamp 1667941163
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1667941163
transform 1 0 11684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_122
timestamp 1667941163
transform 1 0 12328 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_129
timestamp 1667941163
transform 1 0 12972 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_148
timestamp 1667941163
transform 1 0 14720 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_156
timestamp 1667941163
transform 1 0 15456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_161
timestamp 1667941163
transform 1 0 15916 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_174
timestamp 1667941163
transform 1 0 17112 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_181
timestamp 1667941163
transform 1 0 17756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1667941163
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_239
timestamp 1667941163
transform 1 0 23092 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1667941163
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_313
timestamp 1667941163
transform 1 0 29900 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_327
timestamp 1667941163
transform 1 0 31188 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_339
timestamp 1667941163
transform 1 0 32292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_351
timestamp 1667941163
transform 1 0 33396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_396
timestamp 1667941163
transform 1 0 37536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_400
timestamp 1667941163
transform 1 0 37904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_26
timestamp 1667941163
transform 1 0 3496 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_34
timestamp 1667941163
transform 1 0 4232 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_46
timestamp 1667941163
transform 1 0 5336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1667941163
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_68
timestamp 1667941163
transform 1 0 7360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_75
timestamp 1667941163
transform 1 0 8004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1667941163
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_89
timestamp 1667941163
transform 1 0 9292 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1667941163
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1667941163
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_128
timestamp 1667941163
transform 1 0 12880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1667941163
transform 1 0 13524 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_143
timestamp 1667941163
transform 1 0 14260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_185
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_195
timestamp 1667941163
transform 1 0 19044 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_203
timestamp 1667941163
transform 1 0 19780 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1667941163
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1667941163
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_256
timestamp 1667941163
transform 1 0 24656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_268
timestamp 1667941163
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_300
timestamp 1667941163
transform 1 0 28704 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_312
timestamp 1667941163
transform 1 0 29808 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_324
timestamp 1667941163
transform 1 0 30912 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_10
timestamp 1667941163
transform 1 0 2024 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1667941163
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1667941163
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_48
timestamp 1667941163
transform 1 0 5520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_55
timestamp 1667941163
transform 1 0 6164 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_59
timestamp 1667941163
transform 1 0 6532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_69
timestamp 1667941163
transform 1 0 7452 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_75
timestamp 1667941163
transform 1 0 8004 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1667941163
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_101
timestamp 1667941163
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_112
timestamp 1667941163
transform 1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_119
timestamp 1667941163
transform 1 0 12052 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1667941163
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1667941163
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_154
timestamp 1667941163
transform 1 0 15272 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_166
timestamp 1667941163
transform 1 0 16376 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_178
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_210
timestamp 1667941163
transform 1 0 20424 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_222
timestamp 1667941163
transform 1 0 21528 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_230
timestamp 1667941163
transform 1 0 22264 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_235
timestamp 1667941163
transform 1 0 22724 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_247
timestamp 1667941163
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_258
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_270
timestamp 1667941163
transform 1 0 25944 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_282
timestamp 1667941163
transform 1 0 27048 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_291
timestamp 1667941163
transform 1 0 27876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_303
timestamp 1667941163
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1667941163
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_29
timestamp 1667941163
transform 1 0 3772 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1667941163
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_68
timestamp 1667941163
transform 1 0 7360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_80
timestamp 1667941163
transform 1 0 8464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_86
timestamp 1667941163
transform 1 0 9016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_90
timestamp 1667941163
transform 1 0 9384 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_96
timestamp 1667941163
transform 1 0 9936 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1667941163
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1667941163
transform 1 0 11960 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_191
timestamp 1667941163
transform 1 0 18676 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_198
timestamp 1667941163
transform 1 0 19320 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_210
timestamp 1667941163
transform 1 0 20424 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_218
timestamp 1667941163
transform 1 0 21160 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_244
timestamp 1667941163
transform 1 0 23552 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_254
timestamp 1667941163
transform 1 0 24472 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_266
timestamp 1667941163
transform 1 0 25576 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_9
timestamp 1667941163
transform 1 0 1932 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_17
timestamp 1667941163
transform 1 0 2668 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1667941163
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_33
timestamp 1667941163
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1667941163
transform 1 0 5428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1667941163
transform 1 0 6072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_58
timestamp 1667941163
transform 1 0 6440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_62
timestamp 1667941163
transform 1 0 6808 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_68
timestamp 1667941163
transform 1 0 7360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_92
timestamp 1667941163
transform 1 0 9568 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_105
timestamp 1667941163
transform 1 0 10764 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1667941163
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1667941163
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_169
timestamp 1667941163
transform 1 0 16652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_183
timestamp 1667941163
transform 1 0 17940 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_202
timestamp 1667941163
transform 1 0 19688 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_214
timestamp 1667941163
transform 1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_220
timestamp 1667941163
transform 1 0 21344 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_232
timestamp 1667941163
transform 1 0 22448 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1667941163
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_268
timestamp 1667941163
transform 1 0 25760 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_293
timestamp 1667941163
transform 1 0 28060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1667941163
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_315
timestamp 1667941163
transform 1 0 30084 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_327
timestamp 1667941163
transform 1 0 31188 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_339
timestamp 1667941163
transform 1 0 32292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_351
timestamp 1667941163
transform 1 0 33396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_19
timestamp 1667941163
transform 1 0 2852 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_26
timestamp 1667941163
transform 1 0 3496 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_61
timestamp 1667941163
transform 1 0 6716 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_65
timestamp 1667941163
transform 1 0 7084 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_73
timestamp 1667941163
transform 1 0 7820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_79
timestamp 1667941163
transform 1 0 8372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_86
timestamp 1667941163
transform 1 0 9016 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_92
timestamp 1667941163
transform 1 0 9568 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1667941163
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_103
timestamp 1667941163
transform 1 0 10580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_128
timestamp 1667941163
transform 1 0 12880 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_139
timestamp 1667941163
transform 1 0 13892 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_151
timestamp 1667941163
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_184
timestamp 1667941163
transform 1 0 18032 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_192
timestamp 1667941163
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_203
timestamp 1667941163
transform 1 0 19780 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1667941163
transform 1 0 22264 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_247
timestamp 1667941163
transform 1 0 23828 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_259
timestamp 1667941163
transform 1 0 24932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_271
timestamp 1667941163
transform 1 0 26036 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1667941163
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_285
timestamp 1667941163
transform 1 0 27324 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_289
timestamp 1667941163
transform 1 0 27692 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_301
timestamp 1667941163
transform 1 0 28796 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_313
timestamp 1667941163
transform 1 0 29900 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_325
timestamp 1667941163
transform 1 0 31004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1667941163
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_353
timestamp 1667941163
transform 1 0 33580 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_365
timestamp 1667941163
transform 1 0 34684 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_377
timestamp 1667941163
transform 1 0 35788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1667941163
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_401
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_12
timestamp 1667941163
transform 1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_19
timestamp 1667941163
transform 1 0 2852 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1667941163
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_35
timestamp 1667941163
transform 1 0 4324 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_43
timestamp 1667941163
transform 1 0 5060 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1667941163
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_54
timestamp 1667941163
transform 1 0 6072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_61
timestamp 1667941163
transform 1 0 6716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_70
timestamp 1667941163
transform 1 0 7544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_74
timestamp 1667941163
transform 1 0 7912 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 1667941163
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1667941163
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_98
timestamp 1667941163
transform 1 0 10120 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_107
timestamp 1667941163
transform 1 0 10948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_113
timestamp 1667941163
transform 1 0 11500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_117
timestamp 1667941163
transform 1 0 11868 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_129
timestamp 1667941163
transform 1 0 12972 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1667941163
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_151
timestamp 1667941163
transform 1 0 14996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_158
timestamp 1667941163
transform 1 0 15640 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_166
timestamp 1667941163
transform 1 0 16376 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1667941163
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185
timestamp 1667941163
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1667941163
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_217
timestamp 1667941163
transform 1 0 21068 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_222
timestamp 1667941163
transform 1 0 21528 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_234
timestamp 1667941163
transform 1 0 22632 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1667941163
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_393
timestamp 1667941163
transform 1 0 37260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_397
timestamp 1667941163
transform 1 0 37628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1667941163
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_16
timestamp 1667941163
transform 1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_20
timestamp 1667941163
transform 1 0 2944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_24
timestamp 1667941163
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_31
timestamp 1667941163
transform 1 0 3956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_38
timestamp 1667941163
transform 1 0 4600 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_46
timestamp 1667941163
transform 1 0 5336 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1667941163
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_89
timestamp 1667941163
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_128
timestamp 1667941163
transform 1 0 12880 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_136
timestamp 1667941163
transform 1 0 13616 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_142
timestamp 1667941163
transform 1 0 14168 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_154
timestamp 1667941163
transform 1 0 15272 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1667941163
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_177
timestamp 1667941163
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_183
timestamp 1667941163
transform 1 0 17940 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_190
timestamp 1667941163
transform 1 0 18584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_197
timestamp 1667941163
transform 1 0 19228 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_201
timestamp 1667941163
transform 1 0 19596 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_211
timestamp 1667941163
transform 1 0 20516 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_215
timestamp 1667941163
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_301
timestamp 1667941163
transform 1 0 28796 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_307
timestamp 1667941163
transform 1 0 29348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_319
timestamp 1667941163
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1667941163
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_400
timestamp 1667941163
transform 1 0 37904 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_406
timestamp 1667941163
transform 1 0 38456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_8
timestamp 1667941163
transform 1 0 1840 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_51
timestamp 1667941163
transform 1 0 5796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1667941163
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1667941163
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_185
timestamp 1667941163
transform 1 0 18124 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1667941163
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_234
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1667941163
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_30
timestamp 1667941163
transform 1 0 3864 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1667941163
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_62
timestamp 1667941163
transform 1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_66
timestamp 1667941163
transform 1 0 7176 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_90
timestamp 1667941163
transform 1 0 9384 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_102
timestamp 1667941163
transform 1 0 10488 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_118
timestamp 1667941163
transform 1 0 11960 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_130
timestamp 1667941163
transform 1 0 13064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_134
timestamp 1667941163
transform 1 0 13432 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_155
timestamp 1667941163
transform 1 0 15364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_191
timestamp 1667941163
transform 1 0 18676 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_210
timestamp 1667941163
transform 1 0 20424 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_214
timestamp 1667941163
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_235
timestamp 1667941163
transform 1 0 22724 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_242
timestamp 1667941163
transform 1 0 23368 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_260
timestamp 1667941163
transform 1 0 25024 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1667941163
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_401
timestamp 1667941163
transform 1 0 37996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1667941163
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_37
timestamp 1667941163
transform 1 0 4508 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1667941163
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_105
timestamp 1667941163
transform 1 0 10764 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_128
timestamp 1667941163
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_147
timestamp 1667941163
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_171
timestamp 1667941163
transform 1 0 16836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_183
timestamp 1667941163
transform 1 0 17940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_202
timestamp 1667941163
transform 1 0 19688 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_214
timestamp 1667941163
transform 1 0 20792 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_226
timestamp 1667941163
transform 1 0 21896 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_236
timestamp 1667941163
transform 1 0 22816 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_243
timestamp 1667941163
transform 1 0 23460 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1667941163
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1667941163
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_271
timestamp 1667941163
transform 1 0 26036 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_283
timestamp 1667941163
transform 1 0 27140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_295
timestamp 1667941163
transform 1 0 28244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_313
timestamp 1667941163
transform 1 0 29900 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_317
timestamp 1667941163
transform 1 0 30268 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_329
timestamp 1667941163
transform 1 0 31372 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_341
timestamp 1667941163
transform 1 0 32476 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_353
timestamp 1667941163
transform 1 0 33580 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1667941163
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_25
timestamp 1667941163
transform 1 0 3404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_33
timestamp 1667941163
transform 1 0 4140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_98
timestamp 1667941163
transform 1 0 10120 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1667941163
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_192
timestamp 1667941163
transform 1 0 18768 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_204
timestamp 1667941163
transform 1 0 19872 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_208
timestamp 1667941163
transform 1 0 20240 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_212
timestamp 1667941163
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1667941163
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_240
timestamp 1667941163
transform 1 0 23184 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_252
timestamp 1667941163
transform 1 0 24288 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_259
timestamp 1667941163
transform 1 0 24932 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_271
timestamp 1667941163
transform 1 0 26036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_314
timestamp 1667941163
transform 1 0 29992 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_327
timestamp 1667941163
transform 1 0 31188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_401
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_52
timestamp 1667941163
transform 1 0 5888 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1667941163
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_124
timestamp 1667941163
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_134
timestamp 1667941163
transform 1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1667941163
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_262
timestamp 1667941163
transform 1 0 25208 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_270
timestamp 1667941163
transform 1 0 25944 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_284
timestamp 1667941163
transform 1 0 27232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_292
timestamp 1667941163
transform 1 0 27968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_299
timestamp 1667941163
transform 1 0 28612 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1667941163
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_9
timestamp 1667941163
transform 1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_13
timestamp 1667941163
transform 1 0 2300 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_35
timestamp 1667941163
transform 1 0 4324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_47
timestamp 1667941163
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_83
timestamp 1667941163
transform 1 0 8740 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1667941163
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_132
timestamp 1667941163
transform 1 0 13248 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1667941163
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1667941163
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_174
timestamp 1667941163
transform 1 0 17112 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_186
timestamp 1667941163
transform 1 0 18216 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_194
timestamp 1667941163
transform 1 0 18952 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_198
timestamp 1667941163
transform 1 0 19320 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_210
timestamp 1667941163
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1667941163
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1667941163
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_253
timestamp 1667941163
transform 1 0 24380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_260
timestamp 1667941163
transform 1 0 25024 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1667941163
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_297
timestamp 1667941163
transform 1 0 28428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp 1667941163
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_321
timestamp 1667941163
transform 1 0 30636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1667941163
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp 1667941163
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_37
timestamp 1667941163
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_58
timestamp 1667941163
transform 1 0 6440 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1667941163
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_103
timestamp 1667941163
transform 1 0 10580 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_127
timestamp 1667941163
transform 1 0 12788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_182
timestamp 1667941163
transform 1 0 17848 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_201
timestamp 1667941163
transform 1 0 19596 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_215
timestamp 1667941163
transform 1 0 20884 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_227
timestamp 1667941163
transform 1 0 21988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_239
timestamp 1667941163
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1667941163
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_286
timestamp 1667941163
transform 1 0 27416 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1667941163
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_314
timestamp 1667941163
transform 1 0 29992 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1667941163
transform 1 0 1840 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_20
timestamp 1667941163
transform 1 0 2944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_28
timestamp 1667941163
transform 1 0 3680 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1667941163
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_117
timestamp 1667941163
transform 1 0 11868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp 1667941163
transform 1 0 13800 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_153
timestamp 1667941163
transform 1 0 15180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1667941163
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_192
timestamp 1667941163
transform 1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_199
timestamp 1667941163
transform 1 0 19412 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_208
timestamp 1667941163
transform 1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_212
timestamp 1667941163
transform 1 0 20608 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1667941163
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1667941163
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_245
timestamp 1667941163
transform 1 0 23644 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_257
timestamp 1667941163
transform 1 0 24748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_269
timestamp 1667941163
transform 1 0 25852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 1667941163
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_289
timestamp 1667941163
transform 1 0 27692 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_299
timestamp 1667941163
transform 1 0 28612 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_311
timestamp 1667941163
transform 1 0 29716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_323
timestamp 1667941163
transform 1 0 30820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_401
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_9
timestamp 1667941163
transform 1 0 1932 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1667941163
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_51
timestamp 1667941163
transform 1 0 5796 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_59
timestamp 1667941163
transform 1 0 6532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_102
timestamp 1667941163
transform 1 0 10488 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_114
timestamp 1667941163
transform 1 0 11592 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_126
timestamp 1667941163
transform 1 0 12696 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_149
timestamp 1667941163
transform 1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_173
timestamp 1667941163
transform 1 0 17020 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_185
timestamp 1667941163
transform 1 0 18124 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1667941163
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_202
timestamp 1667941163
transform 1 0 19688 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_214
timestamp 1667941163
transform 1 0 20792 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_222
timestamp 1667941163
transform 1 0 21528 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_228
timestamp 1667941163
transform 1 0 22080 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_240
timestamp 1667941163
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_281
timestamp 1667941163
transform 1 0 26956 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1667941163
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_295
timestamp 1667941163
transform 1 0 28244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_314
timestamp 1667941163
transform 1 0 29992 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_326
timestamp 1667941163
transform 1 0 31096 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_338
timestamp 1667941163
transform 1 0 32200 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_350
timestamp 1667941163
transform 1 0 33304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_28
timestamp 1667941163
transform 1 0 3680 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_40
timestamp 1667941163
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1667941163
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_144
timestamp 1667941163
transform 1 0 14352 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_156
timestamp 1667941163
transform 1 0 15456 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_189
timestamp 1667941163
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_260
timestamp 1667941163
transform 1 0 25024 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_264
timestamp 1667941163
transform 1 0 25392 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_286
timestamp 1667941163
transform 1 0 27416 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_298
timestamp 1667941163
transform 1 0 28520 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_310
timestamp 1667941163
transform 1 0 29624 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_322
timestamp 1667941163
transform 1 0 30728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1667941163
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_382
timestamp 1667941163
transform 1 0 36248 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1667941163
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_7
timestamp 1667941163
transform 1 0 1748 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_11
timestamp 1667941163
transform 1 0 2116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1667941163
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_48
timestamp 1667941163
transform 1 0 5520 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_63
timestamp 1667941163
transform 1 0 6900 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_70
timestamp 1667941163
transform 1 0 7544 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_122
timestamp 1667941163
transform 1 0 12328 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_128
timestamp 1667941163
transform 1 0 12880 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_163
timestamp 1667941163
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_175
timestamp 1667941163
transform 1 0 17204 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_214
timestamp 1667941163
transform 1 0 20792 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_220
timestamp 1667941163
transform 1 0 21344 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_224
timestamp 1667941163
transform 1 0 21712 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_232
timestamp 1667941163
transform 1 0 22448 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1667941163
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1667941163
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1667941163
transform 1 0 26036 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_278
timestamp 1667941163
transform 1 0 26680 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_290
timestamp 1667941163
transform 1 0 27784 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1667941163
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_314
timestamp 1667941163
transform 1 0 29992 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_322
timestamp 1667941163
transform 1 0 30728 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_338
timestamp 1667941163
transform 1 0 32200 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_350
timestamp 1667941163
transform 1 0 33304 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1667941163
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_397
timestamp 1667941163
transform 1 0 37628 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_402
timestamp 1667941163
transform 1 0 38088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1667941163
transform 1 0 38456 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_10
timestamp 1667941163
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_35
timestamp 1667941163
transform 1 0 4324 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_43
timestamp 1667941163
transform 1 0 5060 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_48
timestamp 1667941163
transform 1 0 5520 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_62
timestamp 1667941163
transform 1 0 6808 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_68
timestamp 1667941163
transform 1 0 7360 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_89
timestamp 1667941163
transform 1 0 9292 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_101
timestamp 1667941163
transform 1 0 10396 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1667941163
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_124
timestamp 1667941163
transform 1 0 12512 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_152
timestamp 1667941163
transform 1 0 15088 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1667941163
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_191
timestamp 1667941163
transform 1 0 18676 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_203
timestamp 1667941163
transform 1 0 19780 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_244
timestamp 1667941163
transform 1 0 23552 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_251
timestamp 1667941163
transform 1 0 24196 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_257
timestamp 1667941163
transform 1 0 24748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_266
timestamp 1667941163
transform 1 0 25576 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_325
timestamp 1667941163
transform 1 0 31004 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_330
timestamp 1667941163
transform 1 0 31464 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_13
timestamp 1667941163
transform 1 0 2300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1667941163
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_35
timestamp 1667941163
transform 1 0 4324 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_39
timestamp 1667941163
transform 1 0 4692 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_63
timestamp 1667941163
transform 1 0 6900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_75
timestamp 1667941163
transform 1 0 8004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_98
timestamp 1667941163
transform 1 0 10120 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_110
timestamp 1667941163
transform 1 0 11224 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_122
timestamp 1667941163
transform 1 0 12328 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1667941163
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_187
timestamp 1667941163
transform 1 0 18308 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_208
timestamp 1667941163
transform 1 0 20240 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_228
timestamp 1667941163
transform 1 0 22080 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_235
timestamp 1667941163
transform 1 0 22724 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_242
timestamp 1667941163
transform 1 0 23368 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1667941163
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_268
timestamp 1667941163
transform 1 0 25760 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_275
timestamp 1667941163
transform 1 0 26404 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_282
timestamp 1667941163
transform 1 0 27048 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_294
timestamp 1667941163
transform 1 0 28152 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1667941163
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_8
timestamp 1667941163
transform 1 0 1840 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_20
timestamp 1667941163
transform 1 0 2944 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_26
timestamp 1667941163
transform 1 0 3496 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1667941163
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_131
timestamp 1667941163
transform 1 0 13156 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_152
timestamp 1667941163
transform 1 0 15088 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1667941163
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_182
timestamp 1667941163
transform 1 0 17848 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_186
timestamp 1667941163
transform 1 0 18216 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_190
timestamp 1667941163
transform 1 0 18584 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_197
timestamp 1667941163
transform 1 0 19228 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_204
timestamp 1667941163
transform 1 0 19872 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1667941163
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_230
timestamp 1667941163
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_245
timestamp 1667941163
transform 1 0 23644 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_260
timestamp 1667941163
transform 1 0 25024 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_264
timestamp 1667941163
transform 1 0 25392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_286
timestamp 1667941163
transform 1 0 27416 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_295
timestamp 1667941163
transform 1 0 28244 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_306
timestamp 1667941163
transform 1 0 29256 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_318
timestamp 1667941163
transform 1 0 30360 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1667941163
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_9
timestamp 1667941163
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1667941163
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_44
timestamp 1667941163
transform 1 0 5152 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_52
timestamp 1667941163
transform 1 0 5888 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1667941163
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_147
timestamp 1667941163
transform 1 0 14628 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_168
timestamp 1667941163
transform 1 0 16560 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_180
timestamp 1667941163
transform 1 0 17664 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_187
timestamp 1667941163
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_202
timestamp 1667941163
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_219
timestamp 1667941163
transform 1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_226
timestamp 1667941163
transform 1 0 21896 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_240
timestamp 1667941163
transform 1 0 23184 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1667941163
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_264
timestamp 1667941163
transform 1 0 25392 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1667941163
transform 1 0 26036 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_278
timestamp 1667941163
transform 1 0 26680 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_285
timestamp 1667941163
transform 1 0 27324 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1667941163
transform 1 0 28060 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_297
timestamp 1667941163
transform 1 0 28428 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1667941163
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_316
timestamp 1667941163
transform 1 0 30176 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_328
timestamp 1667941163
transform 1 0 31280 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_23
timestamp 1667941163
transform 1 0 3220 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_29
timestamp 1667941163
transform 1 0 3772 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1667941163
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_85
timestamp 1667941163
transform 1 0 8924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 1667941163
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_144
timestamp 1667941163
transform 1 0 14352 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_156
timestamp 1667941163
transform 1 0 15456 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_191
timestamp 1667941163
transform 1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_198
timestamp 1667941163
transform 1 0 19320 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_229
timestamp 1667941163
transform 1 0 22172 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_251
timestamp 1667941163
transform 1 0 24196 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_268
timestamp 1667941163
transform 1 0 25760 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1667941163
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_299
timestamp 1667941163
transform 1 0 28612 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_303
timestamp 1667941163
transform 1 0 28980 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_324
timestamp 1667941163
transform 1 0 30912 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_11
timestamp 1667941163
transform 1 0 2116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1667941163
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_120
timestamp 1667941163
transform 1 0 12144 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_132
timestamp 1667941163
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_191
timestamp 1667941163
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_202
timestamp 1667941163
transform 1 0 19688 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_208
timestamp 1667941163
transform 1 0 20240 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_212
timestamp 1667941163
transform 1 0 20608 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_219
timestamp 1667941163
transform 1 0 21252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_226
timestamp 1667941163
transform 1 0 21896 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_237
timestamp 1667941163
transform 1 0 22908 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_244
timestamp 1667941163
transform 1 0 23552 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_258
timestamp 1667941163
transform 1 0 24840 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_281
timestamp 1667941163
transform 1 0 26956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_293
timestamp 1667941163
transform 1 0 28060 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_297
timestamp 1667941163
transform 1 0 28428 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1667941163
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_314
timestamp 1667941163
transform 1 0 29992 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_326
timestamp 1667941163
transform 1 0 31096 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_338
timestamp 1667941163
transform 1 0 32200 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_350
timestamp 1667941163
transform 1 0 33304 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1667941163
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_21
timestamp 1667941163
transform 1 0 3036 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1667941163
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1667941163
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_138
timestamp 1667941163
transform 1 0 13800 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_145
timestamp 1667941163
transform 1 0 14444 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_157
timestamp 1667941163
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1667941163
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_191
timestamp 1667941163
transform 1 0 18676 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_201
timestamp 1667941163
transform 1 0 19596 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_208
timestamp 1667941163
transform 1 0 20240 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1667941163
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_248
timestamp 1667941163
transform 1 0 23920 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1667941163
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_272
timestamp 1667941163
transform 1 0 26128 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_296
timestamp 1667941163
transform 1 0 28336 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_308
timestamp 1667941163
transform 1 0 29440 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_320
timestamp 1667941163
transform 1 0 30544 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_328
timestamp 1667941163
transform 1 0 31280 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_333
timestamp 1667941163
transform 1 0 31740 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_402
timestamp 1667941163
transform 1 0 38088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_406
timestamp 1667941163
transform 1 0 38456 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1667941163
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_35
timestamp 1667941163
transform 1 0 4324 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_39
timestamp 1667941163
transform 1 0 4692 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_51
timestamp 1667941163
transform 1 0 5796 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_63
timestamp 1667941163
transform 1 0 6900 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_75
timestamp 1667941163
transform 1 0 8004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_119
timestamp 1667941163
transform 1 0 12052 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_131
timestamp 1667941163
transform 1 0 13156 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_159
timestamp 1667941163
transform 1 0 15732 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_183
timestamp 1667941163
transform 1 0 17940 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_190
timestamp 1667941163
transform 1 0 18584 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_238
timestamp 1667941163
transform 1 0 23000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1667941163
transform 1 0 24840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_272
timestamp 1667941163
transform 1 0 26128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_279
timestamp 1667941163
transform 1 0 26772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_286
timestamp 1667941163
transform 1 0 27416 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_293
timestamp 1667941163
transform 1 0 28060 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_300
timestamp 1667941163
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_314
timestamp 1667941163
transform 1 0 29992 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_339
timestamp 1667941163
transform 1 0 32292 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_343
timestamp 1667941163
transform 1 0 32660 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_355
timestamp 1667941163
transform 1 0 33764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1667941163
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_20
timestamp 1667941163
transform 1 0 2944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_28
timestamp 1667941163
transform 1 0 3680 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1667941163
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_97
timestamp 1667941163
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1667941163
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_147
timestamp 1667941163
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1667941163
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_191
timestamp 1667941163
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_198
timestamp 1667941163
transform 1 0 19320 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_210
timestamp 1667941163
transform 1 0 20424 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_214
timestamp 1667941163
transform 1 0 20792 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_218
timestamp 1667941163
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_240
timestamp 1667941163
transform 1 0 23184 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_253
timestamp 1667941163
transform 1 0 24380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_260
timestamp 1667941163
transform 1 0 25024 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_264
timestamp 1667941163
transform 1 0 25392 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1667941163
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_292
timestamp 1667941163
transform 1 0 27968 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_299
timestamp 1667941163
transform 1 0 28612 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_306
timestamp 1667941163
transform 1 0 29256 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_318
timestamp 1667941163
transform 1 0 30360 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1667941163
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_7
timestamp 1667941163
transform 1 0 1748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_11
timestamp 1667941163
transform 1 0 2116 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_17
timestamp 1667941163
transform 1 0 2668 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1667941163
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_66
timestamp 1667941163
transform 1 0 7176 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_78
timestamp 1667941163
transform 1 0 8280 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_131
timestamp 1667941163
transform 1 0 13156 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1667941163
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_146
timestamp 1667941163
transform 1 0 14536 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_152
timestamp 1667941163
transform 1 0 15088 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_174
timestamp 1667941163
transform 1 0 17112 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1667941163
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_218
timestamp 1667941163
transform 1 0 21160 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_225
timestamp 1667941163
transform 1 0 21804 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1667941163
transform 1 0 22448 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_236
timestamp 1667941163
transform 1 0 22816 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1667941163
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_258
timestamp 1667941163
transform 1 0 24840 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_266
timestamp 1667941163
transform 1 0 25576 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_285
timestamp 1667941163
transform 1 0 27324 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_295
timestamp 1667941163
transform 1 0 28244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1667941163
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_314
timestamp 1667941163
transform 1 0 29992 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_326
timestamp 1667941163
transform 1 0 31096 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_331
timestamp 1667941163
transform 1 0 31556 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_343
timestamp 1667941163
transform 1 0 32660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_355
timestamp 1667941163
transform 1 0 33764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_20
timestamp 1667941163
transform 1 0 2944 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_26
timestamp 1667941163
transform 1 0 3496 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_38
timestamp 1667941163
transform 1 0 4600 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_50
timestamp 1667941163
transform 1 0 5704 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_80
timestamp 1667941163
transform 1 0 8464 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_87
timestamp 1667941163
transform 1 0 9108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_94
timestamp 1667941163
transform 1 0 9752 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_98
timestamp 1667941163
transform 1 0 10120 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1667941163
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_138
timestamp 1667941163
transform 1 0 13800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_142
timestamp 1667941163
transform 1 0 14168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_163
timestamp 1667941163
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_191
timestamp 1667941163
transform 1 0 18676 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_203
timestamp 1667941163
transform 1 0 19780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1667941163
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_233
timestamp 1667941163
transform 1 0 22540 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_241
timestamp 1667941163
transform 1 0 23276 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_256
timestamp 1667941163
transform 1 0 24656 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_264
timestamp 1667941163
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_275
timestamp 1667941163
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_291
timestamp 1667941163
transform 1 0 27876 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_303
timestamp 1667941163
transform 1 0 28980 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_315
timestamp 1667941163
transform 1 0 30084 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_319
timestamp 1667941163
transform 1 0 30452 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_323
timestamp 1667941163
transform 1 0 30820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_8
timestamp 1667941163
transform 1 0 1840 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1667941163
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_113
timestamp 1667941163
transform 1 0 11500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1667941163
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_186
timestamp 1667941163
transform 1 0 18216 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_190
timestamp 1667941163
transform 1 0 18584 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1667941163
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_203
timestamp 1667941163
transform 1 0 19780 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_207
timestamp 1667941163
transform 1 0 20148 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_211
timestamp 1667941163
transform 1 0 20516 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_218
timestamp 1667941163
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_235
timestamp 1667941163
transform 1 0 22724 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_242
timestamp 1667941163
transform 1 0 23368 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1667941163
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_268
timestamp 1667941163
transform 1 0 25760 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_278
timestamp 1667941163
transform 1 0 26680 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_286
timestamp 1667941163
transform 1 0 27416 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_300
timestamp 1667941163
transform 1 0 28704 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_9
timestamp 1667941163
transform 1 0 1932 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_13
timestamp 1667941163
transform 1 0 2300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_25
timestamp 1667941163
transform 1 0 3404 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_37
timestamp 1667941163
transform 1 0 4508 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 1667941163
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_135
timestamp 1667941163
transform 1 0 13524 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_147
timestamp 1667941163
transform 1 0 14628 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_159
timestamp 1667941163
transform 1 0 15732 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_192
timestamp 1667941163
transform 1 0 18768 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_200
timestamp 1667941163
transform 1 0 19504 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_213
timestamp 1667941163
transform 1 0 20700 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_240
timestamp 1667941163
transform 1 0 23184 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_257
timestamp 1667941163
transform 1 0 24748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_264
timestamp 1667941163
transform 1 0 25392 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_268
timestamp 1667941163
transform 1 0 25760 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1667941163
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_287
timestamp 1667941163
transform 1 0 27508 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_296
timestamp 1667941163
transform 1 0 28336 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_303
timestamp 1667941163
transform 1 0 28980 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_310
timestamp 1667941163
transform 1 0 29624 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_322
timestamp 1667941163
transform 1 0 30728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1667941163
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_163
timestamp 1667941163
transform 1 0 16100 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_175
timestamp 1667941163
transform 1 0 17204 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_187
timestamp 1667941163
transform 1 0 18308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_201
timestamp 1667941163
transform 1 0 19596 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_205
timestamp 1667941163
transform 1 0 19964 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_218
timestamp 1667941163
transform 1 0 21160 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_228
timestamp 1667941163
transform 1 0 22080 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_234
timestamp 1667941163
transform 1 0 22632 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_241
timestamp 1667941163
transform 1 0 23276 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1667941163
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_258
timestamp 1667941163
transform 1 0 24840 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_273
timestamp 1667941163
transform 1 0 26220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_280
timestamp 1667941163
transform 1 0 26864 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_287
timestamp 1667941163
transform 1 0 27508 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_294
timestamp 1667941163
transform 1 0 28152 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_320
timestamp 1667941163
transform 1 0 30544 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_332
timestamp 1667941163
transform 1 0 31648 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_344
timestamp 1667941163
transform 1 0 32752 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 1667941163
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_370
timestamp 1667941163
transform 1 0 35144 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_382
timestamp 1667941163
transform 1 0 36248 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_394
timestamp 1667941163
transform 1 0 37352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_8
timestamp 1667941163
transform 1 0 1840 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_20
timestamp 1667941163
transform 1 0 2944 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1667941163
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_64
timestamp 1667941163
transform 1 0 6992 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_96
timestamp 1667941163
transform 1 0 9936 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1667941163
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_142
timestamp 1667941163
transform 1 0 14168 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_154
timestamp 1667941163
transform 1 0 15272 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1667941163
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_191
timestamp 1667941163
transform 1 0 18676 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_203
timestamp 1667941163
transform 1 0 19780 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_209
timestamp 1667941163
transform 1 0 20332 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_213
timestamp 1667941163
transform 1 0 20700 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1667941163
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_241
timestamp 1667941163
transform 1 0 23276 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_248
timestamp 1667941163
transform 1 0 23920 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_255
timestamp 1667941163
transform 1 0 24564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_262
timestamp 1667941163
transform 1 0 25208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_269
timestamp 1667941163
transform 1 0 25852 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1667941163
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_286
timestamp 1667941163
transform 1 0 27416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_300
timestamp 1667941163
transform 1 0 28704 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_307
timestamp 1667941163
transform 1 0 29348 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_316
timestamp 1667941163
transform 1 0 30176 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_328
timestamp 1667941163
transform 1 0 31280 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_7
timestamp 1667941163
transform 1 0 1748 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_11
timestamp 1667941163
transform 1 0 2116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_19
timestamp 1667941163
transform 1 0 2852 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_23
timestamp 1667941163
transform 1 0 3220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_34
timestamp 1667941163
transform 1 0 4232 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_42
timestamp 1667941163
transform 1 0 4968 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_66
timestamp 1667941163
transform 1 0 7176 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_73
timestamp 1667941163
transform 1 0 7820 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_81
timestamp 1667941163
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_111
timestamp 1667941163
transform 1 0 11316 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_115
timestamp 1667941163
transform 1 0 11684 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_137
timestamp 1667941163
transform 1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_169
timestamp 1667941163
transform 1 0 16652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1667941163
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_225
timestamp 1667941163
transform 1 0 21804 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_244
timestamp 1667941163
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_258
timestamp 1667941163
transform 1 0 24840 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_272
timestamp 1667941163
transform 1 0 26128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_287
timestamp 1667941163
transform 1 0 27508 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1667941163
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_16
timestamp 1667941163
transform 1 0 2576 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_28
timestamp 1667941163
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_40
timestamp 1667941163
transform 1 0 4784 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_48
timestamp 1667941163
transform 1 0 5520 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1667941163
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_71
timestamp 1667941163
transform 1 0 7636 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_83
timestamp 1667941163
transform 1 0 8740 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_131
timestamp 1667941163
transform 1 0 13156 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_155
timestamp 1667941163
transform 1 0 15364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_191
timestamp 1667941163
transform 1 0 18676 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_199
timestamp 1667941163
transform 1 0 19412 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_212
timestamp 1667941163
transform 1 0 20608 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 1667941163
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_230
timestamp 1667941163
transform 1 0 22264 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_238
timestamp 1667941163
transform 1 0 23000 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_252
timestamp 1667941163
transform 1 0 24288 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_269
timestamp 1667941163
transform 1 0 25852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1667941163
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_286
timestamp 1667941163
transform 1 0 27416 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_401
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_25
timestamp 1667941163
transform 1 0 3404 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_40
timestamp 1667941163
transform 1 0 4784 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_46
timestamp 1667941163
transform 1 0 5336 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_56
timestamp 1667941163
transform 1 0 6256 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_63
timestamp 1667941163
transform 1 0 6900 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_70
timestamp 1667941163
transform 1 0 7544 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1667941163
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_116
timestamp 1667941163
transform 1 0 11776 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_128
timestamp 1667941163
transform 1 0 12880 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_146
timestamp 1667941163
transform 1 0 14536 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_152
timestamp 1667941163
transform 1 0 15088 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_164
timestamp 1667941163
transform 1 0 16192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_170
timestamp 1667941163
transform 1 0 16744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1667941163
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_212
timestamp 1667941163
transform 1 0 20608 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_229
timestamp 1667941163
transform 1 0 22172 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_236
timestamp 1667941163
transform 1 0 22816 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_243
timestamp 1667941163
transform 1 0 23460 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1667941163
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_264
timestamp 1667941163
transform 1 0 25392 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_270
timestamp 1667941163
transform 1 0 25944 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_280
timestamp 1667941163
transform 1 0 26864 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_297
timestamp 1667941163
transform 1 0 28428 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1667941163
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_9
timestamp 1667941163
transform 1 0 1932 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_35
timestamp 1667941163
transform 1 0 4324 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_41
timestamp 1667941163
transform 1 0 4876 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_45
timestamp 1667941163
transform 1 0 5244 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1667941163
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_92
timestamp 1667941163
transform 1 0 9568 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_104
timestamp 1667941163
transform 1 0 10672 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_118
timestamp 1667941163
transform 1 0 11960 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_130
timestamp 1667941163
transform 1 0 13064 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_152
timestamp 1667941163
transform 1 0 15088 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1667941163
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_192
timestamp 1667941163
transform 1 0 18768 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_204
timestamp 1667941163
transform 1 0 19872 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1667941163
transform 1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_230
timestamp 1667941163
transform 1 0 22264 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_241
timestamp 1667941163
transform 1 0 23276 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_245
timestamp 1667941163
transform 1 0 23644 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_252
timestamp 1667941163
transform 1 0 24288 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_271
timestamp 1667941163
transform 1 0 26036 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1667941163
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1667941163
transform 1 0 27416 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_310
timestamp 1667941163
transform 1 0 29624 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_322
timestamp 1667941163
transform 1 0 30728 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1667941163
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_34
timestamp 1667941163
transform 1 0 4232 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_46
timestamp 1667941163
transform 1 0 5336 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_58
timestamp 1667941163
transform 1 0 6440 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1667941163
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_114
timestamp 1667941163
transform 1 0 11592 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1667941163
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_154
timestamp 1667941163
transform 1 0 15272 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_160
timestamp 1667941163
transform 1 0 15824 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_181
timestamp 1667941163
transform 1 0 17756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1667941163
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_227
timestamp 1667941163
transform 1 0 21988 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_231
timestamp 1667941163
transform 1 0 22356 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_239
timestamp 1667941163
transform 1 0 23092 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1667941163
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_264
timestamp 1667941163
transform 1 0 25392 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_271
timestamp 1667941163
transform 1 0 26036 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_275
timestamp 1667941163
transform 1 0 26404 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_285
timestamp 1667941163
transform 1 0 27324 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_298
timestamp 1667941163
transform 1 0 28520 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1667941163
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_314
timestamp 1667941163
transform 1 0 29992 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_397
timestamp 1667941163
transform 1 0 37628 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_402
timestamp 1667941163
transform 1 0 38088 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1667941163
transform 1 0 38456 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_8
timestamp 1667941163
transform 1 0 1840 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_47
timestamp 1667941163
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_62
timestamp 1667941163
transform 1 0 6808 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_74
timestamp 1667941163
transform 1 0 7912 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_79
timestamp 1667941163
transform 1 0 8372 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_91
timestamp 1667941163
transform 1 0 9476 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_103
timestamp 1667941163
transform 1 0 10580 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_118
timestamp 1667941163
transform 1 0 11960 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_124
timestamp 1667941163
transform 1 0 12512 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_128
timestamp 1667941163
transform 1 0 12880 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_136
timestamp 1667941163
transform 1 0 13616 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_158
timestamp 1667941163
transform 1 0 15640 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1667941163
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_191
timestamp 1667941163
transform 1 0 18676 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_203
timestamp 1667941163
transform 1 0 19780 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_211
timestamp 1667941163
transform 1 0 20516 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1667941163
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_234
timestamp 1667941163
transform 1 0 22632 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_241
timestamp 1667941163
transform 1 0 23276 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_248
timestamp 1667941163
transform 1 0 23920 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_255
timestamp 1667941163
transform 1 0 24564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_262
timestamp 1667941163
transform 1 0 25208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_269
timestamp 1667941163
transform 1 0 25852 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1667941163
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_286
timestamp 1667941163
transform 1 0 27416 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_300
timestamp 1667941163
transform 1 0 28704 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_307
timestamp 1667941163
transform 1 0 29348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_314
timestamp 1667941163
transform 1 0 29992 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_321
timestamp 1667941163
transform 1 0 30636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1667941163
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_25
timestamp 1667941163
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_34
timestamp 1667941163
transform 1 0 4232 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_46
timestamp 1667941163
transform 1 0 5336 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_52
timestamp 1667941163
transform 1 0 5888 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_73
timestamp 1667941163
transform 1 0 7820 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_81
timestamp 1667941163
transform 1 0 8556 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_103
timestamp 1667941163
transform 1 0 10580 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_128
timestamp 1667941163
transform 1 0 12880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_135
timestamp 1667941163
transform 1 0 13524 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_167
timestamp 1667941163
transform 1 0 16468 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 1667941163
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_202
timestamp 1667941163
transform 1 0 19688 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_206
timestamp 1667941163
transform 1 0 20056 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_210
timestamp 1667941163
transform 1 0 20424 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_217
timestamp 1667941163
transform 1 0 21068 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_224
timestamp 1667941163
transform 1 0 21712 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1667941163
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_238
timestamp 1667941163
transform 1 0 23000 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_244
timestamp 1667941163
transform 1 0 23552 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1667941163
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_258
timestamp 1667941163
transform 1 0 24840 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_271
timestamp 1667941163
transform 1 0 26036 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_285
timestamp 1667941163
transform 1 0 27324 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_298
timestamp 1667941163
transform 1 0 28520 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1667941163
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_314
timestamp 1667941163
transform 1 0 29992 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_328
timestamp 1667941163
transform 1 0 31280 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_340
timestamp 1667941163
transform 1 0 32384 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_352
timestamp 1667941163
transform 1 0 33488 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_397
timestamp 1667941163
transform 1 0 37628 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1667941163
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_9
timestamp 1667941163
transform 1 0 1932 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_19
timestamp 1667941163
transform 1 0 2852 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_28
timestamp 1667941163
transform 1 0 3680 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_40
timestamp 1667941163
transform 1 0 4784 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1667941163
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_85
timestamp 1667941163
transform 1 0 8924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_90
timestamp 1667941163
transform 1 0 9384 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_102
timestamp 1667941163
transform 1 0 10488 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_109
timestamp 1667941163
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_121
timestamp 1667941163
transform 1 0 12236 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_144
timestamp 1667941163
transform 1 0 14352 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_156
timestamp 1667941163
transform 1 0 15456 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_191
timestamp 1667941163
transform 1 0 18676 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_202
timestamp 1667941163
transform 1 0 19688 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_209
timestamp 1667941163
transform 1 0 20332 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_216
timestamp 1667941163
transform 1 0 20976 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1667941163
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_242
timestamp 1667941163
transform 1 0 23368 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_268
timestamp 1667941163
transform 1 0 25760 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_275
timestamp 1667941163
transform 1 0 26404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_286
timestamp 1667941163
transform 1 0 27416 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_299
timestamp 1667941163
transform 1 0 28612 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_312
timestamp 1667941163
transform 1 0 29808 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_319
timestamp 1667941163
transform 1 0 30452 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_326
timestamp 1667941163
transform 1 0 31096 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1667941163
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_342
timestamp 1667941163
transform 1 0 32568 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_354
timestamp 1667941163
transform 1 0 33672 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_366
timestamp 1667941163
transform 1 0 34776 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_378
timestamp 1667941163
transform 1 0 35880 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1667941163
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_70
timestamp 1667941163
transform 1 0 7544 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_78
timestamp 1667941163
transform 1 0 8280 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1667941163
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_116
timestamp 1667941163
transform 1 0 11776 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_131
timestamp 1667941163
transform 1 0 13156 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1667941163
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1667941163
transform 1 0 14444 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_149
timestamp 1667941163
transform 1 0 14812 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_161
timestamp 1667941163
transform 1 0 15916 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_169
timestamp 1667941163
transform 1 0 16652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_190
timestamp 1667941163
transform 1 0 18584 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_201
timestamp 1667941163
transform 1 0 19596 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_205
timestamp 1667941163
transform 1 0 19964 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_218
timestamp 1667941163
transform 1 0 21160 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_226
timestamp 1667941163
transform 1 0 21896 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_241
timestamp 1667941163
transform 1 0 23276 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1667941163
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_264
timestamp 1667941163
transform 1 0 25392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_284
timestamp 1667941163
transform 1 0 27232 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_305
timestamp 1667941163
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_328
timestamp 1667941163
transform 1 0 31280 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_335
timestamp 1667941163
transform 1 0 31924 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_342
timestamp 1667941163
transform 1 0 32568 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_354
timestamp 1667941163
transform 1 0 33672 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1667941163
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_385
timestamp 1667941163
transform 1 0 36524 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_8
timestamp 1667941163
transform 1 0 1840 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_19
timestamp 1667941163
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_31
timestamp 1667941163
transform 1 0 3956 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_42
timestamp 1667941163
transform 1 0 4968 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_63
timestamp 1667941163
transform 1 0 6900 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_67
timestamp 1667941163
transform 1 0 7268 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_74
timestamp 1667941163
transform 1 0 7912 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_88
timestamp 1667941163
transform 1 0 9200 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_92
timestamp 1667941163
transform 1 0 9568 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_96
timestamp 1667941163
transform 1 0 9936 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_103
timestamp 1667941163
transform 1 0 10580 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_146
timestamp 1667941163
transform 1 0 14536 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_153
timestamp 1667941163
transform 1 0 15180 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1667941163
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_191
timestamp 1667941163
transform 1 0 18676 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_202
timestamp 1667941163
transform 1 0 19688 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_209
timestamp 1667941163
transform 1 0 20332 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_216
timestamp 1667941163
transform 1 0 20976 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_230
timestamp 1667941163
transform 1 0 22264 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_244
timestamp 1667941163
transform 1 0 23552 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_248
timestamp 1667941163
transform 1 0 23920 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_270
timestamp 1667941163
transform 1 0 25944 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 1667941163
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_290
timestamp 1667941163
transform 1 0 27784 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_312
timestamp 1667941163
transform 1 0 29808 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_343
timestamp 1667941163
transform 1 0 32660 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_351
timestamp 1667941163
transform 1 0 33396 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_363
timestamp 1667941163
transform 1 0 34500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_371
timestamp 1667941163
transform 1 0 35236 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_377
timestamp 1667941163
transform 1 0 35788 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_50
timestamp 1667941163
transform 1 0 5704 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_71
timestamp 1667941163
transform 1 0 7636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_89
timestamp 1667941163
transform 1 0 9292 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_93
timestamp 1667941163
transform 1 0 9660 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_100
timestamp 1667941163
transform 1 0 10304 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1667941163
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_146
timestamp 1667941163
transform 1 0 14536 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1667941163
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_174
timestamp 1667941163
transform 1 0 17112 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_182
timestamp 1667941163
transform 1 0 17848 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_190
timestamp 1667941163
transform 1 0 18584 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_202
timestamp 1667941163
transform 1 0 19688 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_217
timestamp 1667941163
transform 1 0 21068 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1667941163
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_244
timestamp 1667941163
transform 1 0 23552 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_270
timestamp 1667941163
transform 1 0 25944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1667941163
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1667941163
transform 1 0 27416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_294
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_330
timestamp 1667941163
transform 1 0 31464 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_349
timestamp 1667941163
transform 1 0 33212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_399
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0384_
timestamp 1667941163
transform 1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0385_
timestamp 1667941163
transform 1 0 5796 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0386_
timestamp 1667941163
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0387_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0388_
timestamp 1667941163
transform 1 0 21068 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0389_
timestamp 1667941163
transform 1 0 19780 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0390_
timestamp 1667941163
transform 1 0 5888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0391_
timestamp 1667941163
transform 1 0 18952 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0392_
timestamp 1667941163
transform 1 0 18676 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0393_
timestamp 1667941163
transform 1 0 8832 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0394_
timestamp 1667941163
transform 1 0 20976 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0395_
timestamp 1667941163
transform 1 0 20884 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0396_
timestamp 1667941163
transform 1 0 19412 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0397_
timestamp 1667941163
transform 1 0 30360 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0398_
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0399_
timestamp 1667941163
transform 1 0 23276 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0400_
timestamp 1667941163
transform 1 0 23368 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0401_
timestamp 1667941163
transform 1 0 19044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0402_
timestamp 1667941163
transform 1 0 3680 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0403_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9016 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0404_
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0405_
timestamp 1667941163
transform 1 0 6532 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0406_
timestamp 1667941163
transform 1 0 11684 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0407_
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0408_
timestamp 1667941163
transform 1 0 7268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0409_
timestamp 1667941163
transform 1 0 19504 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0410_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0411_
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0412_
timestamp 1667941163
transform 1 0 10672 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0413_
timestamp 1667941163
transform 1 0 2300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0414_
timestamp 1667941163
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0415_
timestamp 1667941163
transform 1 0 5152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0416_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 17756 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0418_
timestamp 1667941163
transform 1 0 21620 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0419_
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0420_
timestamp 1667941163
transform 1 0 12696 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0421_
timestamp 1667941163
transform 1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 4600 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 21804 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0424_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0425_
timestamp 1667941163
transform 1 0 23184 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0426_
timestamp 1667941163
transform 1 0 11592 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0427_
timestamp 1667941163
transform 1 0 19044 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 6716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0430_
timestamp 1667941163
transform 1 0 22264 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0431_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0432_
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0433_
timestamp 1667941163
transform 1 0 20608 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 28336 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 28152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0436_
timestamp 1667941163
transform 1 0 16652 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0437_
timestamp 1667941163
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0438_
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0439_
timestamp 1667941163
transform 1 0 9108 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 13248 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 27324 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0442_
timestamp 1667941163
transform 1 0 27140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0443_
timestamp 1667941163
transform 1 0 19872 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0444_
timestamp 1667941163
transform 1 0 18308 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0445_
timestamp 1667941163
transform 1 0 24564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 23736 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform 1 0 23644 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0448_
timestamp 1667941163
transform 1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0449_
timestamp 1667941163
transform 1 0 21252 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1667941163
transform 1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1667941163
transform 1 0 19596 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1667941163
transform 1 0 28888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1667941163
transform 1 0 22908 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1667941163
transform 1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1667941163
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0456_
timestamp 1667941163
transform 1 0 23092 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1667941163
transform 1 0 28980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0458_
timestamp 1667941163
transform 1 0 27968 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0459_
timestamp 1667941163
transform 1 0 23920 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 27140 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0462_
timestamp 1667941163
transform 1 0 27784 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0463_
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0464_
timestamp 1667941163
transform 1 0 19688 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0465_
timestamp 1667941163
transform 1 0 27968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 22632 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0468_
timestamp 1667941163
transform 1 0 23736 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0469_
timestamp 1667941163
transform 1 0 25576 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0470_
timestamp 1667941163
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0471_
timestamp 1667941163
transform 1 0 19044 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 27232 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0474_
timestamp 1667941163
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0475_
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0476_
timestamp 1667941163
transform 1 0 25208 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1667941163
transform 1 0 24932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 14536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform 1 0 18032 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1667941163
transform 1 0 26128 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1667941163
transform 1 0 25760 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 27784 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 25944 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform 1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform 1 0 28428 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 30820 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 17112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform 1 0 19136 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform 1 0 24288 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 18400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 19688 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 23368 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 20608 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 8004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 2760 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 13248 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 19688 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30176 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 31648 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0508_
timestamp 1667941163
transform 1 0 11684 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0509_
timestamp 1667941163
transform 1 0 10304 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 8372 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0511_
timestamp 1667941163
transform 1 0 11500 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0512_
timestamp 1667941163
transform 1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 5704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 8096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0515_
timestamp 1667941163
transform 1 0 5060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform 1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1667941163
transform 1 0 3312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 3956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 5336 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0520_
timestamp 1667941163
transform 1 0 4416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0521_
timestamp 1667941163
transform 1 0 3772 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 19780 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0524_
timestamp 1667941163
transform 1 0 24380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0526_
timestamp 1667941163
transform 1 0 15548 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 22448 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0529_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0530_
timestamp 1667941163
transform 1 0 25208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 22448 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0533_
timestamp 1667941163
transform 1 0 23092 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 24656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0535_
timestamp 1667941163
transform 1 0 23092 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 21068 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0538_
timestamp 1667941163
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0539_
timestamp 1667941163
transform 1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 26496 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 18952 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0542_
timestamp 1667941163
transform 1 0 15364 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0544_
timestamp 1667941163
transform 1 0 28152 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 24932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1667941163
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 13524 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0550_
timestamp 1667941163
transform 1 0 25576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1667941163
transform 1 0 26312 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 4692 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 8372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform 1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0556_
timestamp 1667941163
transform 1 0 4968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1667941163
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 3956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 9844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1667941163
transform 1 0 24748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 23460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1667941163
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 15640 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform 1 0 22448 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0568_
timestamp 1667941163
transform 1 0 6808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0569_
timestamp 1667941163
transform 1 0 7636 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 29072 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 27784 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform 1 0 26404 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0574_
timestamp 1667941163
transform 1 0 7544 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0575_
timestamp 1667941163
transform 1 0 6624 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 28612 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1667941163
transform 1 0 28428 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 28980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1667941163
transform 1 0 24932 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 27140 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 28704 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 27784 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 26128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 24288 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 27140 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 19412 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 27784 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 18676 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 29716 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 27140 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 21804 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 23828 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 20516 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 25760 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 26772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 27048 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 10304 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 15088 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0611_
timestamp 1667941163
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0613_
timestamp 1667941163
transform 1 0 26128 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 2392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 35972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 28980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1667941163
transform 1 0 3956 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0618_
timestamp 1667941163
transform 1 0 37812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 33120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 30360 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 29716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 29072 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 4968 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1667941163
transform 1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 28244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 31464 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 14536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 2668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 7268 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 26312 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 6992 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 27140 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 23828 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 1840 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 27140 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 29716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 32292 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 14720 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 12880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 30544 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1667941163
transform 1 0 28520 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 11776 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 14444 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 25760 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1667941163
transform 1 0 19412 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 29348 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 13248 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 19688 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 28888 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 20148 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 29716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 29072 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1667941163
transform 1 0 5796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 32292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 25484 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 33764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1667941163
transform 1 0 23276 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 26128 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 30360 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 14536 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 30360 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 28336 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 19780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 11408 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 31832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 27876 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 14996 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 18952 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 29992 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 22632 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 17480 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 28428 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 28520 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 20056 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 1840 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 20700 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 4692 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 3956 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 9108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 20976 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 30360 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 27968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 7636 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 37260 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 14904 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 11684 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 26404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 29900 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 23736 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 2208 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0713_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24472 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _0714_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19964 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _0715_
timestamp 1667941163
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 10212 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 3036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 3220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 2576 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 3496 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 3220 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 19688 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 18308 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 18308 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0726_
timestamp 1667941163
transform 1 0 20608 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 25208 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 25576 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 23736 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 24564 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 22724 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 20792 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0737_
timestamp 1667941163
transform 1 0 19044 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 20332 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 20792 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 20700 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 22080 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 14260 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 19688 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 22356 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 23092 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 14168 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 22080 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0748_
timestamp 1667941163
transform 1 0 12880 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 3680 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 12328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 10304 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 13616 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 9292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0759_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11868 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 11684 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 14720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 6532 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 2208 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 8096 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 4416 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 5244 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0770_
timestamp 1667941163
transform 1 0 22724 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 23000 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 24932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 25208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 23092 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 22172 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 24748 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 20240 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 20424 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 20884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0781_
timestamp 1667941163
transform 1 0 21988 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 22632 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 23552 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 21620 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 25208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 25760 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 23368 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 23644 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 23184 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 21988 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 20976 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0792_
timestamp 1667941163
transform 1 0 17940 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 12236 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 19964 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 19964 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 20976 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 8740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0803_
timestamp 1667941163
transform 1 0 12880 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 8096 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 6808 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0814_
timestamp 1667941163
transform 1 0 11868 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 6532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 9660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 2576 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 4600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 4324 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 7268 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 18584 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 19044 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0825_
timestamp 1667941163
transform 1 0 21528 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 21528 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 3312 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 2576 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 2576 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 3404 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 3956 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 13524 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 12880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 20056 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 5244 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 1840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 2024 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 2300 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 5612 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 9476 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 4416 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0844_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6808 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0845_
timestamp 1667941163
transform 1 0 6348 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0846_
timestamp 1667941163
transform 1 0 2024 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0847_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2392 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0848_
timestamp 1667941163
transform 1 0 2392 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0849_
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0850_
timestamp 1667941163
transform 1 0 12788 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0851_
timestamp 1667941163
transform 1 0 16468 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0852_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0853_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0854_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0855_
timestamp 1667941163
transform 1 0 15916 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0856_
timestamp 1667941163
transform 1 0 16928 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0857_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0858_
timestamp 1667941163
transform 1 0 16836 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0859_
timestamp 1667941163
transform 1 0 16836 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0860_
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0861_
timestamp 1667941163
transform 1 0 11960 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0862_
timestamp 1667941163
transform 1 0 14260 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0863_
timestamp 1667941163
transform 1 0 16836 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0864_
timestamp 1667941163
transform 1 0 14260 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0865_
timestamp 1667941163
transform 1 0 16744 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0866_
timestamp 1667941163
transform 1 0 12696 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0867_
timestamp 1667941163
transform 1 0 14628 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0868_
timestamp 1667941163
transform 1 0 13800 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0869_
timestamp 1667941163
transform 1 0 16376 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0870_
timestamp 1667941163
transform 1 0 10948 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0871_
timestamp 1667941163
transform 1 0 16744 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0872_
timestamp 1667941163
transform 1 0 6072 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0873_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0874_
timestamp 1667941163
transform 1 0 1656 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0875_
timestamp 1667941163
transform 1 0 1748 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0876_
timestamp 1667941163
transform 1 0 6256 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1667941163
transform 1 0 3956 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0878_
timestamp 1667941163
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0879_
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0880_
timestamp 1667941163
transform 1 0 10580 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0881_
timestamp 1667941163
transform 1 0 13524 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0882_
timestamp 1667941163
transform 1 0 9752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0883_
timestamp 1667941163
transform 1 0 7268 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0884_
timestamp 1667941163
transform 1 0 10948 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0885_
timestamp 1667941163
transform 1 0 14720 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0886_
timestamp 1667941163
transform 1 0 4232 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0887_
timestamp 1667941163
transform 1 0 8188 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0888_
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0889_
timestamp 1667941163
transform 1 0 12052 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0890_
timestamp 1667941163
transform 1 0 11960 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1667941163
transform 1 0 6808 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 4232 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0893_
timestamp 1667941163
transform 1 0 3956 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0894_
timestamp 1667941163
transform 1 0 5060 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0895_
timestamp 1667941163
transform 1 0 3956 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0896_
timestamp 1667941163
transform 1 0 9016 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0897_
timestamp 1667941163
transform 1 0 8188 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0898_
timestamp 1667941163
transform 1 0 16928 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0899_
timestamp 1667941163
transform 1 0 16560 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0900_
timestamp 1667941163
transform 1 0 15824 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0901_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1667941163
transform 1 0 11684 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0903_
timestamp 1667941163
transform 1 0 16836 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0904_
timestamp 1667941163
transform 1 0 13248 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0905_
timestamp 1667941163
transform 1 0 12236 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0906_
timestamp 1667941163
transform 1 0 12236 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0907_
timestamp 1667941163
transform 1 0 3956 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 8096 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0909_
timestamp 1667941163
transform 1 0 8924 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0910_
timestamp 1667941163
transform 1 0 16836 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0911_
timestamp 1667941163
transform 1 0 16836 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0912_
timestamp 1667941163
transform 1 0 13248 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0913_
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 11868 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0915_
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0916_
timestamp 1667941163
transform 1 0 14720 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0917_
timestamp 1667941163
transform 1 0 16836 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform 1 0 16836 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1667941163
transform 1 0 15916 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0920_
timestamp 1667941163
transform 1 0 13156 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0921_
timestamp 1667941163
transform 1 0 11592 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 4600 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0923_
timestamp 1667941163
transform 1 0 9384 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 9108 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0926_
timestamp 1667941163
transform 1 0 14076 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0927_
timestamp 1667941163
transform 1 0 16560 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 13340 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0929_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1667941163
transform 1 0 11040 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 6808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 6900 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0934_
timestamp 1667941163
transform 1 0 10396 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0935_
timestamp 1667941163
transform 1 0 7728 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0936_
timestamp 1667941163
transform 1 0 9108 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0937_
timestamp 1667941163
transform 1 0 3956 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform 1 0 3956 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 1656 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1667941163
transform 1 0 4600 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0942_
timestamp 1667941163
transform 1 0 15088 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1667941163
transform 1 0 16836 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0944_
timestamp 1667941163
transform 1 0 11776 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0945_
timestamp 1667941163
transform 1 0 11224 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0946_
timestamp 1667941163
transform 1 0 4140 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1667941163
transform 1 0 1564 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0951_
timestamp 1667941163
transform 1 0 6716 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0952_
timestamp 1667941163
transform 1 0 9660 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0953_
timestamp 1667941163
transform 1 0 12420 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0954_
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0955_
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1667941163
transform 1 0 5060 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1667941163
transform 1 0 3404 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0958_
timestamp 1667941163
transform 1 0 6532 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0959_
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0960_
timestamp 1667941163
transform 1 0 10212 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0961_
timestamp 1667941163
transform 1 0 6256 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1667941163
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1667941163
transform 1 0 2944 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1667941163
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0991_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19872 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1667941163
transform 1 0 37352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 21988 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 37812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1667941163
transform 1 0 29716 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1667941163
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 24840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 20792 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1667941163
transform 1 0 22632 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1000_
timestamp 1667941163
transform 1 0 27600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1001_
timestamp 1667941163
transform 1 0 31372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 31280 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 26312 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 12052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 1564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1007_
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1008_
timestamp 1667941163
transform 1 0 13156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 2300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1011_
timestamp 1667941163
transform 1 0 26312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 14260 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 32384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 9016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 37628 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1016_
timestamp 1667941163
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 27140 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 37812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform 1 0 27140 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 27140 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 28796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 28980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 6716 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 34684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1028_
timestamp 1667941163
transform 1 0 32292 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 33304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1667941163
transform 1 0 32384 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform 1 0 3956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 5428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 4508 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1667941163
transform 1 0 35328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 37812 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1667941163
transform 1 0 37812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1667941163
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1044_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8280 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1045__142 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1045_
timestamp 1667941163
transform 1 0 15088 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1046_
timestamp 1667941163
transform 1 0 11684 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1047_
timestamp 1667941163
transform 1 0 2208 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1048_
timestamp 1667941163
transform 1 0 11684 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1049_
timestamp 1667941163
transform 1 0 15456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1050_
timestamp 1667941163
transform 1 0 9476 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1052_
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1053_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25484 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1054_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1055_
timestamp 1667941163
transform 1 0 29716 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1055__143
timestamp 1667941163
transform 1 0 29900 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1056_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1057_
timestamp 1667941163
transform 1 0 21896 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1058_
timestamp 1667941163
transform 1 0 24840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1059_
timestamp 1667941163
transform 1 0 22632 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1060_
timestamp 1667941163
transform 1 0 22080 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1061_
timestamp 1667941163
transform 1 0 26496 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1062__144
timestamp 1667941163
transform 1 0 31464 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1062_
timestamp 1667941163
transform 1 0 28980 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1063_
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1064_
timestamp 1667941163
transform 1 0 26036 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1065_
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1066_
timestamp 1667941163
transform 1 0 20700 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1067_
timestamp 1667941163
transform 1 0 24840 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1068__145
timestamp 1667941163
transform 1 0 31188 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1068_
timestamp 1667941163
transform 1 0 31004 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1069_
timestamp 1667941163
transform 1 0 26680 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1070_
timestamp 1667941163
transform 1 0 27600 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1071_
timestamp 1667941163
transform 1 0 27876 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1072_
timestamp 1667941163
transform 1 0 29716 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1073__146
timestamp 1667941163
transform 1 0 28428 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1073_
timestamp 1667941163
transform 1 0 27600 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1074_
timestamp 1667941163
transform 1 0 28244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1075_
timestamp 1667941163
transform 1 0 27140 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 27508 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1077__147
timestamp 1667941163
transform 1 0 5612 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1077_
timestamp 1667941163
transform 1 0 5428 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1078_
timestamp 1667941163
transform 1 0 23184 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1079_
timestamp 1667941163
transform 1 0 24564 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1080_
timestamp 1667941163
transform 1 0 22540 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1081_
timestamp 1667941163
transform 1 0 9108 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1081__148
timestamp 1667941163
transform 1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1082_
timestamp 1667941163
transform 1 0 20608 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1083_
timestamp 1667941163
transform 1 0 6624 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1084_
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1085_
timestamp 1667941163
transform 1 0 2392 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1085__149
timestamp 1667941163
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1086_
timestamp 1667941163
transform 1 0 25576 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1087_
timestamp 1667941163
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1088_
timestamp 1667941163
transform 1 0 9936 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1089__150
timestamp 1667941163
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1089_
timestamp 1667941163
transform 1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1090_
timestamp 1667941163
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1091_
timestamp 1667941163
transform 1 0 4048 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1092_
timestamp 1667941163
transform 1 0 8004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1093_
timestamp 1667941163
transform 1 0 27140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1093__151
timestamp 1667941163
transform 1 0 26956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1094_
timestamp 1667941163
transform 1 0 13248 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1095_
timestamp 1667941163
transform 1 0 25024 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform 1 0 12052 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1097_
timestamp 1667941163
transform 1 0 28520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1097__152
timestamp 1667941163
transform 1 0 28704 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1098_
timestamp 1667941163
transform 1 0 17296 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1099_
timestamp 1667941163
transform 1 0 26220 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1100_
timestamp 1667941163
transform 1 0 18952 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1101_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1102_
timestamp 1667941163
transform 1 0 20332 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1102__153
timestamp 1667941163
transform 1 0 20424 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1103_
timestamp 1667941163
transform 1 0 23552 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1104_
timestamp 1667941163
transform 1 0 23184 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1105_
timestamp 1667941163
transform 1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1106_
timestamp 1667941163
transform 1 0 23092 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1107_
timestamp 1667941163
transform 1 0 14904 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1108__154
timestamp 1667941163
transform 1 0 24288 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1108_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1109_
timestamp 1667941163
transform 1 0 23644 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1110_
timestamp 1667941163
transform 1 0 14444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1111_
timestamp 1667941163
transform 1 0 23184 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1112_
timestamp 1667941163
transform 1 0 20056 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1113_
timestamp 1667941163
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1114__155
timestamp 1667941163
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1114_
timestamp 1667941163
transform 1 0 3956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 6624 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1116_
timestamp 1667941163
transform 1 0 6624 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1117_
timestamp 1667941163
transform 1 0 6532 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1118_
timestamp 1667941163
transform 1 0 7728 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1119_
timestamp 1667941163
transform 1 0 9200 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1120__156
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1120_
timestamp 1667941163
transform 1 0 10396 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1121_
timestamp 1667941163
transform 1 0 24380 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1122_
timestamp 1667941163
transform 1 0 27784 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1123_
timestamp 1667941163
transform 1 0 8464 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1124_
timestamp 1667941163
transform 1 0 21988 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1125_
timestamp 1667941163
transform 1 0 7452 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1126_
timestamp 1667941163
transform 1 0 26220 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1127_
timestamp 1667941163
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1128__157
timestamp 1667941163
transform 1 0 25760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1128_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1129_
timestamp 1667941163
transform 1 0 2392 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1130_
timestamp 1667941163
transform 1 0 10948 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1131_
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 18216 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1133_
timestamp 1667941163
transform 1 0 19688 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1134_
timestamp 1667941163
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1135_
timestamp 1667941163
transform 1 0 2300 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1136_
timestamp 1667941163
transform 1 0 25392 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1137_
timestamp 1667941163
transform 1 0 20332 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1138_
timestamp 1667941163
transform 1 0 20240 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1139_
timestamp 1667941163
transform 1 0 19780 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1140__158
timestamp 1667941163
transform 1 0 26404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1140_
timestamp 1667941163
transform 1 0 25760 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1141_
timestamp 1667941163
transform 1 0 17204 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1142_
timestamp 1667941163
transform 1 0 30084 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1143_
timestamp 1667941163
transform 1 0 24196 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 25760 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1145_
timestamp 1667941163
transform 1 0 20056 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1146_
timestamp 1667941163
transform 1 0 27140 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1147_
timestamp 1667941163
transform 1 0 26128 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1148_
timestamp 1667941163
transform 1 0 25116 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1149_
timestamp 1667941163
transform 1 0 25576 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1150_
timestamp 1667941163
transform 1 0 25760 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1151_
timestamp 1667941163
transform 1 0 12512 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1152__159
timestamp 1667941163
transform 1 0 27600 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1152_
timestamp 1667941163
transform 1 0 27508 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1153_
timestamp 1667941163
transform 1 0 15824 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1154_
timestamp 1667941163
transform 1 0 11684 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1155_
timestamp 1667941163
transform 1 0 20516 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 19596 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1157_
timestamp 1667941163
transform 1 0 23552 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1158_
timestamp 1667941163
transform 1 0 27508 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1159_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1160_
timestamp 1667941163
transform 1 0 25852 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1161_
timestamp 1667941163
transform 1 0 22356 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1162_
timestamp 1667941163
transform 1 0 24656 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1163_
timestamp 1667941163
transform 1 0 24564 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1164__160
timestamp 1667941163
transform 1 0 29716 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1164_
timestamp 1667941163
transform 1 0 28796 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 27140 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1167_
timestamp 1667941163
transform 1 0 23552 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 28152 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1169_
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1170_
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1171_
timestamp 1667941163
transform 1 0 27784 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1172_
timestamp 1667941163
transform 1 0 30360 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _1173_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22264 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1174_
timestamp 1667941163
transform 1 0 10672 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1175__161
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1175_
timestamp 1667941163
transform 1 0 26128 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1176_
timestamp 1667941163
transform 1 0 24288 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1177_
timestamp 1667941163
transform 1 0 25484 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1178_
timestamp 1667941163
transform 1 0 23828 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1179_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1180_
timestamp 1667941163
transform 1 0 24564 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1181_
timestamp 1667941163
transform 1 0 22908 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1182_
timestamp 1667941163
transform 1 0 19504 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1183_
timestamp 1667941163
transform 1 0 27968 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1184_
timestamp 1667941163
transform 1 0 23092 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1185_
timestamp 1667941163
transform 1 0 9200 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1186_
timestamp 1667941163
transform 1 0 10028 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1187_
timestamp 1667941163
transform 1 0 5244 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1187__162
timestamp 1667941163
transform 1 0 5336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1188_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1189_
timestamp 1667941163
transform 1 0 25484 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1190_
timestamp 1667941163
transform 1 0 26036 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1191_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1192_
timestamp 1667941163
transform 1 0 29440 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1193_
timestamp 1667941163
transform 1 0 28796 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1194_
timestamp 1667941163
transform 1 0 9568 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1195_
timestamp 1667941163
transform 1 0 12144 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1196_
timestamp 1667941163
transform 1 0 29992 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1197_
timestamp 1667941163
transform 1 0 17756 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1198_
timestamp 1667941163
transform 1 0 16744 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1199_
timestamp 1667941163
transform 1 0 23184 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1199__163
timestamp 1667941163
transform 1 0 23368 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1200_
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1201_
timestamp 1667941163
transform 1 0 23552 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1202_
timestamp 1667941163
transform 1 0 9108 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1203_
timestamp 1667941163
transform 1 0 22724 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1204_
timestamp 1667941163
transform 1 0 20332 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1205_
timestamp 1667941163
transform 1 0 2300 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1206_
timestamp 1667941163
transform 1 0 15180 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1207_
timestamp 1667941163
transform 1 0 7452 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1208_
timestamp 1667941163
transform 1 0 4232 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1209_
timestamp 1667941163
transform 1 0 6532 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1210_
timestamp 1667941163
transform 1 0 2300 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1211_
timestamp 1667941163
transform 1 0 2668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1211__164
timestamp 1667941163
transform 1 0 3128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1212_
timestamp 1667941163
transform 1 0 21804 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1213_
timestamp 1667941163
transform 1 0 22356 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1214_
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1215_
timestamp 1667941163
transform 1 0 11316 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1216_
timestamp 1667941163
transform 1 0 23460 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1217_
timestamp 1667941163
transform 1 0 21804 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1218_
timestamp 1667941163
transform 1 0 6624 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1219_
timestamp 1667941163
transform 1 0 17664 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1220_
timestamp 1667941163
transform 1 0 21528 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1221_
timestamp 1667941163
transform 1 0 27876 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1222_
timestamp 1667941163
transform 1 0 1840 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1223_
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1223__165
timestamp 1667941163
transform 1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1224_
timestamp 1667941163
transform 1 0 10028 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1225_
timestamp 1667941163
transform 1 0 10396 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1226_
timestamp 1667941163
transform 1 0 6348 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1227_
timestamp 1667941163
transform 1 0 24564 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1228_
timestamp 1667941163
transform 1 0 22080 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1229_
timestamp 1667941163
transform 1 0 30176 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1230_
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1231_
timestamp 1667941163
transform 1 0 20976 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1232_
timestamp 1667941163
transform 1 0 30268 0 1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1233_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1234_
timestamp 1667941163
transform 1 0 4140 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1235_
timestamp 1667941163
transform 1 0 19596 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1235__166
timestamp 1667941163
transform 1 0 19688 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1236_
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1237_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1238_
timestamp 1667941163
transform 1 0 21988 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1239_
timestamp 1667941163
transform 1 0 22632 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1240_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1241_
timestamp 1667941163
transform 1 0 4508 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1242_
timestamp 1667941163
transform 1 0 7360 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1243_
timestamp 1667941163
transform 1 0 20608 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1244_
timestamp 1667941163
transform 1 0 4048 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10212 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk
timestamp 1667941163
transform 1 0 5888 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 7728 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 4140 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 9108 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 11868 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 14168 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 11316 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 6164 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 10212 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 6624 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 10304 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 15364 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 17480 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 14260 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12880 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1667941163
transform 1 0 1564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1667941163
transform 1 0 37444 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 26956 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1667941163
transform 1 0 37444 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform 1 0 1564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 29716 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1667941163
transform 1 0 37444 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 4692 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 16100 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 38088 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 1564 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 38088 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 26312 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 14904 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 10304 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 38088 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 38088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 36708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1667941163
transform 1 0 37444 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 38088 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 1564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 2668 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 36616 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 1564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 37352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 2208 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1667941163
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1667941163
transform 1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1667941163
transform 1 0 35512 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1667941163
transform 1 0 37444 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1667941163
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1667941163
transform 1 0 38088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1667941163
transform 1 0 32292 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1667941163
transform 1 0 31004 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 5796 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1667941163
transform 1 0 2576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 38088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 37996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 33028 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 33764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 1564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 10856 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform 1 0 27784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 17480 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 30452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  sb_1__0__141
timestamp 1667941163
transform 1 0 38088 0 1 20672
box -38 -48 314 592
<< labels >>
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 2 nsew signal input
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 3 nsew signal input
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 4 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 5 nsew signal input
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 6 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_left_in[14]
port 7 nsew signal input
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 8 nsew signal input
flabel metal3 s 39200 8168 39800 8288 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 9 nsew signal input
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 10 nsew signal input
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 11 nsew signal input
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 12 nsew signal input
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chanx_left_in[2]
port 13 nsew signal input
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 14 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 15 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 16 nsew signal input
flabel metal2 s 28354 200 28410 800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 17 nsew signal input
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chanx_left_in[7]
port 18 nsew signal input
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 19 nsew signal input
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chanx_left_in[9]
port 20 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 21 nsew signal tristate
flabel metal2 s 20626 200 20682 800 0 FreeSans 224 90 0 0 chanx_left_out[10]
port 22 nsew signal tristate
flabel metal3 s 39200 27888 39800 28008 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 23 nsew signal tristate
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 24 nsew signal tristate
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_left_out[13]
port 25 nsew signal tristate
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 26 nsew signal tristate
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 27 nsew signal tristate
flabel metal2 s 17406 200 17462 800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 28 nsew signal tristate
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 29 nsew signal tristate
flabel metal2 s 10966 200 11022 800 0 FreeSans 224 90 0 0 chanx_left_out[18]
port 30 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 31 nsew signal tristate
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 32 nsew signal tristate
flabel metal3 s 39200 12928 39800 13048 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 33 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 34 nsew signal tristate
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 35 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 36 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 37 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 38 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 39 nsew signal tristate
flabel metal3 s 39200 16328 39800 16448 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 40 nsew signal input
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 41 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 42 nsew signal input
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 43 nsew signal input
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 44 nsew signal input
flabel metal3 s 200 4088 800 4208 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 45 nsew signal input
flabel metal3 s 39200 17688 39800 17808 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 46 nsew signal input
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 47 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 48 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 49 nsew signal input
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 50 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chanx_right_in[2]
port 51 nsew signal input
flabel metal2 s 18694 39200 18750 39800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 52 nsew signal input
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 chanx_right_in[4]
port 53 nsew signal input
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 54 nsew signal input
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 55 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 56 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 57 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 58 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 59 nsew signal tristate
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 60 nsew signal tristate
flabel metal3 s 200 14968 800 15088 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 61 nsew signal tristate
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 62 nsew signal tristate
flabel metal2 s 10966 39200 11022 39800 0 FreeSans 224 90 0 0 chanx_right_out[13]
port 63 nsew signal tristate
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 64 nsew signal tristate
flabel metal3 s 200 21768 800 21888 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 65 nsew signal tristate
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 66 nsew signal tristate
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 67 nsew signal tristate
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chanx_right_out[18]
port 68 nsew signal tristate
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 69 nsew signal tristate
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 70 nsew signal tristate
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 71 nsew signal tristate
flabel metal3 s 39200 4768 39800 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 72 nsew signal tristate
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 73 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 74 nsew signal tristate
flabel metal2 s 17406 39200 17462 39800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 75 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 76 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 77 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_top_in[0]
port 78 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 79 nsew signal input
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chany_top_in[11]
port 80 nsew signal input
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chany_top_in[12]
port 81 nsew signal input
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_top_in[13]
port 82 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_top_in[14]
port 83 nsew signal input
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_top_in[15]
port 84 nsew signal input
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_top_in[16]
port 85 nsew signal input
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_top_in[17]
port 86 nsew signal input
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 87 nsew signal input
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_top_in[1]
port 88 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_top_in[2]
port 89 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chany_top_in[3]
port 90 nsew signal input
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_in[4]
port 91 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_top_in[5]
port 92 nsew signal input
flabel metal3 s 200 18368 800 18488 0 FreeSans 480 0 0 0 chany_top_in[6]
port 93 nsew signal input
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_top_in[7]
port 94 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_top_in[8]
port 95 nsew signal input
flabel metal2 s 14186 39200 14242 39800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 96 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_top_out[0]
port 97 nsew signal tristate
flabel metal2 s 3882 200 3938 800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 98 nsew signal tristate
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chany_top_out[11]
port 99 nsew signal tristate
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_top_out[12]
port 100 nsew signal tristate
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_top_out[13]
port 101 nsew signal tristate
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chany_top_out[14]
port 102 nsew signal tristate
flabel metal2 s 32862 200 32918 800 0 FreeSans 224 90 0 0 chany_top_out[15]
port 103 nsew signal tristate
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_top_out[16]
port 104 nsew signal tristate
flabel metal3 s 39200 9528 39800 9648 0 FreeSans 480 0 0 0 chany_top_out[17]
port 105 nsew signal tristate
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_top_out[18]
port 106 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_top_out[2]
port 108 nsew signal tristate
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 109 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_top_out[4]
port 110 nsew signal tristate
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_top_out[5]
port 111 nsew signal tristate
flabel metal3 s 200 2048 800 2168 0 FreeSans 480 0 0 0 chany_top_out[6]
port 112 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_top_out[7]
port 113 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[8]
port 114 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 115 nsew signal tristate
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 116 nsew signal input
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 117 nsew signal input
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 118 nsew signal input
flabel metal3 s 200 29928 800 30048 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 119 nsew signal input
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 120 nsew signal input
flabel metal2 s 1950 200 2006 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 121 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 122 nsew signal input
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 123 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 124 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 125 nsew signal input
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 pReset
port 126 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 prog_clk
port 127 nsew signal input
flabel metal3 s 200 11568 800 11688 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 128 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 129 nsew signal input
flabel metal2 s 14186 200 14242 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 130 nsew signal input
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 131 nsew signal input
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 132 nsew signal input
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 133 nsew signal input
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 134 nsew signal input
flabel metal2 s 28354 39200 28410 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 135 nsew signal input
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 136 nsew signal input
flabel metal2 s 6458 39200 6514 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 137 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 138 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 139 nsew signal input
flabel metal3 s 200 34688 800 34808 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 140 nsew signal input
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 141 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 143 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 3956 16490 3956 16490 0 _0000_
rlabel metal1 7820 18394 7820 18394 0 _0001_
rlabel metal2 2898 33694 2898 33694 0 _0002_
rlabel metal1 12643 31382 12643 31382 0 _0003_
rlabel metal1 8188 22134 8188 22134 0 _0004_
rlabel metal1 5474 22950 5474 22950 0 _0005_
rlabel metal1 6578 16524 6578 16524 0 _0006_
rlabel metal1 6026 23494 6026 23494 0 _0007_
rlabel metal2 6486 32929 6486 32929 0 _0008_
rlabel metal1 25162 34510 25162 34510 0 _0009_
rlabel metal1 22080 25772 22080 25772 0 _0010_
rlabel metal1 12420 28152 12420 28152 0 _0011_
rlabel metal2 20194 30430 20194 30430 0 _0012_
rlabel metal2 20194 27404 20194 27404 0 _0013_
rlabel metal1 17763 27438 17763 27438 0 _0014_
rlabel metal1 19320 29478 19320 29478 0 _0015_
rlabel metal1 18630 31246 18630 31246 0 _0016_
rlabel metal1 20838 29478 20838 29478 0 _0017_
rlabel metal1 21574 24616 21574 24616 0 _0018_
rlabel metal2 21390 23936 21390 23936 0 _0019_
rlabel metal1 21252 26282 21252 26282 0 _0020_
rlabel metal2 13018 26928 13018 26928 0 _0021_
rlabel metal1 10994 31416 10994 31416 0 _0022_
rlabel metal2 13110 32606 13110 32606 0 _0023_
rlabel metal2 19274 32793 19274 32793 0 _0024_
rlabel metal1 18499 32878 18499 32878 0 _0025_
rlabel metal1 18354 33320 18354 33320 0 _0026_
rlabel metal1 17112 26554 17112 26554 0 _0027_
rlabel metal2 13662 17986 13662 17986 0 _0028_
rlabel metal2 13754 23222 13754 23222 0 _0029_
rlabel metal1 19688 24310 19688 24310 0 _0030_
rlabel metal2 20470 26112 20470 26112 0 _0031_
rlabel metal2 20102 28254 20102 28254 0 _0032_
rlabel metal1 19826 33082 19826 33082 0 _0033_
rlabel metal1 21298 34918 21298 34918 0 _0034_
rlabel metal3 17434 32028 17434 32028 0 _0035_
rlabel metal1 3864 16422 3864 16422 0 _0036_
rlabel metal1 9292 16218 9292 16218 0 _0037_
rlabel metal2 10442 18360 10442 18360 0 _0038_
rlabel metal1 18223 17578 18223 17578 0 _0039_
rlabel metal1 16882 20230 16882 20230 0 _0040_
rlabel metal1 19504 18938 19504 18938 0 _0041_
rlabel metal1 14122 17306 14122 17306 0 _0042_
rlabel metal2 17802 18360 17802 18360 0 _0043_
rlabel metal1 11178 16218 11178 16218 0 _0044_
rlabel metal1 11546 14586 11546 14586 0 _0045_
rlabel metal2 8234 17476 8234 17476 0 _0046_
rlabel metal1 7084 16218 7084 16218 0 _0047_
rlabel metal1 7544 15674 7544 15674 0 _0048_
rlabel metal1 15594 22440 15594 22440 0 _0049_
rlabel metal1 9844 21114 9844 21114 0 _0050_
rlabel metal2 4738 17884 4738 17884 0 _0051_
rlabel metal1 4876 21454 4876 21454 0 _0052_
rlabel metal1 3227 19754 3227 19754 0 _0053_
rlabel metal1 4278 17238 4278 17238 0 _0054_
rlabel metal1 6585 20842 6585 20842 0 _0055_
rlabel metal1 17119 21930 17119 21930 0 _0056_
rlabel metal2 19182 26520 19182 26520 0 _0057_
rlabel metal2 22126 32096 22126 32096 0 _0058_
rlabel metal1 12650 28567 12650 28567 0 _0059_
rlabel metal1 4409 25942 4409 25942 0 _0060_
rlabel metal2 2714 35785 2714 35785 0 _0061_
rlabel metal1 2668 35462 2668 35462 0 _0062_
rlabel metal1 4179 34646 4179 34646 0 _0063_
rlabel metal1 4370 34170 4370 34170 0 _0064_
rlabel metal2 8142 35122 8142 35122 0 _0065_
rlabel metal1 11415 32810 11415 32810 0 _0066_
rlabel metal1 18630 35802 18630 35802 0 _0067_
rlabel metal1 6801 23766 6801 23766 0 _0068_
rlabel metal2 4646 24344 4646 24344 0 _0069_
rlabel metal2 3358 26282 3358 26282 0 _0070_
rlabel metal2 4738 28526 4738 28526 0 _0071_
rlabel metal1 4048 32198 4048 32198 0 _0072_
rlabel metal1 14674 32878 14674 32878 0 _0073_
rlabel metal1 10396 29002 10396 29002 0 _0074_
rlabel metal1 5796 27302 5796 27302 0 _0075_
rlabel metal1 8609 20910 8609 20910 0 _0076_
rlabel metal1 5152 17306 5152 17306 0 _0077_
rlabel metal2 3358 17272 3358 17272 0 _0078_
rlabel metal1 2346 16422 2346 16422 0 _0079_
rlabel metal1 3680 25670 3680 25670 0 _0080_
rlabel metal1 3135 27370 3135 27370 0 _0081_
rlabel metal2 13662 28254 13662 28254 0 _0082_
rlabel metal1 17947 24174 17947 24174 0 _0083_
rlabel metal2 18446 24174 18446 24174 0 _0084_
rlabel metal2 18446 17816 18446 17816 0 _0085_
rlabel metal1 19235 21590 19235 21590 0 _0086_
rlabel metal1 18315 20910 18315 20910 0 _0087_
rlabel metal1 18354 33449 18354 33449 0 _0088_
rlabel metal2 21574 35122 21574 35122 0 _0089_
rlabel metal1 20194 34680 20194 34680 0 _0090_
rlabel metal1 18262 35095 18262 35095 0 _0091_
rlabel metal1 21206 36176 21206 36176 0 _0092_
rlabel metal1 14819 33898 14819 33898 0 _0093_
rlabel metal1 20010 30022 20010 30022 0 _0094_
rlabel metal1 19787 31382 19787 31382 0 _0095_
rlabel metal1 19918 32198 19918 32198 0 _0096_
rlabel metal1 18453 31790 18453 31790 0 _0097_
rlabel metal1 20792 35802 20792 35802 0 _0098_
rlabel metal1 16613 34986 16613 34986 0 _0099_
rlabel metal2 14398 33864 14398 33864 0 _0100_
rlabel metal1 18039 29614 18039 29614 0 _0101_
rlabel metal1 13669 34986 13669 34986 0 _0102_
rlabel metal2 18170 36380 18170 36380 0 _0103_
rlabel metal1 9345 25194 9345 25194 0 _0104_
rlabel metal2 13754 33864 13754 33864 0 _0105_
rlabel metal1 3128 12954 3128 12954 0 _0106_
rlabel metal1 1932 17510 1932 17510 0 _0107_
rlabel metal1 2116 12410 2116 12410 0 _0108_
rlabel metal1 4370 12954 4370 12954 0 _0109_
rlabel metal1 12604 15130 12604 15130 0 _0110_
rlabel metal2 2898 17000 2898 17000 0 _0111_
rlabel metal1 10902 20774 10902 20774 0 _0112_
rlabel metal2 13754 17306 13754 17306 0 _0113_
rlabel metal1 9982 15674 9982 15674 0 _0114_
rlabel metal1 7130 16014 7130 16014 0 _0115_
rlabel metal1 11776 18394 11776 18394 0 _0116_
rlabel metal1 14996 16558 14996 16558 0 _0117_
rlabel metal2 13202 15776 13202 15776 0 _0118_
rlabel metal1 2254 34612 2254 34612 0 _0119_
rlabel metal2 20930 29444 20930 29444 0 _0120_
rlabel metal1 21344 26350 21344 26350 0 _0121_
rlabel metal1 12558 16558 12558 16558 0 _0122_
rlabel metal1 13938 17136 13938 17136 0 _0123_
rlabel metal2 2622 15980 2622 15980 0 _0124_
rlabel metal1 21988 32402 21988 32402 0 _0125_
rlabel metal2 31878 35836 31878 35836 0 _0126_
rlabel metal1 11132 34714 11132 34714 0 _0127_
rlabel metal1 11316 35666 11316 35666 0 _0128_
rlabel metal1 5336 13294 5336 13294 0 _0129_
rlabel metal1 4186 11764 4186 11764 0 _0130_
rlabel metal1 4232 9554 4232 9554 0 _0131_
rlabel metal2 24426 14212 24426 14212 0 _0132_
rlabel metal1 15134 11118 15134 11118 0 _0133_
rlabel metal1 25438 9996 25438 9996 0 _0134_
rlabel metal1 23598 18394 23598 18394 0 _0135_
rlabel metal1 22816 10030 22816 10030 0 _0136_
rlabel metal2 21022 8058 21022 8058 0 _0137_
rlabel metal2 16330 16252 16330 16252 0 _0138_
rlabel metal1 29026 25228 29026 25228 0 _0139_
rlabel metal1 13984 10642 13984 10642 0 _0140_
rlabel metal2 26542 11322 26542 11322 0 _0141_
rlabel metal1 9154 14042 9154 14042 0 _0142_
rlabel metal1 4600 8942 4600 8942 0 _0143_
rlabel metal1 24242 20570 24242 20570 0 _0144_
rlabel metal1 4416 12206 4416 12206 0 _0145_
rlabel metal2 22126 24429 22126 24429 0 _0146_
rlabel metal2 7866 10948 7866 10948 0 _0147_
rlabel metal1 27278 33422 27278 33422 0 _0148_
rlabel metal1 7222 31994 7222 31994 0 _0149_
rlabel metal1 28842 27574 28842 27574 0 _0150_
rlabel metal1 26082 31314 26082 31314 0 _0151_
rlabel metal1 19826 18394 19826 18394 0 _0152_
rlabel metal1 1794 23732 1794 23732 0 _0153_
rlabel metal1 2622 16593 2622 16593 0 _0154_
rlabel metal1 20838 21522 20838 21522 0 _0155_
rlabel metal1 18814 32878 18814 32878 0 _0156_
rlabel metal1 7820 10710 7820 10710 0 _0157_
rlabel metal1 15272 12070 15272 12070 0 _0158_
rlabel metal1 11178 9622 11178 9622 0 _0159_
rlabel metal1 2300 9962 2300 9962 0 _0160_
rlabel metal2 11914 11152 11914 11152 0 _0161_
rlabel metal2 15686 11152 15686 11152 0 _0162_
rlabel metal2 9706 10846 9706 10846 0 _0163_
rlabel metal2 9246 9758 9246 9758 0 _0164_
rlabel metal2 17986 10438 17986 10438 0 _0165_
rlabel metal1 26450 24786 26450 24786 0 _0166_
rlabel metal1 24840 24106 24840 24106 0 _0167_
rlabel metal1 28750 25942 28750 25942 0 _0168_
rlabel metal1 22172 18258 22172 18258 0 _0169_
rlabel metal2 21390 17884 21390 17884 0 _0170_
rlabel metal1 25070 23732 25070 23732 0 _0171_
rlabel metal1 22402 24310 22402 24310 0 _0172_
rlabel metal1 22310 18700 22310 18700 0 _0173_
rlabel metal2 26726 34136 26726 34136 0 _0174_
rlabel metal2 29854 35224 29854 35224 0 _0175_
rlabel metal2 20562 36210 20562 36210 0 _0176_
rlabel metal1 26266 32776 26266 32776 0 _0177_
rlabel metal2 27922 35224 27922 35224 0 _0178_
rlabel metal1 20746 34646 20746 34646 0 _0179_
rlabel metal1 24748 33558 24748 33558 0 _0180_
rlabel metal1 30774 23018 30774 23018 0 _0181_
rlabel metal1 27094 34510 27094 34510 0 _0182_
rlabel metal1 27830 32776 27830 32776 0 _0183_
rlabel metal1 27692 33354 27692 33354 0 _0184_
rlabel metal1 29394 30294 29394 30294 0 _0185_
rlabel metal2 27830 30668 27830 30668 0 _0186_
rlabel metal2 29026 28628 29026 28628 0 _0187_
rlabel metal1 27048 29138 27048 29138 0 _0188_
rlabel metal1 28244 28594 28244 28594 0 _0189_
rlabel metal1 5658 32776 5658 32776 0 _0190_
rlabel metal1 25484 33626 25484 33626 0 _0191_
rlabel metal2 27462 34272 27462 34272 0 _0192_
rlabel metal2 23460 31892 23460 31892 0 _0193_
rlabel metal1 8510 10778 8510 10778 0 _0194_
rlabel metal1 21482 24072 21482 24072 0 _0195_
rlabel metal1 6486 12274 6486 12274 0 _0196_
rlabel metal1 16514 13192 16514 13192 0 _0197_
rlabel metal1 3220 14382 3220 14382 0 _0198_
rlabel metal2 25806 20638 25806 20638 0 _0199_
rlabel metal1 3542 13498 3542 13498 0 _0200_
rlabel metal2 10166 15912 10166 15912 0 _0201_
rlabel metal2 3082 8636 3082 8636 0 _0202_
rlabel metal1 9246 10234 9246 10234 0 _0203_
rlabel metal1 4554 10642 4554 10642 0 _0204_
rlabel metal1 8050 11730 8050 11730 0 _0205_
rlabel metal1 26864 11322 26864 11322 0 _0206_
rlabel metal1 13524 10778 13524 10778 0 _0207_
rlabel metal1 25162 11866 25162 11866 0 _0208_
rlabel metal1 11822 11798 11822 11798 0 _0209_
rlabel metal1 28796 25466 28796 25466 0 _0210_
rlabel metal1 16836 16218 16836 16218 0 _0211_
rlabel metal2 26450 26860 26450 26860 0 _0212_
rlabel metal2 19182 16558 19182 16558 0 _0213_
rlabel metal2 22310 10404 22310 10404 0 _0214_
rlabel metal2 20838 8772 20838 8772 0 _0215_
rlabel metal1 23782 19244 23782 19244 0 _0216_
rlabel metal1 23046 11186 23046 11186 0 _0217_
rlabel metal1 21114 10642 21114 10642 0 _0218_
rlabel metal1 22954 11730 22954 11730 0 _0219_
rlabel metal1 14996 10642 14996 10642 0 _0220_
rlabel metal1 25162 10234 25162 10234 0 _0221_
rlabel metal2 24610 14824 24610 14824 0 _0222_
rlabel metal2 14674 11900 14674 11900 0 _0223_
rlabel metal2 23414 13736 23414 13736 0 _0224_
rlabel metal1 20102 10778 20102 10778 0 _0225_
rlabel metal1 5152 11798 5152 11798 0 _0226_
rlabel metal1 4002 8398 4002 8398 0 _0227_
rlabel metal1 6072 13498 6072 13498 0 _0228_
rlabel metal2 6854 13464 6854 13464 0 _0229_
rlabel metal1 6394 10642 6394 10642 0 _0230_
rlabel metal2 8234 14756 8234 14756 0 _0231_
rlabel metal1 10074 35258 10074 35258 0 _0232_
rlabel metal2 10902 35972 10902 35972 0 _0233_
rlabel metal2 27462 36125 27462 36125 0 _0234_
rlabel via2 13386 35139 13386 35139 0 _0235_
rlabel metal1 8602 36346 8602 36346 0 _0236_
rlabel via1 22126 35989 22126 35989 0 _0237_
rlabel metal2 7682 15912 7682 15912 0 _0238_
rlabel metal2 26450 21114 26450 21114 0 _0239_
rlabel metal2 24794 23154 24794 23154 0 _0240_
rlabel metal2 23138 18122 23138 18122 0 _0241_
rlabel metal1 2346 9690 2346 9690 0 _0242_
rlabel metal2 11178 11288 11178 11288 0 _0243_
rlabel metal1 20194 30362 20194 30362 0 _0244_
rlabel metal2 18446 14382 18446 14382 0 _0245_
rlabel metal2 19918 21080 19918 21080 0 _0246_
rlabel metal1 24794 32776 24794 32776 0 _0247_
rlabel metal2 2898 27336 2898 27336 0 _0248_
rlabel metal2 25622 30906 25622 30906 0 _0249_
rlabel metal1 20286 23766 20286 23766 0 _0250_
rlabel metal1 20286 24854 20286 24854 0 _0251_
rlabel metal2 20010 11934 20010 11934 0 _0252_
rlabel metal1 26036 23494 26036 23494 0 _0253_
rlabel metal2 17434 10200 17434 10200 0 _0254_
rlabel metal1 30912 35802 30912 35802 0 _0255_
rlabel metal2 24426 22814 24426 22814 0 _0256_
rlabel metal1 26128 35802 26128 35802 0 _0257_
rlabel via2 19826 25211 19826 25211 0 _0258_
rlabel metal2 27370 27166 27370 27166 0 _0259_
rlabel metal2 28566 34816 28566 34816 0 _0260_
rlabel metal1 25852 34510 25852 34510 0 _0261_
rlabel metal1 25576 29206 25576 29206 0 _0262_
rlabel metal1 25806 28458 25806 28458 0 _0263_
rlabel metal1 13294 12614 13294 12614 0 _0264_
rlabel metal2 27738 14382 27738 14382 0 _0265_
rlabel metal1 15548 12138 15548 12138 0 _0266_
rlabel metal1 11178 13974 11178 13974 0 _0267_
rlabel metal2 19182 28662 19182 28662 0 _0268_
rlabel metal1 19826 14280 19826 14280 0 _0269_
rlabel metal2 23782 28798 23782 28798 0 _0270_
rlabel metal2 27738 30056 27738 30056 0 _0271_
rlabel metal1 24932 15402 24932 15402 0 _0272_
rlabel metal2 26082 30838 26082 30838 0 _0273_
rlabel metal1 21206 32334 21206 32334 0 _0274_
rlabel via1 24882 32470 24882 32470 0 _0275_
rlabel metal1 24288 35258 24288 35258 0 _0276_
rlabel metal1 28474 32538 28474 32538 0 _0277_
rlabel metal1 26680 27574 26680 27574 0 _0278_
rlabel metal2 24794 25738 24794 25738 0 _0279_
rlabel metal1 23920 23494 23920 23494 0 _0280_
rlabel metal1 28244 24582 28244 24582 0 _0281_
rlabel metal2 22770 23528 22770 23528 0 _0282_
rlabel metal1 27554 32538 27554 32538 0 _0283_
rlabel metal2 28014 21726 28014 21726 0 _0284_
rlabel metal2 30590 19550 30590 19550 0 _0285_
rlabel metal1 21482 24684 21482 24684 0 _0286_
rlabel metal1 10948 10778 10948 10778 0 _0287_
rlabel metal2 22678 16048 22678 16048 0 _0288_
rlabel metal2 24518 27710 24518 27710 0 _0289_
rlabel metal2 25714 29342 25714 29342 0 _0290_
rlabel metal1 23828 24854 23828 24854 0 _0291_
rlabel metal2 17066 16558 17066 16558 0 _0292_
rlabel metal2 24794 30328 24794 30328 0 _0293_
rlabel metal1 23184 16490 23184 16490 0 _0294_
rlabel metal1 19090 27370 19090 27370 0 _0295_
rlabel metal1 29072 34170 29072 34170 0 _0296_
rlabel metal1 24012 31994 24012 31994 0 _0297_
rlabel metal2 9430 14552 9430 14552 0 _0298_
rlabel metal2 10212 12852 10212 12852 0 _0299_
rlabel metal2 5474 11288 5474 11288 0 _0300_
rlabel metal1 19872 11050 19872 11050 0 _0301_
rlabel metal1 26496 22678 26496 22678 0 _0302_
rlabel metal2 26266 20808 26266 20808 0 _0303_
rlabel metal1 16928 15062 16928 15062 0 _0304_
rlabel metal1 28980 20502 28980 20502 0 _0305_
rlabel metal2 29026 19550 29026 19550 0 _0306_
rlabel metal2 9798 13464 9798 13464 0 _0307_
rlabel metal2 13386 13294 13386 13294 0 _0308_
rlabel metal2 26174 13532 26174 13532 0 _0309_
rlabel metal1 18354 14314 18354 14314 0 _0310_
rlabel metal1 16974 15368 16974 15368 0 _0311_
rlabel metal1 23368 12886 23368 12886 0 _0312_
rlabel metal1 24334 26554 24334 26554 0 _0313_
rlabel metal1 23046 25466 23046 25466 0 _0314_
rlabel metal1 7498 12614 7498 12614 0 _0315_
rlabel metal2 22954 15640 22954 15640 0 _0316_
rlabel metal1 20608 16150 20608 16150 0 _0317_
rlabel metal2 4738 14110 4738 14110 0 _0318_
rlabel metal1 13340 13498 13340 13498 0 _0319_
rlabel metal2 8234 10336 8234 10336 0 _0320_
rlabel metal1 5336 14586 5336 14586 0 _0321_
rlabel metal1 6256 15062 6256 15062 0 _0322_
rlabel metal2 2898 6664 2898 6664 0 _0323_
rlabel metal2 2990 13056 2990 13056 0 _0324_
rlabel metal1 21068 27098 21068 27098 0 _0325_
rlabel metal2 21942 24650 21942 24650 0 _0326_
rlabel metal2 18446 11934 18446 11934 0 _0327_
rlabel metal2 11546 15912 11546 15912 0 _0328_
rlabel metal2 24702 28390 24702 28390 0 _0329_
rlabel metal1 22080 12138 22080 12138 0 _0330_
rlabel metal1 6900 14314 6900 14314 0 _0331_
rlabel metal1 17848 12886 17848 12886 0 _0332_
rlabel metal1 21620 29546 21620 29546 0 _0333_
rlabel metal2 9338 36261 9338 36261 0 _0334_
rlabel metal2 3818 16014 3818 16014 0 _0335_
rlabel metal2 20562 20060 20562 20060 0 _0336_
rlabel metal2 10258 15470 10258 15470 0 _0337_
rlabel metal1 11224 33626 11224 33626 0 _0338_
rlabel metal1 6624 34714 6624 34714 0 _0339_
rlabel metal1 24150 25942 24150 25942 0 _0340_
rlabel metal1 22678 36074 22678 36074 0 _0341_
rlabel metal2 12742 34748 12742 34748 0 _0342_
rlabel metal2 24242 36873 24242 36873 0 _0343_
rlabel via2 26358 32555 26358 32555 0 _0344_
rlabel metal2 30498 36210 30498 36210 0 _0345_
rlabel metal1 19228 24718 19228 24718 0 _0346_
rlabel metal1 5980 14586 5980 14586 0 _0347_
rlabel metal2 19826 17884 19826 17884 0 _0348_
rlabel metal1 21620 28118 21620 28118 0 _0349_
rlabel metal1 21666 19414 21666 19414 0 _0350_
rlabel metal2 13938 29648 13938 29648 0 _0351_
rlabel metal2 22494 15810 22494 15810 0 _0352_
rlabel metal2 22034 15181 22034 15181 0 _0353_
rlabel metal1 4784 12886 4784 12886 0 _0354_
rlabel metal1 7130 12886 7130 12886 0 _0355_
rlabel metal1 19688 31790 19688 31790 0 _0356_
rlabel metal1 5106 16150 5106 16150 0 _0357_
rlabel metal3 1234 28628 1234 28628 0 ccff_head
rlabel metal1 6394 37094 6394 37094 0 ccff_tail
rlabel metal2 12926 1588 12926 1588 0 chanx_left_in[0]
rlabel metal2 19366 1588 19366 1588 0 chanx_left_in[10]
rlabel metal3 1188 26588 1188 26588 0 chanx_left_in[11]
rlabel metal3 1188 6868 1188 6868 0 chanx_left_in[12]
rlabel via2 37490 30685 37490 30685 0 chanx_left_in[13]
rlabel metal1 11684 2958 11684 2958 0 chanx_left_in[14]
rlabel metal1 27186 36176 27186 36176 0 chanx_left_in[15]
rlabel metal2 38134 8347 38134 8347 0 chanx_left_in[16]
rlabel metal3 1188 748 1188 748 0 chanx_left_in[17]
rlabel metal2 37490 35513 37490 35513 0 chanx_left_in[18]
rlabel metal3 1050 19108 1050 19108 0 chanx_left_in[1]
rlabel metal2 29946 35156 29946 35156 0 chanx_left_in[2]
rlabel metal3 1050 23188 1050 23188 0 chanx_left_in[3]
rlabel metal1 12328 37298 12328 37298 0 chanx_left_in[4]
rlabel metal1 37352 11118 37352 11118 0 chanx_left_in[5]
rlabel metal2 28382 1554 28382 1554 0 chanx_left_in[6]
rlabel metal1 4784 37230 4784 37230 0 chanx_left_in[7]
rlabel metal1 36202 37230 36202 37230 0 chanx_left_in[8]
rlabel metal1 37490 37230 37490 37230 0 chanx_left_in[9]
rlabel metal3 1234 5508 1234 5508 0 chanx_left_out[0]
rlabel metal2 20654 1520 20654 1520 0 chanx_left_out[10]
rlabel via2 38226 27931 38226 27931 0 chanx_left_out[11]
rlabel metal3 38740 12308 38740 12308 0 chanx_left_out[12]
rlabel metal1 15640 37094 15640 37094 0 chanx_left_out[13]
rlabel metal2 39330 2336 39330 2336 0 chanx_left_out[14]
rlabel metal1 33488 37094 33488 37094 0 chanx_left_out[15]
rlabel metal2 17434 1520 17434 1520 0 chanx_left_out[16]
rlabel metal1 3726 37094 3726 37094 0 chanx_left_out[17]
rlabel metal2 10994 1520 10994 1520 0 chanx_left_out[18]
rlabel metal3 1234 15708 1234 15708 0 chanx_left_out[1]
rlabel metal2 25162 1520 25162 1520 0 chanx_left_out[2]
rlabel metal2 38226 13073 38226 13073 0 chanx_left_out[3]
rlabel via2 38226 27285 38226 27285 0 chanx_left_out[4]
rlabel metal2 34822 1520 34822 1520 0 chanx_left_out[5]
rlabel metal2 14858 1520 14858 1520 0 chanx_left_out[6]
rlabel metal1 32752 36890 32752 36890 0 chanx_left_out[7]
rlabel metal1 20148 37094 20148 37094 0 chanx_left_out[8]
rlabel metal2 33534 1520 33534 1520 0 chanx_left_out[9]
rlabel metal2 38134 16439 38134 16439 0 chanx_right_in[0]
rlabel metal1 7866 37230 7866 37230 0 chanx_right_in[10]
rlabel metal2 38318 24021 38318 24021 0 chanx_right_in[11]
rlabel metal1 16330 36788 16330 36788 0 chanx_right_in[12]
rlabel metal2 38134 32759 38134 32759 0 chanx_right_in[13]
rlabel metal3 1188 4148 1188 4148 0 chanx_right_in[14]
rlabel metal2 38318 18003 38318 18003 0 chanx_right_in[15]
rlabel metal3 1234 31348 1234 31348 0 chanx_right_in[16]
rlabel metal3 1188 35428 1188 35428 0 chanx_right_in[17]
rlabel metal2 38318 32215 38318 32215 0 chanx_right_in[18]
rlabel metal2 37490 1921 37490 1921 0 chanx_right_in[1]
rlabel metal1 21666 37298 21666 37298 0 chanx_right_in[2]
rlabel metal1 17066 37196 17066 37196 0 chanx_right_in[3]
rlabel metal2 30958 38260 30958 38260 0 chanx_right_in[4]
rlabel metal2 38134 37145 38134 37145 0 chanx_right_in[5]
rlabel metal1 26312 37230 26312 37230 0 chanx_right_in[6]
rlabel metal2 9706 1588 9706 1588 0 chanx_right_in[7]
rlabel metal3 1188 17068 1188 17068 0 chanx_right_in[8]
rlabel metal3 1142 7548 1142 7548 0 chanx_right_in[9]
rlabel metal2 31602 1520 31602 1520 0 chanx_right_out[0]
rlabel metal2 38226 2057 38226 2057 0 chanx_right_out[10]
rlabel metal3 1234 15028 1234 15028 0 chanx_right_out[11]
rlabel metal2 38226 7633 38226 7633 0 chanx_right_out[12]
rlabel metal2 11086 37145 11086 37145 0 chanx_right_out[13]
rlabel metal2 1794 38131 1794 38131 0 chanx_right_out[14]
rlabel metal3 1234 21828 1234 21828 0 chanx_right_out[15]
rlabel metal2 16146 1520 16146 1520 0 chanx_right_out[16]
rlabel metal3 1234 25228 1234 25228 0 chanx_right_out[17]
rlabel metal1 34822 37094 34822 37094 0 chanx_right_out[18]
rlabel metal2 22586 1520 22586 1520 0 chanx_right_out[1]
rlabel metal2 29670 1520 29670 1520 0 chanx_right_out[2]
rlabel via2 38226 24565 38226 24565 0 chanx_right_out[3]
rlabel metal2 38226 4913 38226 4913 0 chanx_right_out[4]
rlabel metal1 27876 37094 27876 37094 0 chanx_right_out[5]
rlabel metal1 37352 36346 37352 36346 0 chanx_right_out[6]
rlabel metal1 17572 37094 17572 37094 0 chanx_right_out[7]
rlabel metal2 690 1792 690 1792 0 chanx_right_out[8]
rlabel metal2 5198 1520 5198 1520 0 chanx_right_out[9]
rlabel metal1 15134 37196 15134 37196 0 chany_top_in[0]
rlabel metal1 9798 36754 9798 36754 0 chany_top_in[10]
rlabel metal2 38318 21335 38318 21335 0 chany_top_in[11]
rlabel via2 38318 14365 38318 14365 0 chany_top_in[12]
rlabel metal1 38134 36754 38134 36754 0 chany_top_in[13]
rlabel metal1 3404 3026 3404 3026 0 chany_top_in[14]
rlabel metal2 37490 2873 37490 2873 0 chany_top_in[15]
rlabel metal2 38318 15895 38318 15895 0 chany_top_in[16]
rlabel metal3 1234 27268 1234 27268 0 chany_top_in[17]
rlabel metal2 2622 38209 2622 38209 0 chany_top_in[18]
rlabel metal2 36754 1894 36754 1894 0 chany_top_in[1]
rlabel metal3 1234 20468 1234 20468 0 chany_top_in[2]
rlabel metal1 920 36142 920 36142 0 chany_top_in[3]
rlabel metal1 36846 36176 36846 36176 0 chany_top_in[4]
rlabel metal2 8418 1588 8418 1588 0 chany_top_in[5]
rlabel metal3 1234 18428 1234 18428 0 chany_top_in[6]
rlabel metal2 23874 1588 23874 1588 0 chany_top_in[7]
rlabel metal2 38042 1367 38042 1367 0 chany_top_in[8]
rlabel metal1 14352 37230 14352 37230 0 chany_top_in[9]
rlabel metal2 30314 1520 30314 1520 0 chany_top_out[0]
rlabel metal2 3910 1520 3910 1520 0 chany_top_out[10]
rlabel metal3 1234 13668 1234 13668 0 chany_top_out[11]
rlabel metal2 38226 4301 38226 4301 0 chany_top_out[12]
rlabel metal2 38226 29393 38226 29393 0 chany_top_out[13]
rlabel metal2 32890 1520 32890 1520 0 chany_top_out[15]
rlabel metal3 1234 23868 1234 23868 0 chany_top_out[16]
rlabel metal2 38226 9741 38226 9741 0 chany_top_out[17]
rlabel metal3 1234 32028 1234 32028 0 chany_top_out[18]
rlabel via2 38226 22491 38226 22491 0 chany_top_out[1]
rlabel metal2 38226 34221 38226 34221 0 chany_top_out[2]
rlabel metal2 36110 1520 36110 1520 0 chany_top_out[3]
rlabel metal2 38226 36057 38226 36057 0 chany_top_out[4]
rlabel metal3 1234 33388 1234 33388 0 chany_top_out[5]
rlabel metal3 1602 2108 1602 2108 0 chany_top_out[6]
rlabel metal3 1234 12308 1234 12308 0 chany_top_out[7]
rlabel metal2 46 1656 46 1656 0 chany_top_out[8]
rlabel metal2 25806 1520 25806 1520 0 chany_top_out[9]
rlabel metal1 14720 21590 14720 21590 0 clknet_0_prog_clk
rlabel metal1 2484 20366 2484 20366 0 clknet_4_0_0_prog_clk
rlabel metal2 2714 33184 2714 33184 0 clknet_4_10_0_prog_clk
rlabel metal2 8970 33218 8970 33218 0 clknet_4_11_0_prog_clk
rlabel metal1 15088 31382 15088 31382 0 clknet_4_12_0_prog_clk
rlabel metal1 14352 27506 14352 27506 0 clknet_4_13_0_prog_clk
rlabel metal2 14674 35360 14674 35360 0 clknet_4_14_0_prog_clk
rlabel metal2 15962 32674 15962 32674 0 clknet_4_15_0_prog_clk
rlabel metal2 7314 17952 7314 17952 0 clknet_4_1_0_prog_clk
rlabel metal2 2438 23188 2438 23188 0 clknet_4_2_0_prog_clk
rlabel metal1 5796 21114 5796 21114 0 clknet_4_3_0_prog_clk
rlabel metal2 12006 17476 12006 17476 0 clknet_4_4_0_prog_clk
rlabel metal1 14536 21522 14536 21522 0 clknet_4_5_0_prog_clk
rlabel metal1 13340 20434 13340 20434 0 clknet_4_6_0_prog_clk
rlabel metal1 13938 23086 13938 23086 0 clknet_4_7_0_prog_clk
rlabel metal2 4002 27744 4002 27744 0 clknet_4_8_0_prog_clk
rlabel metal2 11270 27744 11270 27744 0 clknet_4_9_0_prog_clk
rlabel metal2 2898 37145 2898 37145 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 9982 37230 9982 37230 0 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 27370 37196 27370 37196 0 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1234 29988 1234 29988 0 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 6486 1588 6486 1588 0 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 1978 1894 1978 1894 0 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal1 1794 6732 1794 6732 0 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal1 19642 37196 19642 37196 0 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 18078 1588 18078 1588 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 35604 36754 35604 36754 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 10810 26095 10810 26095 0 mem_left_track_1.DFFR_0_.D
rlabel metal1 19780 21998 19780 21998 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 13662 17544 13662 17544 0 mem_left_track_1.DFFR_1_.Q
rlabel metal2 21666 26010 21666 26010 0 mem_left_track_1.DFFR_2_.Q
rlabel metal1 17526 12206 17526 12206 0 mem_left_track_1.DFFR_3_.Q
rlabel metal1 6348 20774 6348 20774 0 mem_left_track_1.DFFR_4_.Q
rlabel metal1 1978 19720 1978 19720 0 mem_left_track_1.DFFR_5_.Q
rlabel metal1 3542 19686 3542 19686 0 mem_left_track_1.DFFR_6_.Q
rlabel metal1 2438 12818 2438 12818 0 mem_left_track_1.DFFR_7_.Q
rlabel metal1 12788 35598 12788 35598 0 mem_left_track_17.DFFR_0_.D
rlabel metal2 14214 34833 14214 34833 0 mem_left_track_17.DFFR_0_.Q
rlabel metal3 10787 16116 10787 16116 0 mem_left_track_17.DFFR_1_.Q
rlabel metal2 16054 34085 16054 34085 0 mem_left_track_17.DFFR_2_.Q
rlabel metal2 12650 34748 12650 34748 0 mem_left_track_17.DFFR_3_.Q
rlabel metal1 15410 34680 15410 34680 0 mem_left_track_17.DFFR_4_.Q
rlabel metal1 3496 35258 3496 35258 0 mem_left_track_17.DFFR_5_.Q
rlabel metal1 4554 17850 4554 17850 0 mem_left_track_17.DFFR_6_.Q
rlabel metal1 19090 20502 19090 20502 0 mem_left_track_17.DFFR_7_.Q
rlabel metal2 16560 27370 16560 27370 0 mem_left_track_25.DFFR_0_.Q
rlabel metal1 21068 15470 21068 15470 0 mem_left_track_25.DFFR_1_.Q
rlabel metal1 20654 19346 20654 19346 0 mem_left_track_25.DFFR_2_.Q
rlabel metal1 3956 14382 3956 14382 0 mem_left_track_25.DFFR_3_.Q
rlabel metal2 5382 25500 5382 25500 0 mem_left_track_25.DFFR_4_.Q
rlabel metal2 17526 24633 17526 24633 0 mem_left_track_25.DFFR_5_.Q
rlabel metal2 7360 18292 7360 18292 0 mem_left_track_25.DFFR_6_.Q
rlabel metal1 13662 18122 13662 18122 0 mem_left_track_25.DFFR_7_.Q
rlabel via2 13754 27013 13754 27013 0 mem_left_track_33.DFFR_0_.Q
rlabel metal1 17158 32776 17158 32776 0 mem_left_track_33.DFFR_1_.Q
rlabel metal1 17158 32504 17158 32504 0 mem_left_track_33.DFFR_2_.Q
rlabel metal1 18630 32300 18630 32300 0 mem_left_track_33.DFFR_3_.Q
rlabel metal1 19734 32368 19734 32368 0 mem_left_track_33.DFFR_4_.Q
rlabel metal1 13156 20502 13156 20502 0 mem_left_track_9.DFFR_0_.Q
rlabel metal1 14582 13872 14582 13872 0 mem_left_track_9.DFFR_1_.Q
rlabel metal1 12742 13974 12742 13974 0 mem_left_track_9.DFFR_2_.Q
rlabel metal1 17204 29206 17204 29206 0 mem_left_track_9.DFFR_3_.Q
rlabel metal1 18400 29070 18400 29070 0 mem_left_track_9.DFFR_4_.Q
rlabel metal2 13294 34850 13294 34850 0 mem_right_track_0.DFFR_0_.D
rlabel metal1 22494 32878 22494 32878 0 mem_right_track_0.DFFR_0_.Q
rlabel via2 2622 9571 2622 9571 0 mem_right_track_0.DFFR_1_.Q
rlabel metal1 20654 17204 20654 17204 0 mem_right_track_0.DFFR_2_.Q
rlabel metal1 15778 21386 15778 21386 0 mem_right_track_0.DFFR_3_.Q
rlabel metal1 8096 16626 8096 16626 0 mem_right_track_0.DFFR_4_.Q
rlabel metal1 13846 22032 13846 22032 0 mem_right_track_0.DFFR_5_.Q
rlabel metal1 19458 16592 19458 16592 0 mem_right_track_16.DFFR_0_.D
rlabel metal1 18952 19482 18952 19482 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 16698 16592 16698 16592 0 mem_right_track_16.DFFR_1_.Q
rlabel metal2 18354 19414 18354 19414 0 mem_right_track_16.DFFR_2_.Q
rlabel metal1 17158 19482 17158 19482 0 mem_right_track_16.DFFR_3_.Q
rlabel metal2 15226 17238 15226 17238 0 mem_right_track_16.DFFR_4_.Q
rlabel metal1 10304 17102 10304 17102 0 mem_right_track_16.DFFR_5_.Q
rlabel metal2 11178 17510 11178 17510 0 mem_right_track_16.DFFR_6_.Q
rlabel metal1 4922 19890 4922 19890 0 mem_right_track_16.DFFR_7_.Q
rlabel metal1 5474 14382 5474 14382 0 mem_right_track_24.DFFR_0_.Q
rlabel metal2 18814 15776 18814 15776 0 mem_right_track_24.DFFR_1_.Q
rlabel metal2 17250 22984 17250 22984 0 mem_right_track_24.DFFR_2_.Q
rlabel metal1 7406 21454 7406 21454 0 mem_right_track_24.DFFR_3_.Q
rlabel metal2 12742 13396 12742 13396 0 mem_right_track_24.DFFR_4_.Q
rlabel metal2 13570 18326 13570 18326 0 mem_right_track_24.DFFR_5_.Q
rlabel metal1 13202 18938 13202 18938 0 mem_right_track_24.DFFR_6_.Q
rlabel metal1 15548 18938 15548 18938 0 mem_right_track_24.DFFR_7_.Q
rlabel metal1 14950 29070 14950 29070 0 mem_right_track_32.DFFR_0_.Q
rlabel metal1 17250 10642 17250 10642 0 mem_right_track_32.DFFR_1_.Q
rlabel metal1 17296 30294 17296 30294 0 mem_right_track_32.DFFR_2_.Q
rlabel metal2 18078 26452 18078 26452 0 mem_right_track_32.DFFR_3_.Q
rlabel metal2 18262 25466 18262 25466 0 mem_right_track_32.DFFR_4_.Q
rlabel metal1 14260 33014 14260 33014 0 mem_right_track_8.DFFR_0_.Q
rlabel metal1 16008 17170 16008 17170 0 mem_right_track_8.DFFR_1_.Q
rlabel metal1 17434 27982 17434 27982 0 mem_right_track_8.DFFR_2_.Q
rlabel metal1 17664 25806 17664 25806 0 mem_right_track_8.DFFR_3_.Q
rlabel metal2 18630 25568 18630 25568 0 mem_right_track_8.DFFR_4_.Q
rlabel metal2 16514 24140 16514 24140 0 mem_right_track_8.DFFR_5_.Q
rlabel metal2 14766 22576 14766 22576 0 mem_right_track_8.DFFR_6_.Q
rlabel metal2 5198 13804 5198 13804 0 mem_top_track_0.DFFR_0_.Q
rlabel metal1 3680 20366 3680 20366 0 mem_top_track_0.DFFR_1_.Q
rlabel metal2 2622 12036 2622 12036 0 mem_top_track_0.DFFR_2_.Q
rlabel metal1 6670 17544 6670 17544 0 mem_top_track_0.DFFR_3_.Q
rlabel metal1 7866 17510 7866 17510 0 mem_top_track_0.DFFR_4_.Q
rlabel metal1 15042 12206 15042 12206 0 mem_top_track_0.DFFR_5_.Q
rlabel metal2 15594 35394 15594 35394 0 mem_top_track_10.DFFR_0_.D
rlabel metal2 18538 35734 18538 35734 0 mem_top_track_10.DFFR_0_.Q
rlabel metal1 12742 35224 12742 35224 0 mem_top_track_10.DFFR_1_.Q
rlabel metal2 15686 13413 15686 13413 0 mem_top_track_12.DFFR_0_.Q
rlabel metal1 7314 18326 7314 18326 0 mem_top_track_12.DFFR_1_.Q
rlabel metal2 17618 17272 17618 17272 0 mem_top_track_14.DFFR_0_.Q
rlabel metal1 4462 17714 4462 17714 0 mem_top_track_14.DFFR_1_.Q
rlabel metal1 6394 17850 6394 17850 0 mem_top_track_16.DFFR_0_.Q
rlabel metal1 7636 18190 7636 18190 0 mem_top_track_16.DFFR_1_.Q
rlabel metal1 22126 11730 22126 11730 0 mem_top_track_18.DFFR_0_.Q
rlabel metal1 22540 11118 22540 11118 0 mem_top_track_18.DFFR_1_.Q
rlabel metal1 17158 21624 17158 21624 0 mem_top_track_2.DFFR_0_.Q
rlabel metal1 18584 21318 18584 21318 0 mem_top_track_2.DFFR_1_.Q
rlabel metal1 20562 18292 20562 18292 0 mem_top_track_2.DFFR_2_.Q
rlabel metal1 20240 23834 20240 23834 0 mem_top_track_2.DFFR_3_.Q
rlabel metal1 18216 24038 18216 24038 0 mem_top_track_2.DFFR_4_.Q
rlabel metal2 14582 27948 14582 27948 0 mem_top_track_2.DFFR_5_.Q
rlabel metal1 16606 18734 16606 18734 0 mem_top_track_20.DFFR_0_.Q
rlabel metal1 15272 11730 15272 11730 0 mem_top_track_20.DFFR_1_.Q
rlabel metal1 4738 18190 4738 18190 0 mem_top_track_22.DFFR_0_.Q
rlabel metal2 6026 18768 6026 18768 0 mem_top_track_22.DFFR_1_.Q
rlabel metal2 14398 10812 14398 10812 0 mem_top_track_24.DFFR_0_.Q
rlabel metal1 25070 11730 25070 11730 0 mem_top_track_24.DFFR_1_.Q
rlabel metal2 15318 19210 15318 19210 0 mem_top_track_26.DFFR_0_.Q
rlabel metal1 13018 19788 13018 19788 0 mem_top_track_26.DFFR_1_.Q
rlabel metal1 19918 36142 19918 36142 0 mem_top_track_36.DFFR_0_.Q
rlabel metal1 17066 36686 17066 36686 0 mem_top_track_4.DFFR_0_.Q
rlabel via1 17894 36550 17894 36550 0 mem_top_track_4.DFFR_1_.Q
rlabel metal2 18630 34510 18630 34510 0 mem_top_track_4.DFFR_2_.Q
rlabel metal1 17204 35598 17204 35598 0 mem_top_track_4.DFFR_3_.Q
rlabel via2 21022 35445 21022 35445 0 mem_top_track_4.DFFR_4_.Q
rlabel metal1 18630 33286 18630 33286 0 mem_top_track_4.DFFR_5_.Q
rlabel metal2 16422 35734 16422 35734 0 mem_top_track_6.DFFR_0_.Q
rlabel metal1 16836 32810 16836 32810 0 mem_top_track_6.DFFR_1_.Q
rlabel metal2 24150 32640 24150 32640 0 mem_top_track_6.DFFR_2_.Q
rlabel metal1 17296 31382 17296 31382 0 mem_top_track_6.DFFR_3_.Q
rlabel metal2 18630 29920 18630 29920 0 mem_top_track_6.DFFR_4_.Q
rlabel metal2 16698 29274 16698 29274 0 mem_top_track_6.DFFR_5_.Q
rlabel metal1 15732 34442 15732 34442 0 mem_top_track_8.DFFR_0_.Q
rlabel metal2 20654 34952 20654 34952 0 mux_left_track_1.INVTX1_0_.out
rlabel metal1 16974 15980 16974 15980 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 28014 36550 28014 36550 0 mux_left_track_1.INVTX1_2_.out
rlabel metal1 22356 12274 22356 12274 0 mux_left_track_1.INVTX1_3_.out
rlabel metal1 16698 12750 16698 12750 0 mux_left_track_1.INVTX1_4_.out
rlabel metal1 22724 33286 22724 33286 0 mux_left_track_1.INVTX1_5_.out
rlabel metal1 23368 14926 23368 14926 0 mux_left_track_1.INVTX1_6_.out
rlabel metal1 18722 10778 18722 10778 0 mux_left_track_1.INVTX1_7_.out
rlabel metal1 1932 22950 1932 22950 0 mux_left_track_1.INVTX1_8_.out
rlabel metal1 22678 12138 22678 12138 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 19918 23494 19918 23494 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 7360 14314 7360 14314 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 1794 10234 1794 10234 0 mux_left_track_1.out
rlabel via2 7774 36533 7774 36533 0 mux_left_track_17.INVTX1_0_.out
rlabel metal1 26174 11254 26174 11254 0 mux_left_track_17.INVTX1_1_.out
rlabel metal1 25898 36040 25898 36040 0 mux_left_track_17.INVTX1_2_.out
rlabel metal2 9522 36057 9522 36057 0 mux_left_track_17.INVTX1_3_.out
rlabel metal2 21114 34918 21114 34918 0 mux_left_track_17.INVTX1_4_.out
rlabel metal1 9706 9146 9706 9146 0 mux_left_track_17.INVTX1_5_.out
rlabel metal1 8556 31926 8556 31926 0 mux_left_track_17.INVTX1_6_.out
rlabel metal2 6486 36380 6486 36380 0 mux_left_track_17.INVTX1_7_.out
rlabel metal1 2622 14926 2622 14926 0 mux_left_track_17.INVTX1_8_.out
rlabel metal1 25162 36686 25162 36686 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 11316 15062 11316 15062 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 20930 17408 20930 17408 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 20930 36890 20930 36890 0 mux_left_track_17.out
rlabel metal2 4186 16422 4186 16422 0 mux_left_track_25.INVTX1_0_.out
rlabel metal1 22862 15368 22862 15368 0 mux_left_track_25.INVTX1_1_.out
rlabel metal2 21942 15436 21942 15436 0 mux_left_track_25.INVTX1_2_.out
rlabel metal1 2530 13838 2530 13838 0 mux_left_track_25.INVTX1_3_.out
rlabel metal1 25070 31858 25070 31858 0 mux_left_track_25.INVTX1_4_.out
rlabel metal1 20654 11832 20654 11832 0 mux_left_track_25.INVTX1_5_.out
rlabel metal1 18722 16014 18722 16014 0 mux_left_track_25.INVTX1_6_.out
rlabel metal1 16008 30090 16008 30090 0 mux_left_track_25.INVTX1_7_.out
rlabel metal1 2116 8602 2116 8602 0 mux_left_track_25.INVTX1_8_.out
rlabel metal2 17986 14450 17986 14450 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 21896 31858 21896 31858 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 20838 15436 20838 15436 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 37720 12206 37720 12206 0 mux_left_track_25.out
rlabel metal1 31418 9622 31418 9622 0 mux_left_track_33.INVTX1_0_.out
rlabel metal2 21850 15793 21850 15793 0 mux_left_track_33.INVTX1_1_.out
rlabel metal1 29072 20978 29072 20978 0 mux_left_track_33.INVTX1_2_.out
rlabel metal1 28842 19278 28842 19278 0 mux_left_track_33.INVTX1_3_.out
rlabel metal1 27554 28492 27554 28492 0 mux_left_track_33.INVTX1_4_.out
rlabel metal1 20378 34918 20378 34918 0 mux_left_track_33.INVTX1_5_.out
rlabel metal1 28428 34034 28428 34034 0 mux_left_track_33.INVTX1_6_.out
rlabel metal1 25162 35802 25162 35802 0 mux_left_track_33.INVTX1_7_.out
rlabel metal2 24058 20162 24058 20162 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 28014 21386 28014 21386 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 24886 32334 24886 32334 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 21942 9554 21942 9554 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 19136 7854 19136 7854 0 mux_left_track_33.out
rlabel metal1 26496 30158 26496 30158 0 mux_left_track_9.INVTX1_0_.out
rlabel metal1 19872 34918 19872 34918 0 mux_left_track_9.INVTX1_1_.out
rlabel metal1 17434 13838 17434 13838 0 mux_left_track_9.INVTX1_2_.out
rlabel metal1 23920 15402 23920 15402 0 mux_left_track_9.INVTX1_3_.out
rlabel metal1 15502 13362 15502 13362 0 mux_left_track_9.INVTX1_4_.out
rlabel metal1 11500 13838 11500 13838 0 mux_left_track_9.INVTX1_5_.out
rlabel metal1 28152 29682 28152 29682 0 mux_left_track_9.INVTX1_6_.out
rlabel metal1 13018 10234 13018 10234 0 mux_left_track_9.INVTX1_7_.out
rlabel metal2 23690 15317 23690 15317 0 mux_left_track_9.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 21620 12410 21620 12410 0 mux_left_track_9.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 23230 11424 23230 11424 0 mux_left_track_9.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 28474 29206 28474 29206 0 mux_left_track_9.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 31510 28730 31510 28730 0 mux_left_track_9.out
rlabel metal2 2438 29104 2438 29104 0 mux_right_track_0.INVTX1_3_.out
rlabel metal2 2392 8772 2392 8772 0 mux_right_track_0.INVTX1_4_.out
rlabel metal1 11454 9486 11454 9486 0 mux_right_track_0.INVTX1_5_.out
rlabel via1 23966 33558 23966 33558 0 mux_right_track_0.INVTX1_6_.out
rlabel metal2 23460 21420 23460 21420 0 mux_right_track_0.INVTX1_7_.out
rlabel metal2 19826 20910 19826 20910 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 6808 12580 6808 12580 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 25806 20842 25806 20842 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 27140 8466 27140 8466 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 29072 7854 29072 7854 0 mux_right_track_0.out
rlabel metal1 11868 12750 11868 12750 0 mux_right_track_16.INVTX1_4_.out
rlabel metal1 19964 10234 19964 10234 0 mux_right_track_16.INVTX1_5_.out
rlabel metal1 27324 33830 27324 33830 0 mux_right_track_16.INVTX1_6_.out
rlabel metal1 26496 20366 26496 20366 0 mux_right_track_16.INVTX1_7_.out
rlabel metal1 11868 13294 11868 13294 0 mux_right_track_16.INVTX1_8_.out
rlabel metal2 17250 14212 17250 14212 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 12558 13600 12558 13600 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 10258 13838 10258 13838 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 4738 5372 4738 5372 0 mux_right_track_16.out
rlabel metal1 6210 9554 6210 9554 0 mux_right_track_24.INVTX1_4_.out
rlabel metal1 23782 28594 23782 28594 0 mux_right_track_24.INVTX1_5_.out
rlabel metal1 25024 33410 25024 33410 0 mux_right_track_24.INVTX1_6_.out
rlabel metal1 8602 12274 8602 12274 0 mux_right_track_24.INVTX1_7_.out
rlabel metal2 16882 14994 16882 14994 0 mux_right_track_24.INVTX1_8_.out
rlabel metal2 15318 14076 15318 14076 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 17802 14314 17802 14314 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 31878 11356 31878 11356 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 32614 9996 32614 9996 0 mux_right_track_24.out
rlabel metal2 14858 9010 14858 9010 0 mux_right_track_32.INVTX1_4_.out
rlabel metal1 31326 36210 31326 36210 0 mux_right_track_32.INVTX1_5_.out
rlabel metal1 28934 27302 28934 27302 0 mux_right_track_32.INVTX1_6_.out
rlabel metal1 20746 10574 20746 10574 0 mux_right_track_32.INVTX1_7_.out
rlabel metal1 26818 36074 26818 36074 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 19412 10098 19412 10098 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 20654 11628 20654 11628 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 21160 12308 21160 12308 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 17020 7174 17020 7174 0 mux_right_track_32.out
rlabel via2 14674 36091 14674 36091 0 mux_right_track_8.INVTX1_4_.out
rlabel metal1 24426 26860 24426 26860 0 mux_right_track_8.INVTX1_5_.out
rlabel metal1 25576 24786 25576 24786 0 mux_right_track_8.INVTX1_6_.out
rlabel metal2 20746 23800 20746 23800 0 mux_right_track_8.INVTX1_7_.out
rlabel metal1 8372 11594 8372 11594 0 mux_right_track_8.INVTX1_8_.out
rlabel metal2 20102 16218 20102 16218 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 26772 33796 26772 33796 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 23966 11186 23966 11186 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 34960 6766 34960 6766 0 mux_right_track_8.out
rlabel metal1 23092 11662 23092 11662 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 19780 12138 19780 12138 0 mux_top_track_0.INVTX1_1_.out
rlabel metal1 9844 9486 9844 9486 0 mux_top_track_0.INVTX1_3_.out
rlabel metal2 2346 10540 2346 10540 0 mux_top_track_0.INVTX1_5_.out
rlabel metal1 17526 10472 17526 10472 0 mux_top_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 8464 10574 8464 10574 0 mux_top_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 20217 5678 20217 5678 0 mux_top_track_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 24794 5372 24794 5372 0 mux_top_track_0.out
rlabel metal1 24702 34068 24702 34068 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel via2 6210 32861 6210 32861 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 4738 33082 4738 33082 0 mux_top_track_10.out
rlabel metal1 21436 24174 21436 24174 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 6808 12410 6808 12410 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 6164 8942 6164 8942 0 mux_top_track_12.out
rlabel metal1 6578 15538 6578 15538 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 3128 14586 3128 14586 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 4646 13838 4646 13838 0 mux_top_track_14.out
rlabel metal1 8372 11526 8372 11526 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 3542 9520 3542 9520 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 3956 7378 3956 7378 0 mux_top_track_16.out
rlabel metal1 24288 11866 24288 11866 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 21206 10064 21206 10064 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 23874 9996 23874 9996 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 24794 8330 24794 8330 0 mux_top_track_18.out
rlabel metal1 21988 18258 21988 18258 0 mux_top_track_2.INVTX1_1_.out
rlabel metal1 27002 23630 27002 23630 0 mux_top_track_2.INVTX1_3_.out
rlabel metal2 25530 24208 25530 24208 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal2 22770 19346 22770 19346 0 mux_top_track_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 24748 19890 24748 19890 0 mux_top_track_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 36110 22916 36110 22916 0 mux_top_track_2.out
rlabel metal1 22540 12342 22540 12342 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 25346 10880 25346 10880 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15272 10438 15272 10438 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 12466 8092 12466 8092 0 mux_top_track_20.out
rlabel metal1 7728 14042 7728 14042 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 5290 11662 5290 11662 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 2714 11662 2714 11662 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 2116 11118 2116 11118 0 mux_top_track_22.out
rlabel metal2 22862 11866 22862 11866 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 25714 11968 25714 11968 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 34776 7378 34776 7378 0 mux_top_track_24.out
rlabel metal2 19366 16252 19366 16252 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 29210 26758 29210 26758 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 31602 27268 31602 27268 0 mux_top_track_26.out
rlabel metal1 24426 35700 24426 35700 0 mux_top_track_36.INVTX1_1_.out
rlabel metal1 7820 36686 7820 36686 0 mux_top_track_36.INVTX1_2_.out
rlabel metal1 26036 35530 26036 35530 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9246 36074 9246 36074 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 9844 36210 9844 36210 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 7176 32742 7176 32742 0 mux_top_track_36.out
rlabel metal2 29854 21760 29854 21760 0 mux_top_track_4.INVTX1_2_.out
rlabel metal2 21206 35156 21206 35156 0 mux_top_track_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 36869 35054 36869 35054 0 mux_top_track_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 38042 34442 38042 34442 0 mux_top_track_4.out
rlabel metal2 29854 26962 29854 26962 0 mux_top_track_6.INVTX1_0_.out
rlabel metal1 28244 32946 28244 32946 0 mux_top_track_6.INVTX1_2_.out
rlabel metal1 28336 31858 28336 31858 0 mux_top_track_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 32660 4590 32660 4590 0 mux_top_track_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 34408 4590 34408 4590 0 mux_top_track_6.out
rlabel metal2 28198 28832 28198 28832 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 28014 29648 28014 29648 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 35098 30736 35098 30736 0 mux_top_track_8.out
rlabel metal1 1738 27642 1738 27642 0 net1
rlabel metal2 1794 2142 1794 2142 0 net10
rlabel metal1 14950 2380 14950 2380 0 net100
rlabel metal2 33074 36550 33074 36550 0 net101
rlabel metal1 20470 37230 20470 37230 0 net102
rlabel metal2 24886 6460 24886 6460 0 net103
rlabel metal1 32016 2414 32016 2414 0 net104
rlabel metal1 37950 3570 37950 3570 0 net105
rlabel metal1 1610 15436 1610 15436 0 net106
rlabel metal2 34178 8330 34178 8330 0 net107
rlabel metal1 14214 28730 14214 28730 0 net108
rlabel metal1 1978 37230 1978 37230 0 net109
rlabel metal2 37720 19108 37720 19108 0 net11
rlabel metal1 1978 17306 1978 17306 0 net110
rlabel metal2 16882 2618 16882 2618 0 net111
rlabel metal3 1679 24956 1679 24956 0 net112
rlabel metal1 34868 37230 34868 37230 0 net113
rlabel metal1 22678 2448 22678 2448 0 net114
rlabel metal1 29302 20230 29302 20230 0 net115
rlabel metal2 38042 24548 38042 24548 0 net116
rlabel metal2 38042 5916 38042 5916 0 net117
rlabel metal1 27508 36890 27508 36890 0 net118
rlabel metal1 37858 36074 37858 36074 0 net119
rlabel metal1 15042 20264 15042 20264 0 net12
rlabel metal1 17664 37230 17664 37230 0 net120
rlabel metal1 1610 3060 1610 3060 0 net121
rlabel metal1 5290 2448 5290 2448 0 net122
rlabel metal2 30498 3706 30498 3706 0 net123
rlabel metal1 5428 2346 5428 2346 0 net124
rlabel metal1 1702 11322 1702 11322 0 net125
rlabel metal1 37904 4590 37904 4590 0 net126
rlabel metal2 36662 28594 36662 28594 0 net127
rlabel metal1 33212 2414 33212 2414 0 net128
rlabel metal1 1932 24174 1932 24174 0 net129
rlabel metal1 29532 34918 29532 34918 0 net13
rlabel metal2 36478 9724 36478 9724 0 net130
rlabel metal1 1610 32368 1610 32368 0 net131
rlabel metal2 38042 22780 38042 22780 0 net132
rlabel metal2 37858 34374 37858 34374 0 net133
rlabel metal2 35374 3434 35374 3434 0 net134
rlabel metal1 37720 36142 37720 36142 0 net135
rlabel metal1 1610 33558 1610 33558 0 net136
rlabel metal1 2898 2346 2898 2346 0 net137
rlabel metal2 2070 12070 2070 12070 0 net138
rlabel metal1 3910 2482 3910 2482 0 net139
rlabel metal1 2162 24582 2162 24582 0 net14
rlabel metal1 25300 7718 25300 7718 0 net140
rlabel metal2 38318 20689 38318 20689 0 net141
rlabel metal2 15226 5984 15226 5984 0 net142
rlabel metal2 29946 25568 29946 25568 0 net143
rlabel metal1 30314 35598 30314 35598 0 net144
rlabel metal2 31142 23392 31142 23392 0 net145
rlabel metal1 28060 30226 28060 30226 0 net146
rlabel metal2 5566 33184 5566 33184 0 net147
rlabel metal1 8418 10098 8418 10098 0 net148
rlabel metal1 2254 13362 2254 13362 0 net149
rlabel metal2 18446 36584 18446 36584 0 net15
rlabel metal2 2898 8636 2898 8636 0 net150
rlabel metal2 27002 11424 27002 11424 0 net151
rlabel metal1 28658 26010 28658 26010 0 net152
rlabel metal2 20470 9248 20470 9248 0 net153
rlabel metal2 24702 11424 24702 11424 0 net154
rlabel metal1 4324 8466 4324 8466 0 net155
rlabel metal2 10442 36448 10442 36448 0 net156
rlabel metal1 25254 18802 25254 18802 0 net157
rlabel metal1 26174 22066 26174 22066 0 net158
rlabel metal2 27646 14110 27646 14110 0 net159
rlabel metal1 37490 11220 37490 11220 0 net16
rlabel metal1 28934 33592 28934 33592 0 net160
rlabel metal2 26174 15776 26174 15776 0 net161
rlabel metal2 5382 10914 5382 10914 0 net162
rlabel metal1 23368 12274 23368 12274 0 net163
rlabel metal1 2990 12274 2990 12274 0 net164
rlabel metal2 20378 19652 20378 19652 0 net165
rlabel metal1 19596 17306 19596 17306 0 net166
rlabel metal1 28060 2618 28060 2618 0 net17
rlabel metal1 6394 36754 6394 36754 0 net18
rlabel metal2 36386 31756 36386 31756 0 net19
rlabel metal1 18906 3060 18906 3060 0 net2
rlabel metal2 37628 26220 37628 26220 0 net20
rlabel metal2 38226 15062 38226 15062 0 net21
rlabel metal2 8050 31212 8050 31212 0 net22
rlabel metal1 37996 24378 37996 24378 0 net23
rlabel metal2 20194 35564 20194 35564 0 net24
rlabel metal2 37904 26220 37904 26220 0 net25
rlabel metal2 16238 14552 16238 14552 0 net26
rlabel metal1 37398 18394 37398 18394 0 net27
rlabel metal1 3588 31790 3588 31790 0 net28
rlabel metal1 1656 35462 1656 35462 0 net29
rlabel metal1 10764 2482 10764 2482 0 net3
rlabel metal2 33074 33252 33074 33252 0 net30
rlabel metal2 37306 2788 37306 2788 0 net31
rlabel metal1 26634 21522 26634 21522 0 net32
rlabel metal2 19274 36533 19274 36533 0 net33
rlabel metal2 31786 28288 31786 28288 0 net34
rlabel metal1 37766 36550 37766 36550 0 net35
rlabel metal1 23046 36754 23046 36754 0 net36
rlabel metal1 10028 2618 10028 2618 0 net37
rlabel via3 2645 16660 2645 16660 0 net38
rlabel metal2 9154 8432 9154 8432 0 net39
rlabel via3 1909 26452 1909 26452 0 net4
rlabel metal2 14950 36992 14950 36992 0 net40
rlabel metal2 10350 36397 10350 36397 0 net41
rlabel metal2 29762 21114 29762 21114 0 net42
rlabel metal1 37352 14586 37352 14586 0 net43
rlabel metal2 36754 35564 36754 35564 0 net44
rlabel metal1 7268 2890 7268 2890 0 net45
rlabel metal1 37030 2992 37030 2992 0 net46
rlabel metal1 37950 16218 37950 16218 0 net47
rlabel via3 2277 9588 2277 9588 0 net48
rlabel metal1 2714 37128 2714 37128 0 net49
rlabel metal2 12926 8942 12926 8942 0 net5
rlabel metal1 35512 3162 35512 3162 0 net50
rlabel metal2 2254 19482 2254 19482 0 net51
rlabel metal2 7682 36516 7682 36516 0 net52
rlabel metal1 35604 36006 35604 36006 0 net53
rlabel metal1 9154 2312 9154 2312 0 net54
rlabel metal1 1610 17544 1610 17544 0 net55
rlabel metal1 24656 2618 24656 2618 0 net56
rlabel metal1 32706 3366 32706 3366 0 net57
rlabel metal2 19458 35564 19458 35564 0 net58
rlabel metal2 4738 36550 4738 36550 0 net59
rlabel metal1 37766 30838 37766 30838 0 net6
rlabel metal1 12834 36584 12834 36584 0 net60
rlabel metal2 28934 36108 28934 36108 0 net61
rlabel metal1 1932 23086 1932 23086 0 net62
rlabel metal2 9062 2176 9062 2176 0 net63
rlabel metal2 4002 5508 4002 5508 0 net64
rlabel metal1 1886 6630 1886 6630 0 net65
rlabel metal1 25484 35666 25484 35666 0 net66
rlabel metal1 18630 10574 18630 10574 0 net67
rlabel metal1 34132 36618 34132 36618 0 net68
rlabel metal1 25369 6222 25369 6222 0 net69
rlabel metal1 2530 17136 2530 17136 0 net7
rlabel metal2 6854 9588 6854 9588 0 net70
rlabel metal1 7176 2618 7176 2618 0 net71
rlabel metal1 14536 2618 14536 2618 0 net72
rlabel metal1 1932 3706 1932 3706 0 net73
rlabel metal2 30406 26996 30406 26996 0 net74
rlabel metal1 20930 10030 20930 10030 0 net75
rlabel metal2 32062 33014 32062 33014 0 net76
rlabel metal2 32338 35700 32338 35700 0 net77
rlabel metal1 1748 36550 1748 36550 0 net78
rlabel metal2 6118 37094 6118 37094 0 net79
rlabel metal1 32430 36686 32430 36686 0 net8
rlabel metal1 26772 2618 26772 2618 0 net80
rlabel metal1 3910 9520 3910 9520 0 net81
rlabel metal2 3358 34884 3358 34884 0 net82
rlabel metal1 37904 19482 37904 19482 0 net83
rlabel metal2 17802 30702 17802 30702 0 net84
rlabel metal1 1564 5678 1564 5678 0 net85
rlabel metal1 20378 2414 20378 2414 0 net86
rlabel metal2 38042 27268 38042 27268 0 net87
rlabel metal1 37950 12410 37950 12410 0 net88
rlabel metal1 21988 36890 21988 36890 0 net89
rlabel metal2 13294 10268 13294 10268 0 net9
rlabel metal1 37996 4114 37996 4114 0 net90
rlabel metal2 33626 26044 33626 26044 0 net91
rlabel metal1 18124 7718 18124 7718 0 net92
rlabel metal2 2990 34612 2990 34612 0 net93
rlabel metal1 10534 4998 10534 4998 0 net94
rlabel metal2 7222 14722 7222 14722 0 net95
rlabel metal2 25254 2618 25254 2618 0 net96
rlabel metal1 38042 13362 38042 13362 0 net97
rlabel metal2 33074 27914 33074 27914 0 net98
rlabel metal1 33258 2550 33258 2550 0 net99
rlabel via2 37490 6205 37490 6205 0 pReset
rlabel metal3 2108 36788 2108 36788 0 prog_clk
rlabel metal1 1794 8976 1794 8976 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 7130 1588 7130 1588 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 14214 1588 14214 1588 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1234 3468 1234 3468 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 38786 25908 38786 25908 0 right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 21942 1588 21942 1588 0 right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal1 31970 35530 31970 35530 0 right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal1 31234 35088 31234 35088 0 right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal1 1564 36754 1564 36754 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 6256 37230 6256 37230 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 27094 1588 27094 1588 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 2806 9911 2806 9911 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 1234 34748 1234 34748 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 38318 19227 38318 19227 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
