// This is the unpowered netlist.
module sb_1__1_ (bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
    bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    ccff_head,
    ccff_tail,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    pReset,
    prog_clk,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    chanx_left_in,
    chanx_left_out,
    chanx_right_in,
    chanx_right_out,
    chany_bottom_in,
    chany_bottom_out,
    chany_top_in,
    chany_top_out);
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input ccff_head;
 output ccff_tail;
 input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input pReset;
 input prog_clk;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input [0:18] chanx_left_in;
 output [0:18] chanx_left_out;
 input [0:18] chanx_right_in;
 output [0:18] chanx_right_out;
 input [0:18] chany_bottom_in;
 output [0:18] chany_bottom_out;
 input [0:18] chany_top_in;
 output [0:18] chany_top_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire clknet_0_prog_clk;
 wire \mem_bottom_track_1.DFFR_0_.D ;
 wire \mem_bottom_track_1.DFFR_0_.Q ;
 wire \mem_bottom_track_1.DFFR_1_.Q ;
 wire \mem_bottom_track_1.DFFR_2_.Q ;
 wire \mem_bottom_track_1.DFFR_3_.Q ;
 wire \mem_bottom_track_1.DFFR_4_.Q ;
 wire \mem_bottom_track_1.DFFR_5_.Q ;
 wire \mem_bottom_track_1.DFFR_6_.Q ;
 wire \mem_bottom_track_1.DFFR_7_.Q ;
 wire \mem_bottom_track_17.DFFR_0_.D ;
 wire \mem_bottom_track_17.DFFR_0_.Q ;
 wire \mem_bottom_track_17.DFFR_1_.Q ;
 wire \mem_bottom_track_17.DFFR_2_.Q ;
 wire \mem_bottom_track_17.DFFR_3_.Q ;
 wire \mem_bottom_track_17.DFFR_4_.Q ;
 wire \mem_bottom_track_17.DFFR_5_.Q ;
 wire \mem_bottom_track_17.DFFR_6_.Q ;
 wire \mem_bottom_track_17.DFFR_7_.Q ;
 wire \mem_bottom_track_25.DFFR_0_.Q ;
 wire \mem_bottom_track_25.DFFR_1_.Q ;
 wire \mem_bottom_track_25.DFFR_2_.Q ;
 wire \mem_bottom_track_25.DFFR_3_.Q ;
 wire \mem_bottom_track_25.DFFR_4_.Q ;
 wire \mem_bottom_track_25.DFFR_5_.Q ;
 wire \mem_bottom_track_25.DFFR_6_.Q ;
 wire \mem_bottom_track_25.DFFR_7_.Q ;
 wire \mem_bottom_track_33.DFFR_0_.Q ;
 wire \mem_bottom_track_33.DFFR_1_.Q ;
 wire \mem_bottom_track_33.DFFR_2_.Q ;
 wire \mem_bottom_track_33.DFFR_3_.Q ;
 wire \mem_bottom_track_33.DFFR_4_.Q ;
 wire \mem_bottom_track_33.DFFR_5_.Q ;
 wire \mem_bottom_track_9.DFFR_0_.Q ;
 wire \mem_bottom_track_9.DFFR_1_.Q ;
 wire \mem_bottom_track_9.DFFR_2_.Q ;
 wire \mem_bottom_track_9.DFFR_3_.Q ;
 wire \mem_bottom_track_9.DFFR_4_.Q ;
 wire \mem_bottom_track_9.DFFR_5_.Q ;
 wire \mem_bottom_track_9.DFFR_6_.Q ;
 wire \mem_left_track_1.DFFR_0_.Q ;
 wire \mem_left_track_1.DFFR_1_.Q ;
 wire \mem_left_track_1.DFFR_2_.Q ;
 wire \mem_left_track_1.DFFR_3_.Q ;
 wire \mem_left_track_1.DFFR_4_.Q ;
 wire \mem_left_track_1.DFFR_5_.Q ;
 wire \mem_left_track_1.DFFR_6_.Q ;
 wire \mem_left_track_1.DFFR_7_.Q ;
 wire \mem_left_track_17.DFFR_0_.D ;
 wire \mem_left_track_17.DFFR_0_.Q ;
 wire \mem_left_track_17.DFFR_1_.Q ;
 wire \mem_left_track_17.DFFR_2_.Q ;
 wire \mem_left_track_17.DFFR_3_.Q ;
 wire \mem_left_track_17.DFFR_4_.Q ;
 wire \mem_left_track_17.DFFR_5_.Q ;
 wire \mem_left_track_17.DFFR_6_.Q ;
 wire \mem_left_track_17.DFFR_7_.Q ;
 wire \mem_left_track_25.DFFR_0_.Q ;
 wire \mem_left_track_25.DFFR_1_.Q ;
 wire \mem_left_track_25.DFFR_2_.Q ;
 wire \mem_left_track_25.DFFR_3_.Q ;
 wire \mem_left_track_25.DFFR_4_.Q ;
 wire \mem_left_track_25.DFFR_5_.Q ;
 wire \mem_left_track_25.DFFR_6_.Q ;
 wire \mem_left_track_25.DFFR_7_.Q ;
 wire \mem_left_track_33.DFFR_0_.Q ;
 wire \mem_left_track_33.DFFR_1_.Q ;
 wire \mem_left_track_33.DFFR_2_.Q ;
 wire \mem_left_track_33.DFFR_3_.Q ;
 wire \mem_left_track_33.DFFR_4_.Q ;
 wire \mem_left_track_9.DFFR_0_.Q ;
 wire \mem_left_track_9.DFFR_1_.Q ;
 wire \mem_left_track_9.DFFR_2_.Q ;
 wire \mem_left_track_9.DFFR_3_.Q ;
 wire \mem_left_track_9.DFFR_4_.Q ;
 wire \mem_left_track_9.DFFR_5_.Q ;
 wire \mem_left_track_9.DFFR_6_.Q ;
 wire \mem_right_track_0.DFFR_0_.D ;
 wire \mem_right_track_0.DFFR_0_.Q ;
 wire \mem_right_track_0.DFFR_1_.Q ;
 wire \mem_right_track_0.DFFR_2_.Q ;
 wire \mem_right_track_0.DFFR_3_.Q ;
 wire \mem_right_track_0.DFFR_4_.Q ;
 wire \mem_right_track_0.DFFR_5_.Q ;
 wire \mem_right_track_0.DFFR_6_.Q ;
 wire \mem_right_track_0.DFFR_7_.Q ;
 wire \mem_right_track_16.DFFR_0_.D ;
 wire \mem_right_track_16.DFFR_0_.Q ;
 wire \mem_right_track_16.DFFR_1_.Q ;
 wire \mem_right_track_16.DFFR_2_.Q ;
 wire \mem_right_track_16.DFFR_3_.Q ;
 wire \mem_right_track_16.DFFR_4_.Q ;
 wire \mem_right_track_16.DFFR_5_.Q ;
 wire \mem_right_track_16.DFFR_6_.Q ;
 wire \mem_right_track_16.DFFR_7_.Q ;
 wire \mem_right_track_24.DFFR_0_.Q ;
 wire \mem_right_track_24.DFFR_1_.Q ;
 wire \mem_right_track_24.DFFR_2_.Q ;
 wire \mem_right_track_24.DFFR_3_.Q ;
 wire \mem_right_track_24.DFFR_4_.Q ;
 wire \mem_right_track_24.DFFR_5_.Q ;
 wire \mem_right_track_24.DFFR_6_.Q ;
 wire \mem_right_track_24.DFFR_7_.Q ;
 wire \mem_right_track_32.DFFR_0_.Q ;
 wire \mem_right_track_32.DFFR_1_.Q ;
 wire \mem_right_track_32.DFFR_2_.Q ;
 wire \mem_right_track_32.DFFR_3_.Q ;
 wire \mem_right_track_32.DFFR_4_.Q ;
 wire \mem_right_track_8.DFFR_0_.Q ;
 wire \mem_right_track_8.DFFR_1_.Q ;
 wire \mem_right_track_8.DFFR_2_.Q ;
 wire \mem_right_track_8.DFFR_3_.Q ;
 wire \mem_right_track_8.DFFR_4_.Q ;
 wire \mem_right_track_8.DFFR_5_.Q ;
 wire \mem_right_track_8.DFFR_6_.Q ;
 wire \mem_top_track_0.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_1_.Q ;
 wire \mem_top_track_0.DFFR_2_.Q ;
 wire \mem_top_track_0.DFFR_3_.Q ;
 wire \mem_top_track_0.DFFR_4_.Q ;
 wire \mem_top_track_0.DFFR_5_.Q ;
 wire \mem_top_track_0.DFFR_6_.Q ;
 wire \mem_top_track_0.DFFR_7_.Q ;
 wire \mem_top_track_16.DFFR_0_.D ;
 wire \mem_top_track_16.DFFR_0_.Q ;
 wire \mem_top_track_16.DFFR_1_.Q ;
 wire \mem_top_track_16.DFFR_2_.Q ;
 wire \mem_top_track_16.DFFR_3_.Q ;
 wire \mem_top_track_16.DFFR_4_.Q ;
 wire \mem_top_track_16.DFFR_5_.Q ;
 wire \mem_top_track_16.DFFR_6_.Q ;
 wire \mem_top_track_16.DFFR_7_.Q ;
 wire \mem_top_track_24.DFFR_0_.Q ;
 wire \mem_top_track_24.DFFR_1_.Q ;
 wire \mem_top_track_24.DFFR_2_.Q ;
 wire \mem_top_track_24.DFFR_3_.Q ;
 wire \mem_top_track_24.DFFR_4_.Q ;
 wire \mem_top_track_24.DFFR_5_.Q ;
 wire \mem_top_track_24.DFFR_6_.Q ;
 wire \mem_top_track_24.DFFR_7_.Q ;
 wire \mem_top_track_32.DFFR_0_.Q ;
 wire \mem_top_track_32.DFFR_1_.Q ;
 wire \mem_top_track_32.DFFR_2_.Q ;
 wire \mem_top_track_32.DFFR_3_.Q ;
 wire \mem_top_track_32.DFFR_4_.Q ;
 wire \mem_top_track_8.DFFR_0_.Q ;
 wire \mem_top_track_8.DFFR_1_.Q ;
 wire \mem_top_track_8.DFFR_2_.Q ;
 wire \mem_top_track_8.DFFR_3_.Q ;
 wire \mem_top_track_8.DFFR_4_.Q ;
 wire \mem_top_track_8.DFFR_5_.Q ;
 wire \mem_top_track_8.DFFR_6_.Q ;
 wire \mux_bottom_track_1.INVTX1_0_.out ;
 wire \mux_bottom_track_1.INVTX1_10_.out ;
 wire \mux_bottom_track_1.INVTX1_11_.out ;
 wire \mux_bottom_track_1.INVTX1_1_.out ;
 wire \mux_bottom_track_1.INVTX1_2_.out ;
 wire \mux_bottom_track_1.INVTX1_3_.out ;
 wire \mux_bottom_track_1.INVTX1_4_.out ;
 wire \mux_bottom_track_1.INVTX1_5_.out ;
 wire \mux_bottom_track_1.INVTX1_6_.out ;
 wire \mux_bottom_track_1.INVTX1_7_.out ;
 wire \mux_bottom_track_1.INVTX1_8_.out ;
 wire \mux_bottom_track_1.INVTX1_9_.out ;
 wire \mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_bottom_track_1.out ;
 wire \mux_bottom_track_17.INVTX1_0_.out ;
 wire \mux_bottom_track_17.INVTX1_10_.out ;
 wire \mux_bottom_track_17.INVTX1_11_.out ;
 wire \mux_bottom_track_17.INVTX1_1_.out ;
 wire \mux_bottom_track_17.INVTX1_2_.out ;
 wire \mux_bottom_track_17.INVTX1_3_.out ;
 wire \mux_bottom_track_17.INVTX1_4_.out ;
 wire \mux_bottom_track_17.INVTX1_5_.out ;
 wire \mux_bottom_track_17.INVTX1_6_.out ;
 wire \mux_bottom_track_17.INVTX1_7_.out ;
 wire \mux_bottom_track_17.INVTX1_8_.out ;
 wire \mux_bottom_track_17.INVTX1_9_.out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_bottom_track_17.out ;
 wire \mux_bottom_track_25.INVTX1_0_.out ;
 wire \mux_bottom_track_25.INVTX1_10_.out ;
 wire \mux_bottom_track_25.INVTX1_11_.out ;
 wire \mux_bottom_track_25.INVTX1_1_.out ;
 wire \mux_bottom_track_25.INVTX1_2_.out ;
 wire \mux_bottom_track_25.INVTX1_3_.out ;
 wire \mux_bottom_track_25.INVTX1_4_.out ;
 wire \mux_bottom_track_25.INVTX1_5_.out ;
 wire \mux_bottom_track_25.INVTX1_6_.out ;
 wire \mux_bottom_track_25.INVTX1_7_.out ;
 wire \mux_bottom_track_25.INVTX1_8_.out ;
 wire \mux_bottom_track_25.INVTX1_9_.out ;
 wire \mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_bottom_track_25.out ;
 wire \mux_bottom_track_33.INVTX1_0_.out ;
 wire \mux_bottom_track_33.INVTX1_1_.out ;
 wire \mux_bottom_track_33.INVTX1_2_.out ;
 wire \mux_bottom_track_33.INVTX1_3_.out ;
 wire \mux_bottom_track_33.INVTX1_4_.out ;
 wire \mux_bottom_track_33.INVTX1_5_.out ;
 wire \mux_bottom_track_33.INVTX1_6_.out ;
 wire \mux_bottom_track_33.INVTX1_7_.out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_bottom_track_33.out ;
 wire \mux_bottom_track_9.INVTX1_0_.out ;
 wire \mux_bottom_track_9.INVTX1_10_.out ;
 wire \mux_bottom_track_9.INVTX1_11_.out ;
 wire \mux_bottom_track_9.INVTX1_1_.out ;
 wire \mux_bottom_track_9.INVTX1_2_.out ;
 wire \mux_bottom_track_9.INVTX1_3_.out ;
 wire \mux_bottom_track_9.INVTX1_4_.out ;
 wire \mux_bottom_track_9.INVTX1_5_.out ;
 wire \mux_bottom_track_9.INVTX1_6_.out ;
 wire \mux_bottom_track_9.INVTX1_7_.out ;
 wire \mux_bottom_track_9.INVTX1_8_.out ;
 wire \mux_bottom_track_9.INVTX1_9_.out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_bottom_track_9.out ;
 wire \mux_left_track_1.INVTX1_10_.out ;
 wire \mux_left_track_1.INVTX1_11_.out ;
 wire \mux_left_track_1.INVTX1_1_.out ;
 wire \mux_left_track_1.INVTX1_7_.out ;
 wire \mux_left_track_1.INVTX1_8_.out ;
 wire \mux_left_track_1.INVTX1_9_.out ;
 wire \mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_left_track_1.out ;
 wire \mux_left_track_17.INVTX1_10_.out ;
 wire \mux_left_track_17.INVTX1_11_.out ;
 wire \mux_left_track_17.INVTX1_2_.out ;
 wire \mux_left_track_17.INVTX1_7_.out ;
 wire \mux_left_track_17.INVTX1_8_.out ;
 wire \mux_left_track_17.INVTX1_9_.out ;
 wire \mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_left_track_17.out ;
 wire \mux_left_track_25.INVTX1_10_.out ;
 wire \mux_left_track_25.INVTX1_11_.out ;
 wire \mux_left_track_25.INVTX1_2_.out ;
 wire \mux_left_track_25.INVTX1_7_.out ;
 wire \mux_left_track_25.INVTX1_8_.out ;
 wire \mux_left_track_25.INVTX1_9_.out ;
 wire \mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_left_track_25.out ;
 wire \mux_left_track_33.INVTX1_1_.out ;
 wire \mux_left_track_33.INVTX1_5_.out ;
 wire \mux_left_track_33.INVTX1_6_.out ;
 wire \mux_left_track_33.INVTX1_7_.out ;
 wire \mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_left_track_33.out ;
 wire \mux_left_track_9.INVTX1_10_.out ;
 wire \mux_left_track_9.INVTX1_11_.out ;
 wire \mux_left_track_9.INVTX1_3_.out ;
 wire \mux_left_track_9.INVTX1_7_.out ;
 wire \mux_left_track_9.INVTX1_8_.out ;
 wire \mux_left_track_9.INVTX1_9_.out ;
 wire \mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_left_track_9.out ;
 wire \mux_right_track_0.INVTX1_4_.out ;
 wire \mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_right_track_0.out ;
 wire \mux_right_track_16.INVTX1_4_.out ;
 wire \mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_right_track_16.out ;
 wire \mux_right_track_24.INVTX1_4_.out ;
 wire \mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_right_track_24.out ;
 wire \mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_right_track_32.out ;
 wire \mux_right_track_8.INVTX1_4_.out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_right_track_8.out ;
 wire \mux_top_track_0.INVTX1_0_.out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_top_track_0.out ;
 wire \mux_top_track_16.INVTX1_0_.out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_top_track_16.out ;
 wire \mux_top_track_24.INVTX1_0_.out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_top_track_24.out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_top_track_32.out ;
 wire \mux_top_track_8.INVTX1_0_.out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ;
 wire \mux_top_track_8.out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire clknet_4_0_0_prog_clk;
 wire clknet_4_1_0_prog_clk;
 wire clknet_4_2_0_prog_clk;
 wire clknet_4_3_0_prog_clk;
 wire clknet_4_4_0_prog_clk;
 wire clknet_4_5_0_prog_clk;
 wire clknet_4_6_0_prog_clk;
 wire clknet_4_7_0_prog_clk;
 wire clknet_4_8_0_prog_clk;
 wire clknet_4_9_0_prog_clk;
 wire clknet_4_10_0_prog_clk;
 wire clknet_4_11_0_prog_clk;
 wire clknet_4_12_0_prog_clk;
 wire clknet_4_13_0_prog_clk;
 wire clknet_4_14_0_prog_clk;
 wire clknet_4_15_0_prog_clk;

 sky130_fd_sc_hd__inv_2 _0493_ (.A(\mem_left_track_33.DFFR_3_.Q ),
    .Y(_0469_));
 sky130_fd_sc_hd__inv_2 _0494_ (.A(\mem_left_track_33.DFFR_0_.Q ),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_2 _0495_ (.A(\mem_left_track_33.DFFR_2_.Q ),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _0496_ (.A(\mem_left_track_33.DFFR_1_.Q ),
    .Y(_0467_));
 sky130_fd_sc_hd__inv_2 _0497_ (.A(net95),
    .Y(_0462_));
 sky130_fd_sc_hd__inv_2 _0498_ (.A(\mem_left_track_33.DFFR_0_.Q ),
    .Y(_0470_));
 sky130_fd_sc_hd__inv_2 _0499_ (.A(\mem_left_track_33.DFFR_2_.Q ),
    .Y(_0464_));
 sky130_fd_sc_hd__inv_2 _0500_ (.A(\mem_left_track_33.DFFR_1_.Q ),
    .Y(_0463_));
 sky130_fd_sc_hd__inv_2 _0501_ (.A(\mem_left_track_33.DFFR_4_.Q ),
    .Y(_0461_));
 sky130_fd_sc_hd__inv_2 _0502_ (.A(\mem_left_track_33.DFFR_0_.Q ),
    .Y(_0471_));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(\mem_left_track_33.DFFR_2_.Q ),
    .Y(_0466_));
 sky130_fd_sc_hd__inv_2 _0504_ (.A(\mem_left_track_33.DFFR_1_.Q ),
    .Y(_0465_));
 sky130_fd_sc_hd__inv_2 _0505_ (.A(\mem_bottom_track_33.DFFR_3_.Q ),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _0506_ (.A(\mem_bottom_track_33.DFFR_0_.Q ),
    .Y(_0460_));
 sky130_fd_sc_hd__inv_2 _0507_ (.A(\mem_bottom_track_33.DFFR_2_.Q ),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _0508_ (.A(\mem_bottom_track_33.DFFR_1_.Q ),
    .Y(_0455_));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(\mem_bottom_track_33.DFFR_5_.Q ),
    .Y(_0450_));
 sky130_fd_sc_hd__inv_2 _0510_ (.A(\mem_bottom_track_33.DFFR_0_.Q ),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_2 _0511_ (.A(\mem_bottom_track_33.DFFR_2_.Q ),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_2 _0512_ (.A(\mem_bottom_track_33.DFFR_1_.Q ),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _0513_ (.A(\mem_bottom_track_33.DFFR_4_.Q ),
    .Y(_0449_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(\mem_bottom_track_33.DFFR_0_.Q ),
    .Y(_0459_));
 sky130_fd_sc_hd__inv_2 _0515_ (.A(\mem_bottom_track_33.DFFR_2_.Q ),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _0516_ (.A(\mem_bottom_track_33.DFFR_1_.Q ),
    .Y(_0453_));
 sky130_fd_sc_hd__inv_2 _0517_ (.A(\mem_right_track_32.DFFR_3_.Q ),
    .Y(_0445_));
 sky130_fd_sc_hd__inv_2 _0518_ (.A(\mem_right_track_32.DFFR_0_.Q ),
    .Y(_0448_));
 sky130_fd_sc_hd__inv_2 _0519_ (.A(\mem_right_track_32.DFFR_2_.Q ),
    .Y(_0444_));
 sky130_fd_sc_hd__inv_2 _0520_ (.A(\mem_right_track_32.DFFR_1_.Q ),
    .Y(_0443_));
 sky130_fd_sc_hd__inv_2 _0521_ (.A(\mem_bottom_track_1.DFFR_0_.D ),
    .Y(_0438_));
 sky130_fd_sc_hd__inv_2 _0522_ (.A(\mem_right_track_32.DFFR_0_.Q ),
    .Y(_0446_));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(\mem_right_track_32.DFFR_2_.Q ),
    .Y(_0440_));
 sky130_fd_sc_hd__inv_2 _0524_ (.A(\mem_right_track_32.DFFR_1_.Q ),
    .Y(_0439_));
 sky130_fd_sc_hd__inv_2 _0525_ (.A(\mem_right_track_32.DFFR_4_.Q ),
    .Y(_0437_));
 sky130_fd_sc_hd__inv_2 _0526_ (.A(\mem_right_track_32.DFFR_0_.Q ),
    .Y(_0447_));
 sky130_fd_sc_hd__inv_2 _0527_ (.A(\mem_right_track_32.DFFR_2_.Q ),
    .Y(_0442_));
 sky130_fd_sc_hd__inv_2 _0528_ (.A(\mem_right_track_32.DFFR_1_.Q ),
    .Y(_0441_));
 sky130_fd_sc_hd__inv_2 _0529_ (.A(\mem_top_track_32.DFFR_3_.Q ),
    .Y(_0433_));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(\mem_top_track_32.DFFR_0_.Q ),
    .Y(_0436_));
 sky130_fd_sc_hd__inv_2 _0531_ (.A(\mem_top_track_32.DFFR_2_.Q ),
    .Y(_0432_));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(\mem_top_track_32.DFFR_1_.Q ),
    .Y(_0431_));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(\mem_right_track_0.DFFR_0_.D ),
    .Y(_0426_));
 sky130_fd_sc_hd__inv_2 _0534_ (.A(\mem_top_track_32.DFFR_0_.Q ),
    .Y(_0434_));
 sky130_fd_sc_hd__inv_2 _0535_ (.A(\mem_top_track_32.DFFR_2_.Q ),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_2 _0536_ (.A(\mem_top_track_32.DFFR_1_.Q ),
    .Y(_0427_));
 sky130_fd_sc_hd__inv_2 _0537_ (.A(\mem_top_track_32.DFFR_4_.Q ),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_2 _0538_ (.A(\mem_top_track_32.DFFR_0_.Q ),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_2 _0539_ (.A(\mem_top_track_32.DFFR_2_.Q ),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_2 _0540_ (.A(\mem_top_track_32.DFFR_1_.Q ),
    .Y(_0429_));
 sky130_fd_sc_hd__inv_2 _0541_ (.A(\mem_left_track_25.DFFR_4_.Q ),
    .Y(_0421_));
 sky130_fd_sc_hd__inv_2 _0542_ (.A(\mem_left_track_25.DFFR_0_.Q ),
    .Y(_0424_));
 sky130_fd_sc_hd__inv_2 _0543_ (.A(\mem_left_track_25.DFFR_3_.Q ),
    .Y(_0420_));
 sky130_fd_sc_hd__inv_2 _0544_ (.A(\mem_left_track_25.DFFR_2_.Q ),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_2 _0545_ (.A(\mem_left_track_25.DFFR_1_.Q ),
    .Y(_0418_));
 sky130_fd_sc_hd__inv_2 _0546_ (.A(\mem_left_track_25.DFFR_7_.Q ),
    .Y(_0411_));
 sky130_fd_sc_hd__inv_2 _0547_ (.A(\mem_left_track_25.DFFR_6_.Q ),
    .Y(_0410_));
 sky130_fd_sc_hd__inv_2 _0548_ (.A(\mem_left_track_25.DFFR_0_.Q ),
    .Y(_0422_));
 sky130_fd_sc_hd__inv_2 _0549_ (.A(\mem_left_track_25.DFFR_3_.Q ),
    .Y(_0414_));
 sky130_fd_sc_hd__inv_2 _0550_ (.A(\mem_left_track_25.DFFR_2_.Q ),
    .Y(_0413_));
 sky130_fd_sc_hd__inv_2 _0551_ (.A(\mem_left_track_25.DFFR_1_.Q ),
    .Y(_0412_));
 sky130_fd_sc_hd__inv_2 _0552_ (.A(\mem_left_track_25.DFFR_5_.Q ),
    .Y(_0409_));
 sky130_fd_sc_hd__inv_2 _0553_ (.A(\mem_left_track_25.DFFR_0_.Q ),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_2 _0554_ (.A(\mem_left_track_25.DFFR_3_.Q ),
    .Y(_0417_));
 sky130_fd_sc_hd__inv_2 _0555_ (.A(\mem_left_track_25.DFFR_2_.Q ),
    .Y(_0416_));
 sky130_fd_sc_hd__inv_2 _0556_ (.A(\mem_left_track_25.DFFR_1_.Q ),
    .Y(_0415_));
 sky130_fd_sc_hd__inv_2 _0557_ (.A(\mem_left_track_17.DFFR_4_.Q ),
    .Y(_0405_));
 sky130_fd_sc_hd__inv_2 _0558_ (.A(\mem_left_track_17.DFFR_0_.Q ),
    .Y(_0408_));
 sky130_fd_sc_hd__inv_2 _0559_ (.A(\mem_left_track_17.DFFR_3_.Q ),
    .Y(_0404_));
 sky130_fd_sc_hd__inv_2 _0560_ (.A(\mem_left_track_17.DFFR_2_.Q ),
    .Y(_0403_));
 sky130_fd_sc_hd__inv_2 _0561_ (.A(\mem_left_track_17.DFFR_1_.Q ),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _0562_ (.A(\mem_left_track_17.DFFR_7_.Q ),
    .Y(_0395_));
 sky130_fd_sc_hd__inv_2 _0563_ (.A(\mem_left_track_17.DFFR_6_.Q ),
    .Y(_0394_));
 sky130_fd_sc_hd__inv_2 _0564_ (.A(\mem_left_track_17.DFFR_0_.Q ),
    .Y(_0406_));
 sky130_fd_sc_hd__inv_2 _0565_ (.A(\mem_left_track_17.DFFR_3_.Q ),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_2 _0566_ (.A(\mem_left_track_17.DFFR_2_.Q ),
    .Y(_0397_));
 sky130_fd_sc_hd__inv_2 _0567_ (.A(\mem_left_track_17.DFFR_1_.Q ),
    .Y(_0396_));
 sky130_fd_sc_hd__inv_2 _0568_ (.A(\mem_left_track_17.DFFR_5_.Q ),
    .Y(_0393_));
 sky130_fd_sc_hd__inv_2 _0569_ (.A(\mem_left_track_17.DFFR_0_.Q ),
    .Y(_0407_));
 sky130_fd_sc_hd__inv_2 _0570_ (.A(\mem_left_track_17.DFFR_3_.Q ),
    .Y(_0401_));
 sky130_fd_sc_hd__inv_2 _0571_ (.A(\mem_left_track_17.DFFR_2_.Q ),
    .Y(_0400_));
 sky130_fd_sc_hd__inv_2 _0572_ (.A(\mem_left_track_17.DFFR_1_.Q ),
    .Y(_0399_));
 sky130_fd_sc_hd__inv_2 _0573_ (.A(\mem_left_track_9.DFFR_4_.Q ),
    .Y(_0389_));
 sky130_fd_sc_hd__inv_2 _0574_ (.A(\mem_left_track_9.DFFR_0_.Q ),
    .Y(_0392_));
 sky130_fd_sc_hd__inv_2 _0575_ (.A(\mem_left_track_9.DFFR_3_.Q ),
    .Y(_0388_));
 sky130_fd_sc_hd__inv_2 _0576_ (.A(\mem_left_track_9.DFFR_2_.Q ),
    .Y(_0387_));
 sky130_fd_sc_hd__inv_2 _0577_ (.A(\mem_left_track_9.DFFR_1_.Q ),
    .Y(_0386_));
 sky130_fd_sc_hd__inv_2 _0578_ (.A(\mem_left_track_17.DFFR_0_.D ),
    .Y(_0379_));
 sky130_fd_sc_hd__inv_2 _0579_ (.A(\mem_left_track_9.DFFR_6_.Q ),
    .Y(_0378_));
 sky130_fd_sc_hd__inv_2 _0580_ (.A(\mem_left_track_9.DFFR_0_.Q ),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_2 _0581_ (.A(\mem_left_track_9.DFFR_3_.Q ),
    .Y(_0382_));
 sky130_fd_sc_hd__inv_2 _0582_ (.A(\mem_left_track_9.DFFR_2_.Q ),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_2 _0583_ (.A(\mem_left_track_9.DFFR_1_.Q ),
    .Y(_0380_));
 sky130_fd_sc_hd__inv_2 _0584_ (.A(\mem_left_track_9.DFFR_5_.Q ),
    .Y(_0377_));
 sky130_fd_sc_hd__inv_2 _0585_ (.A(\mem_left_track_9.DFFR_0_.Q ),
    .Y(_0391_));
 sky130_fd_sc_hd__inv_2 _0586_ (.A(\mem_left_track_9.DFFR_3_.Q ),
    .Y(_0385_));
 sky130_fd_sc_hd__inv_2 _0587_ (.A(\mem_left_track_9.DFFR_2_.Q ),
    .Y(_0384_));
 sky130_fd_sc_hd__inv_2 _0588_ (.A(\mem_left_track_9.DFFR_1_.Q ),
    .Y(_0383_));
 sky130_fd_sc_hd__inv_2 _0589_ (.A(\mem_left_track_1.DFFR_4_.Q ),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _0590_ (.A(\mem_left_track_1.DFFR_0_.Q ),
    .Y(_0376_));
 sky130_fd_sc_hd__inv_2 _0591_ (.A(\mem_left_track_1.DFFR_3_.Q ),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _0592_ (.A(\mem_left_track_1.DFFR_2_.Q ),
    .Y(_0371_));
 sky130_fd_sc_hd__inv_2 _0593_ (.A(\mem_left_track_1.DFFR_1_.Q ),
    .Y(_0370_));
 sky130_fd_sc_hd__inv_2 _0594_ (.A(\mem_left_track_1.DFFR_7_.Q ),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_2 _0595_ (.A(\mem_left_track_1.DFFR_6_.Q ),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_2 _0596_ (.A(\mem_left_track_1.DFFR_0_.Q ),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _0597_ (.A(\mem_left_track_1.DFFR_3_.Q ),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_2 _0598_ (.A(\mem_left_track_1.DFFR_2_.Q ),
    .Y(_0365_));
 sky130_fd_sc_hd__inv_2 _0599_ (.A(\mem_left_track_1.DFFR_1_.Q ),
    .Y(_0364_));
 sky130_fd_sc_hd__inv_2 _0600_ (.A(\mem_left_track_1.DFFR_5_.Q ),
    .Y(_0361_));
 sky130_fd_sc_hd__inv_2 _0601_ (.A(\mem_left_track_1.DFFR_0_.Q ),
    .Y(_0375_));
 sky130_fd_sc_hd__inv_2 _0602_ (.A(\mem_left_track_1.DFFR_3_.Q ),
    .Y(_0369_));
 sky130_fd_sc_hd__inv_2 _0603_ (.A(\mem_left_track_1.DFFR_2_.Q ),
    .Y(_0368_));
 sky130_fd_sc_hd__inv_2 _0604_ (.A(\mem_left_track_1.DFFR_1_.Q ),
    .Y(_0367_));
 sky130_fd_sc_hd__inv_2 _0605_ (.A(\mem_bottom_track_25.DFFR_4_.Q ),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _0606_ (.A(\mem_bottom_track_25.DFFR_0_.Q ),
    .Y(_0360_));
 sky130_fd_sc_hd__inv_2 _0607_ (.A(\mem_bottom_track_25.DFFR_3_.Q ),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _0608_ (.A(\mem_bottom_track_25.DFFR_2_.Q ),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_2 _0609_ (.A(\mem_bottom_track_25.DFFR_1_.Q ),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _0610_ (.A(\mem_bottom_track_25.DFFR_7_.Q ),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _0611_ (.A(\mem_bottom_track_25.DFFR_6_.Q ),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _0612_ (.A(\mem_bottom_track_25.DFFR_0_.Q ),
    .Y(_0358_));
 sky130_fd_sc_hd__inv_2 _0613_ (.A(\mem_bottom_track_25.DFFR_3_.Q ),
    .Y(_0350_));
 sky130_fd_sc_hd__inv_2 _0614_ (.A(\mem_bottom_track_25.DFFR_2_.Q ),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _0615_ (.A(\mem_bottom_track_25.DFFR_1_.Q ),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _0616_ (.A(\mem_bottom_track_25.DFFR_5_.Q ),
    .Y(_0345_));
 sky130_fd_sc_hd__inv_2 _0617_ (.A(\mem_bottom_track_25.DFFR_0_.Q ),
    .Y(_0359_));
 sky130_fd_sc_hd__inv_2 _0618_ (.A(\mem_bottom_track_25.DFFR_3_.Q ),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_2 _0619_ (.A(\mem_bottom_track_25.DFFR_2_.Q ),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_2 _0620_ (.A(\mem_bottom_track_25.DFFR_1_.Q ),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _0621_ (.A(\mem_bottom_track_17.DFFR_4_.Q ),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _0622_ (.A(\mem_bottom_track_17.DFFR_0_.Q ),
    .Y(_0344_));
 sky130_fd_sc_hd__inv_2 _0623_ (.A(\mem_bottom_track_17.DFFR_3_.Q ),
    .Y(_0340_));
 sky130_fd_sc_hd__inv_2 _0624_ (.A(\mem_bottom_track_17.DFFR_2_.Q ),
    .Y(_0339_));
 sky130_fd_sc_hd__inv_2 _0625_ (.A(\mem_bottom_track_17.DFFR_1_.Q ),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _0626_ (.A(\mem_bottom_track_17.DFFR_7_.Q ),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_2 _0627_ (.A(\mem_bottom_track_17.DFFR_6_.Q ),
    .Y(_0330_));
 sky130_fd_sc_hd__inv_2 _0628_ (.A(\mem_bottom_track_17.DFFR_0_.Q ),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _0629_ (.A(\mem_bottom_track_17.DFFR_3_.Q ),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _0630_ (.A(\mem_bottom_track_17.DFFR_2_.Q ),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _0631_ (.A(\mem_bottom_track_17.DFFR_1_.Q ),
    .Y(_0332_));
 sky130_fd_sc_hd__inv_2 _0632_ (.A(\mem_bottom_track_17.DFFR_5_.Q ),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _0633_ (.A(\mem_bottom_track_17.DFFR_0_.Q ),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_2 _0634_ (.A(\mem_bottom_track_17.DFFR_3_.Q ),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _0635_ (.A(\mem_bottom_track_17.DFFR_2_.Q ),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _0636_ (.A(\mem_bottom_track_17.DFFR_1_.Q ),
    .Y(_0335_));
 sky130_fd_sc_hd__inv_2 _0637_ (.A(\mem_bottom_track_9.DFFR_4_.Q ),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _0638_ (.A(\mem_bottom_track_9.DFFR_0_.Q ),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _0639_ (.A(\mem_bottom_track_9.DFFR_3_.Q ),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_2 _0640_ (.A(\mem_bottom_track_9.DFFR_2_.Q ),
    .Y(_0323_));
 sky130_fd_sc_hd__inv_2 _0641_ (.A(\mem_bottom_track_9.DFFR_1_.Q ),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _0642_ (.A(\mem_bottom_track_17.DFFR_0_.D ),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _0643_ (.A(\mem_bottom_track_9.DFFR_6_.Q ),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_2 _0644_ (.A(\mem_bottom_track_9.DFFR_0_.Q ),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _0645_ (.A(\mem_bottom_track_9.DFFR_3_.Q ),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _0646_ (.A(\mem_bottom_track_9.DFFR_2_.Q ),
    .Y(_0317_));
 sky130_fd_sc_hd__inv_2 _0647_ (.A(\mem_bottom_track_9.DFFR_1_.Q ),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_2 _0648_ (.A(\mem_bottom_track_9.DFFR_5_.Q ),
    .Y(_0313_));
 sky130_fd_sc_hd__inv_2 _0649_ (.A(\mem_bottom_track_9.DFFR_0_.Q ),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _0650_ (.A(\mem_bottom_track_9.DFFR_3_.Q ),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _0651_ (.A(\mem_bottom_track_9.DFFR_2_.Q ),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _0652_ (.A(\mem_bottom_track_9.DFFR_1_.Q ),
    .Y(_0319_));
 sky130_fd_sc_hd__inv_2 _0653_ (.A(\mem_bottom_track_1.DFFR_4_.Q ),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_2 _0654_ (.A(\mem_bottom_track_1.DFFR_0_.Q ),
    .Y(_0312_));
 sky130_fd_sc_hd__inv_2 _0655_ (.A(\mem_bottom_track_1.DFFR_3_.Q ),
    .Y(_0308_));
 sky130_fd_sc_hd__inv_2 _0656_ (.A(\mem_bottom_track_1.DFFR_2_.Q ),
    .Y(_0307_));
 sky130_fd_sc_hd__inv_2 _0657_ (.A(\mem_bottom_track_1.DFFR_1_.Q ),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _0658_ (.A(\mem_bottom_track_1.DFFR_7_.Q ),
    .Y(_0299_));
 sky130_fd_sc_hd__inv_2 _0659_ (.A(\mem_bottom_track_1.DFFR_6_.Q ),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_2 _0660_ (.A(\mem_bottom_track_1.DFFR_0_.Q ),
    .Y(_0310_));
 sky130_fd_sc_hd__inv_2 _0661_ (.A(\mem_bottom_track_1.DFFR_3_.Q ),
    .Y(_0302_));
 sky130_fd_sc_hd__inv_2 _0662_ (.A(\mem_bottom_track_1.DFFR_2_.Q ),
    .Y(_0301_));
 sky130_fd_sc_hd__inv_2 _0663_ (.A(\mem_bottom_track_1.DFFR_1_.Q ),
    .Y(_0300_));
 sky130_fd_sc_hd__inv_2 _0664_ (.A(\mem_bottom_track_1.DFFR_5_.Q ),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_2 _0665_ (.A(\mem_bottom_track_1.DFFR_0_.Q ),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _0666_ (.A(\mem_bottom_track_1.DFFR_3_.Q ),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_2 _0667_ (.A(\mem_bottom_track_1.DFFR_2_.Q ),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_2 _0668_ (.A(\mem_bottom_track_1.DFFR_1_.Q ),
    .Y(_0303_));
 sky130_fd_sc_hd__inv_2 _0669_ (.A(\mem_right_track_24.DFFR_4_.Q ),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _0670_ (.A(\mem_right_track_24.DFFR_0_.Q ),
    .Y(_0296_));
 sky130_fd_sc_hd__inv_2 _0671_ (.A(\mem_right_track_24.DFFR_3_.Q ),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_2 _0672_ (.A(\mem_right_track_24.DFFR_2_.Q ),
    .Y(_0291_));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(\mem_right_track_24.DFFR_1_.Q ),
    .Y(_0290_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(\mem_right_track_24.DFFR_7_.Q ),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _0675_ (.A(\mem_right_track_24.DFFR_6_.Q ),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _0676_ (.A(\mem_right_track_24.DFFR_0_.Q ),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(\mem_right_track_24.DFFR_3_.Q ),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_2 _0678_ (.A(\mem_right_track_24.DFFR_2_.Q ),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _0679_ (.A(\mem_right_track_24.DFFR_1_.Q ),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(\mem_right_track_24.DFFR_5_.Q ),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _0681_ (.A(\mem_right_track_24.DFFR_0_.Q ),
    .Y(_0295_));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(\mem_right_track_24.DFFR_3_.Q ),
    .Y(_0289_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(\mem_right_track_24.DFFR_2_.Q ),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(\mem_right_track_24.DFFR_1_.Q ),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_2 _0685_ (.A(\mem_right_track_16.DFFR_4_.Q ),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _0686_ (.A(\mem_right_track_16.DFFR_0_.Q ),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_2 _0687_ (.A(\mem_right_track_16.DFFR_3_.Q ),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _0688_ (.A(\mem_right_track_16.DFFR_2_.Q ),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_2 _0689_ (.A(\mem_right_track_16.DFFR_1_.Q ),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _0690_ (.A(\mem_right_track_16.DFFR_7_.Q ),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(\mem_right_track_16.DFFR_6_.Q ),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_2 _0692_ (.A(\mem_right_track_16.DFFR_0_.Q ),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _0693_ (.A(\mem_right_track_16.DFFR_3_.Q ),
    .Y(_0270_));
 sky130_fd_sc_hd__inv_2 _0694_ (.A(\mem_right_track_16.DFFR_2_.Q ),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _0695_ (.A(\mem_right_track_16.DFFR_1_.Q ),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _0696_ (.A(\mem_right_track_16.DFFR_5_.Q ),
    .Y(_0265_));
 sky130_fd_sc_hd__inv_2 _0697_ (.A(\mem_right_track_16.DFFR_0_.Q ),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_2 _0698_ (.A(\mem_right_track_16.DFFR_3_.Q ),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(\mem_right_track_16.DFFR_2_.Q ),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(\mem_right_track_16.DFFR_1_.Q ),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(\mem_right_track_8.DFFR_4_.Q ),
    .Y(_0261_));
 sky130_fd_sc_hd__inv_2 _0702_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .Y(_0264_));
 sky130_fd_sc_hd__inv_2 _0703_ (.A(\mem_right_track_8.DFFR_3_.Q ),
    .Y(_0260_));
 sky130_fd_sc_hd__inv_2 _0704_ (.A(\mem_right_track_8.DFFR_2_.Q ),
    .Y(_0259_));
 sky130_fd_sc_hd__inv_2 _0705_ (.A(\mem_right_track_8.DFFR_1_.Q ),
    .Y(_0258_));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(\mem_right_track_16.DFFR_0_.D ),
    .Y(_0251_));
 sky130_fd_sc_hd__inv_2 _0707_ (.A(\mem_right_track_8.DFFR_6_.Q ),
    .Y(_0250_));
 sky130_fd_sc_hd__inv_2 _0708_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_2 _0709_ (.A(\mem_right_track_8.DFFR_3_.Q ),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_2 _0710_ (.A(\mem_right_track_8.DFFR_2_.Q ),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(\mem_right_track_8.DFFR_1_.Q ),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _0712_ (.A(\mem_right_track_8.DFFR_5_.Q ),
    .Y(_0249_));
 sky130_fd_sc_hd__inv_2 _0713_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .Y(_0263_));
 sky130_fd_sc_hd__inv_2 _0714_ (.A(\mem_right_track_8.DFFR_3_.Q ),
    .Y(_0257_));
 sky130_fd_sc_hd__inv_2 _0715_ (.A(\mem_right_track_8.DFFR_2_.Q ),
    .Y(_0256_));
 sky130_fd_sc_hd__inv_2 _0716_ (.A(\mem_right_track_8.DFFR_1_.Q ),
    .Y(_0255_));
 sky130_fd_sc_hd__inv_2 _0717_ (.A(\mem_right_track_0.DFFR_4_.Q ),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _0718_ (.A(\mem_right_track_0.DFFR_0_.Q ),
    .Y(_0248_));
 sky130_fd_sc_hd__inv_2 _0719_ (.A(\mem_right_track_0.DFFR_3_.Q ),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _0720_ (.A(\mem_right_track_0.DFFR_2_.Q ),
    .Y(_0243_));
 sky130_fd_sc_hd__inv_2 _0721_ (.A(\mem_right_track_0.DFFR_1_.Q ),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _0722_ (.A(\mem_right_track_0.DFFR_7_.Q ),
    .Y(_0235_));
 sky130_fd_sc_hd__inv_2 _0723_ (.A(\mem_right_track_0.DFFR_6_.Q ),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _0724_ (.A(\mem_right_track_0.DFFR_0_.Q ),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _0725_ (.A(\mem_right_track_0.DFFR_3_.Q ),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(\mem_right_track_0.DFFR_2_.Q ),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _0727_ (.A(\mem_right_track_0.DFFR_1_.Q ),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(\mem_right_track_0.DFFR_5_.Q ),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(\mem_right_track_0.DFFR_0_.Q ),
    .Y(_0247_));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(\mem_right_track_0.DFFR_3_.Q ),
    .Y(_0241_));
 sky130_fd_sc_hd__inv_2 _0731_ (.A(\mem_right_track_0.DFFR_2_.Q ),
    .Y(_0240_));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(\mem_right_track_0.DFFR_1_.Q ),
    .Y(_0239_));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(\mem_top_track_24.DFFR_4_.Q ),
    .Y(_0229_));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(\mem_top_track_24.DFFR_0_.Q ),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(\mem_top_track_24.DFFR_3_.Q ),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _0736_ (.A(\mem_top_track_24.DFFR_2_.Q ),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _0737_ (.A(\mem_top_track_24.DFFR_1_.Q ),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_2 _0738_ (.A(\mem_top_track_24.DFFR_7_.Q ),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_2 _0739_ (.A(\mem_top_track_24.DFFR_6_.Q ),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_2 _0740_ (.A(\mem_top_track_24.DFFR_0_.Q ),
    .Y(_0230_));
 sky130_fd_sc_hd__inv_2 _0741_ (.A(\mem_top_track_24.DFFR_3_.Q ),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_2 _0742_ (.A(\mem_top_track_24.DFFR_2_.Q ),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(\mem_top_track_24.DFFR_1_.Q ),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(\mem_top_track_24.DFFR_5_.Q ),
    .Y(_0217_));
 sky130_fd_sc_hd__inv_2 _0745_ (.A(\mem_top_track_24.DFFR_0_.Q ),
    .Y(_0231_));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(\mem_top_track_24.DFFR_3_.Q ),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _0747_ (.A(\mem_top_track_24.DFFR_2_.Q ),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(\mem_top_track_24.DFFR_1_.Q ),
    .Y(_0223_));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(\mem_top_track_16.DFFR_4_.Q ),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _0750_ (.A(\mem_top_track_16.DFFR_0_.Q ),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(\mem_top_track_16.DFFR_3_.Q ),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(\mem_top_track_16.DFFR_2_.Q ),
    .Y(_0211_));
 sky130_fd_sc_hd__inv_2 _0753_ (.A(\mem_top_track_16.DFFR_1_.Q ),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(\mem_top_track_16.DFFR_7_.Q ),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_2 _0755_ (.A(\mem_top_track_16.DFFR_6_.Q ),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(\mem_top_track_16.DFFR_0_.Q ),
    .Y(_0214_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(\mem_top_track_16.DFFR_3_.Q ),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(\mem_top_track_16.DFFR_2_.Q ),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(\mem_top_track_16.DFFR_1_.Q ),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_2 _0760_ (.A(\mem_top_track_16.DFFR_5_.Q ),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(\mem_top_track_16.DFFR_0_.Q ),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_2 _0762_ (.A(\mem_top_track_16.DFFR_3_.Q ),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(\mem_top_track_16.DFFR_2_.Q ),
    .Y(_0208_));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(\mem_top_track_16.DFFR_1_.Q ),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(\mem_top_track_8.DFFR_4_.Q ),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(\mem_top_track_8.DFFR_0_.Q ),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(\mem_top_track_8.DFFR_3_.Q ),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(\mem_top_track_8.DFFR_2_.Q ),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _0769_ (.A(\mem_top_track_8.DFFR_1_.Q ),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(\mem_top_track_16.DFFR_0_.D ),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(\mem_top_track_8.DFFR_6_.Q ),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(\mem_top_track_8.DFFR_0_.Q ),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(\mem_top_track_8.DFFR_3_.Q ),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _0774_ (.A(\mem_top_track_8.DFFR_2_.Q ),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(\mem_top_track_8.DFFR_1_.Q ),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(\mem_top_track_8.DFFR_5_.Q ),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(\mem_top_track_8.DFFR_0_.Q ),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(\mem_top_track_8.DFFR_3_.Q ),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(\mem_top_track_8.DFFR_2_.Q ),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(\mem_top_track_8.DFFR_1_.Q ),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _0781_ (.A(\mem_top_track_0.DFFR_4_.Q ),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _0782_ (.A(\mem_top_track_0.DFFR_0_.Q ),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _0783_ (.A(\mem_top_track_0.DFFR_3_.Q ),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _0784_ (.A(\mem_top_track_0.DFFR_2_.Q ),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _0785_ (.A(\mem_top_track_0.DFFR_1_.Q ),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(\mem_top_track_0.DFFR_7_.Q ),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(\mem_top_track_0.DFFR_6_.Q ),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _0788_ (.A(\mem_top_track_0.DFFR_0_.Q ),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(\mem_top_track_0.DFFR_3_.Q ),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(\mem_top_track_0.DFFR_2_.Q ),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _0791_ (.A(\mem_top_track_0.DFFR_1_.Q ),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(\mem_top_track_0.DFFR_5_.Q ),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(\mem_top_track_0.DFFR_0_.Q ),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _0794_ (.A(\mem_top_track_0.DFFR_3_.Q ),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _0795_ (.A(\mem_top_track_0.DFFR_2_.Q ),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _0796_ (.A(\mem_top_track_0.DFFR_1_.Q ),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_top_track_0.out ));
 sky130_fd_sc_hd__inv_2 _0798_ (.A(net91),
    .Y(\mux_top_track_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkinv_2 _0799_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_top_track_8.out ));
 sky130_fd_sc_hd__inv_2 _0800_ (.A(net92),
    .Y(\mux_top_track_8.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_top_track_16.out ));
 sky130_fd_sc_hd__inv_2 _0802_ (.A(net93),
    .Y(\mux_top_track_16.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0803_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_top_track_24.out ));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(net94),
    .Y(\mux_top_track_24.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_right_track_0.out ));
 sky130_fd_sc_hd__inv_2 _0806_ (.A(net89),
    .Y(\mux_right_track_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkinv_2 _0807_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_right_track_8.out ));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(net90),
    .Y(\mux_right_track_8.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0809_ (.A(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_right_track_16.out ));
 sky130_fd_sc_hd__inv_2 _0810_ (.A(net87),
    .Y(\mux_right_track_16.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0811_ (.A(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_right_track_24.out ));
 sky130_fd_sc_hd__inv_2 _0812_ (.A(net88),
    .Y(\mux_right_track_24.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0813_ (.A(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_bottom_track_1.out ));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(net22),
    .Y(\mux_bottom_track_1.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _0815_ (.A(net21),
    .Y(\mux_bottom_track_1.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _0816_ (.A(net6),
    .Y(\mux_bottom_track_1.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0817_ (.A(net3),
    .Y(\mux_bottom_track_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0818_ (.A(net31),
    .Y(\mux_bottom_track_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0819_ (.A(net29),
    .Y(\mux_bottom_track_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0820_ (.A(net40),
    .Y(\mux_bottom_track_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0821_ (.A(net25),
    .Y(\mux_bottom_track_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0822_ (.A(net67),
    .Y(\mux_bottom_track_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0823_ (.A(net78),
    .Y(\mux_bottom_track_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0824_ (.A(net63),
    .Y(\mux_bottom_track_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0825_ (.A(net10),
    .Y(\mux_bottom_track_1.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _0826_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_bottom_track_9.out ));
 sky130_fd_sc_hd__inv_2 _0827_ (.A(net8),
    .Y(\mux_bottom_track_9.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _0828_ (.A(net23),
    .Y(\mux_bottom_track_9.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _0829_ (.A(net16),
    .Y(\mux_bottom_track_9.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(net4),
    .Y(\mux_bottom_track_9.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0831_ (.A(net30),
    .Y(\mux_bottom_track_9.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0832_ (.A(net27),
    .Y(\mux_bottom_track_9.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(net42),
    .Y(\mux_bottom_track_9.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0834_ (.A(net35),
    .Y(\mux_bottom_track_9.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0835_ (.A(net68),
    .Y(\mux_bottom_track_9.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(net80),
    .Y(\mux_bottom_track_9.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(net73),
    .Y(\mux_bottom_track_9.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0838_ (.A(net11),
    .Y(\mux_bottom_track_9.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _0839_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_bottom_track_17.out ));
 sky130_fd_sc_hd__inv_2 _0840_ (.A(net12),
    .Y(\mux_bottom_track_17.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(net24),
    .Y(\mux_bottom_track_17.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _0842_ (.A(net17),
    .Y(\mux_bottom_track_17.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0843_ (.A(net1),
    .Y(\mux_bottom_track_17.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0844_ (.A(net32),
    .Y(\mux_bottom_track_17.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0845_ (.A(net43),
    .Y(\mux_bottom_track_17.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0846_ (.A(net41),
    .Y(\mux_bottom_track_17.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0847_ (.A(net36),
    .Y(\mux_bottom_track_17.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0848_ (.A(net70),
    .Y(\mux_bottom_track_17.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0849_ (.A(net81),
    .Y(\mux_bottom_track_17.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0850_ (.A(net74),
    .Y(\mux_bottom_track_17.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0851_ (.A(net13),
    .Y(\mux_bottom_track_17.INVTX1_11_.out ));
 sky130_fd_sc_hd__clkinv_2 _0852_ (.A(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_bottom_track_25.out ));
 sky130_fd_sc_hd__inv_2 _0853_ (.A(net14),
    .Y(\mux_bottom_track_25.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _0854_ (.A(net7),
    .Y(\mux_bottom_track_25.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _0855_ (.A(net19),
    .Y(\mux_bottom_track_25.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0856_ (.A(net2),
    .Y(\mux_bottom_track_25.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0857_ (.A(net33),
    .Y(\mux_bottom_track_25.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0858_ (.A(net26),
    .Y(\mux_bottom_track_25.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0859_ (.A(net38),
    .Y(\mux_bottom_track_25.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0860_ (.A(net37),
    .Y(\mux_bottom_track_25.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0861_ (.A(net71),
    .Y(\mux_bottom_track_25.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0862_ (.A(net64),
    .Y(\mux_bottom_track_25.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0863_ (.A(net76),
    .Y(\mux_bottom_track_25.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0864_ (.A(net15),
    .Y(\mux_bottom_track_25.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _0865_ (.A(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_left_track_1.out ));
 sky130_fd_sc_hd__inv_2 _0866_ (.A(net53),
    .Y(\mux_left_track_1.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _0867_ (.A(net48),
    .Y(\mux_left_track_1.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _0868_ (.A(net59),
    .Y(\mux_left_track_1.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0869_ (.A(net44),
    .Y(\mux_left_track_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0870_ (.A(net75),
    .Y(\mux_left_track_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0871_ (.A(net84),
    .Y(\mux_left_track_1.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _0872_ (.A(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_left_track_9.out ));
 sky130_fd_sc_hd__inv_2 _0873_ (.A(net49),
    .Y(\mux_left_track_9.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _0874_ (.A(net61),
    .Y(\mux_left_track_9.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _0875_ (.A(net56),
    .Y(\mux_left_track_9.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0876_ (.A(net54),
    .Y(\mux_left_track_9.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0877_ (.A(net72),
    .Y(\mux_left_track_9.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0878_ (.A(net85),
    .Y(\mux_left_track_9.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _0879_ (.A(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_left_track_17.out ));
 sky130_fd_sc_hd__inv_2 _0880_ (.A(net51),
    .Y(\mux_left_track_17.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _0881_ (.A(net62),
    .Y(\mux_left_track_17.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _0882_ (.A(net60),
    .Y(\mux_left_track_17.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0883_ (.A(net55),
    .Y(\mux_left_track_17.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0884_ (.A(net69),
    .Y(\mux_left_track_17.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0885_ (.A(net82),
    .Y(\mux_left_track_17.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _0886_ (.A(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ),
    .Y(\mux_left_track_25.out ));
 sky130_fd_sc_hd__inv_2 _0887_ (.A(net52),
    .Y(\mux_left_track_25.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _0888_ (.A(net46),
    .Y(\mux_left_track_25.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _0889_ (.A(net45),
    .Y(\mux_left_track_25.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _0890_ (.A(net57),
    .Y(\mux_left_track_25.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0891_ (.A(net65),
    .Y(\mux_left_track_25.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0892_ (.A(net83),
    .Y(\mux_left_track_25.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _0893_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(\mux_top_track_32.out ));
 sky130_fd_sc_hd__inv_2 _0894_ (.A(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(\mux_right_track_32.out ));
 sky130_fd_sc_hd__inv_2 _0895_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(\mux_bottom_track_33.out ));
 sky130_fd_sc_hd__inv_2 _0896_ (.A(net20),
    .Y(\mux_bottom_track_33.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0897_ (.A(net18),
    .Y(\mux_bottom_track_33.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0898_ (.A(net34),
    .Y(\mux_bottom_track_33.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _0899_ (.A(net28),
    .Y(\mux_bottom_track_33.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _0900_ (.A(net39),
    .Y(\mux_bottom_track_33.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0901_ (.A(net66),
    .Y(\mux_bottom_track_33.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0902_ (.A(net77),
    .Y(\mux_bottom_track_33.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0903_ (.A(net9),
    .Y(\mux_bottom_track_33.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _0904_ (.A(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(\mux_left_track_33.out ));
 sky130_fd_sc_hd__inv_2 _0905_ (.A(net47),
    .Y(\mux_left_track_33.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _0906_ (.A(net58),
    .Y(\mux_left_track_33.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _0907_ (.A(net79),
    .Y(\mux_left_track_33.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0908_ (.A(net50),
    .Y(\mux_left_track_33.INVTX1_7_.out ));
 sky130_fd_sc_hd__buf_2 _0909_ (.A(net86),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_4 _0910_ (.A(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__buf_4 _0911_ (.A(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__inv_2 _0912_ (.A(_0154_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0913_ (.A(_0154_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0914_ (.A(_0154_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0915_ (.A(_0154_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0916_ (.A(_0154_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0917_ (.A(_0154_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0918_ (.A(_0154_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0919_ (.A(_0154_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0920_ (.A(_0154_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0921_ (.A(_0154_),
    .Y(_0009_));
 sky130_fd_sc_hd__buf_4 _0922_ (.A(_0153_),
    .X(_0155_));
 sky130_fd_sc_hd__inv_2 _0923_ (.A(_0155_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0924_ (.A(_0155_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0925_ (.A(_0155_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0926_ (.A(_0155_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0927_ (.A(_0155_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0928_ (.A(_0155_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _0929_ (.A(_0155_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _0930_ (.A(_0155_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _0931_ (.A(_0155_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _0932_ (.A(_0155_),
    .Y(_0019_));
 sky130_fd_sc_hd__buf_4 _0933_ (.A(_0153_),
    .X(_0156_));
 sky130_fd_sc_hd__inv_2 _0934_ (.A(_0156_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _0935_ (.A(_0156_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0936_ (.A(_0156_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _0937_ (.A(_0156_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _0938_ (.A(_0156_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0939_ (.A(_0156_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _0940_ (.A(_0156_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _0941_ (.A(_0156_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _0942_ (.A(_0156_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0943_ (.A(_0156_),
    .Y(_0029_));
 sky130_fd_sc_hd__buf_4 _0944_ (.A(_0153_),
    .X(_0157_));
 sky130_fd_sc_hd__inv_2 _0945_ (.A(_0157_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0946_ (.A(_0157_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _0947_ (.A(_0157_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _0948_ (.A(_0157_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _0949_ (.A(_0157_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _0950_ (.A(_0157_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _0951_ (.A(_0157_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _0952_ (.A(_0157_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _0953_ (.A(_0157_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _0954_ (.A(_0157_),
    .Y(_0039_));
 sky130_fd_sc_hd__buf_6 _0955_ (.A(_0153_),
    .X(_0158_));
 sky130_fd_sc_hd__inv_2 _0956_ (.A(_0158_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _0957_ (.A(_0158_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _0958_ (.A(_0158_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _0959_ (.A(_0158_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _0960_ (.A(_0158_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _0961_ (.A(_0158_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _0962_ (.A(_0158_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _0963_ (.A(_0158_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _0964_ (.A(_0158_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _0965_ (.A(_0158_),
    .Y(_0049_));
 sky130_fd_sc_hd__buf_4 _0966_ (.A(_0153_),
    .X(_0159_));
 sky130_fd_sc_hd__inv_2 _0967_ (.A(_0159_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _0968_ (.A(_0159_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _0969_ (.A(_0159_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(_0159_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _0971_ (.A(_0159_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _0972_ (.A(_0159_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _0973_ (.A(_0159_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _0974_ (.A(_0159_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _0975_ (.A(_0159_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _0976_ (.A(_0159_),
    .Y(_0059_));
 sky130_fd_sc_hd__buf_4 _0977_ (.A(_0153_),
    .X(_0160_));
 sky130_fd_sc_hd__inv_2 _0978_ (.A(_0160_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _0979_ (.A(_0160_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _0980_ (.A(_0160_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _0981_ (.A(_0160_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _0982_ (.A(_0160_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _0983_ (.A(_0160_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _0984_ (.A(_0160_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _0985_ (.A(_0160_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _0986_ (.A(_0160_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _0987_ (.A(_0160_),
    .Y(_0069_));
 sky130_fd_sc_hd__clkbuf_8 _0988_ (.A(_0153_),
    .X(_0161_));
 sky130_fd_sc_hd__inv_2 _0989_ (.A(_0161_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(_0161_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(_0161_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _0992_ (.A(_0161_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _0993_ (.A(_0161_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _0994_ (.A(_0161_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _0995_ (.A(_0161_),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _0996_ (.A(_0161_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _0997_ (.A(_0161_),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _0998_ (.A(_0161_),
    .Y(_0079_));
 sky130_fd_sc_hd__buf_4 _0999_ (.A(_0152_),
    .X(_0162_));
 sky130_fd_sc_hd__inv_2 _1000_ (.A(_0162_),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1001_ (.A(_0162_),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1002_ (.A(_0162_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1003_ (.A(_0162_),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _1004_ (.A(_0162_),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1005_ (.A(_0162_),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _1006_ (.A(_0162_),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1007_ (.A(_0162_),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(_0162_),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _1009_ (.A(_0162_),
    .Y(_0089_));
 sky130_fd_sc_hd__buf_4 _1010_ (.A(_0152_),
    .X(_0163_));
 sky130_fd_sc_hd__inv_2 _1011_ (.A(_0163_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1012_ (.A(_0163_),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _1013_ (.A(_0163_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1014_ (.A(_0163_),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _1015_ (.A(_0163_),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _1016_ (.A(_0163_),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _1017_ (.A(_0163_),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _1018_ (.A(_0163_),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _1019_ (.A(_0163_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1020_ (.A(_0163_),
    .Y(_0099_));
 sky130_fd_sc_hd__buf_4 _1021_ (.A(_0152_),
    .X(_0164_));
 sky130_fd_sc_hd__inv_2 _1022_ (.A(_0164_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1023_ (.A(_0164_),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _1024_ (.A(_0164_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _1025_ (.A(_0164_),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _1026_ (.A(_0164_),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1027_ (.A(_0164_),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(_0164_),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _1029_ (.A(_0164_),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _1030_ (.A(_0164_),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _1031_ (.A(_0164_),
    .Y(_0109_));
 sky130_fd_sc_hd__buf_4 _1032_ (.A(_0152_),
    .X(_0165_));
 sky130_fd_sc_hd__inv_2 _1033_ (.A(_0165_),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _1034_ (.A(_0165_),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _1035_ (.A(_0165_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(_0165_),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _1037_ (.A(_0165_),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1038_ (.A(_0165_),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _1039_ (.A(_0165_),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1040_ (.A(_0165_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1041_ (.A(_0165_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1042_ (.A(_0165_),
    .Y(_0119_));
 sky130_fd_sc_hd__buf_6 _1043_ (.A(_0152_),
    .X(_0166_));
 sky130_fd_sc_hd__inv_2 _1044_ (.A(_0166_),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1045_ (.A(_0166_),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _1046_ (.A(_0166_),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _1047_ (.A(_0166_),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _1048_ (.A(_0166_),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(_0166_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(_0166_),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(_0166_),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(_0166_),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(_0166_),
    .Y(_0129_));
 sky130_fd_sc_hd__buf_4 _1054_ (.A(_0152_),
    .X(_0167_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(_0167_),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(_0167_),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _1057_ (.A(_0167_),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(_0167_),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(_0167_),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _1060_ (.A(_0167_),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _1061_ (.A(_0167_),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(_0167_),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(_0167_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1064_ (.A(_0167_),
    .Y(_0139_));
 sky130_fd_sc_hd__buf_4 _1065_ (.A(_0152_),
    .X(_0168_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(_0168_),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(_0168_),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(_0168_),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(_0168_),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(_0168_),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _1071_ (.A(_0168_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _1072_ (.A(_0168_),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(_0168_),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _1074_ (.A(_0168_),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1075_ (.A(_0168_),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(_0153_),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(_0153_),
    .Y(_0151_));
 sky130_fd_sc_hd__dfrtp_1 _1078_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_top_track_0.DFFR_6_.Q ),
    .RESET_B(_0000_),
    .Q(\mem_top_track_0.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1079_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_top_track_0.DFFR_5_.Q ),
    .RESET_B(_0001_),
    .Q(\mem_top_track_0.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1080_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_top_track_0.DFFR_4_.Q ),
    .RESET_B(_0002_),
    .Q(\mem_top_track_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1081_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_top_track_0.DFFR_3_.Q ),
    .RESET_B(_0003_),
    .Q(\mem_top_track_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1082_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_top_track_0.DFFR_2_.Q ),
    .RESET_B(_0004_),
    .Q(\mem_top_track_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1083_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_top_track_0.DFFR_1_.Q ),
    .RESET_B(_0005_),
    .Q(\mem_top_track_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1084_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_top_track_0.DFFR_0_.Q ),
    .RESET_B(_0006_),
    .Q(\mem_top_track_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1085_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net5),
    .RESET_B(_0007_),
    .Q(\mem_top_track_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1086_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_top_track_8.DFFR_6_.Q ),
    .RESET_B(_0008_),
    .Q(\mem_top_track_16.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_1 _1087_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_top_track_8.DFFR_5_.Q ),
    .RESET_B(_0009_),
    .Q(\mem_top_track_8.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1088_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_top_track_8.DFFR_4_.Q ),
    .RESET_B(_0010_),
    .Q(\mem_top_track_8.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1089_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_top_track_8.DFFR_3_.Q ),
    .RESET_B(_0011_),
    .Q(\mem_top_track_8.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1090_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_top_track_8.DFFR_2_.Q ),
    .RESET_B(_0012_),
    .Q(\mem_top_track_8.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _1091_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_top_track_8.DFFR_1_.Q ),
    .RESET_B(_0013_),
    .Q(\mem_top_track_8.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1092_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_top_track_8.DFFR_0_.Q ),
    .RESET_B(_0014_),
    .Q(\mem_top_track_8.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1093_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_top_track_0.DFFR_7_.Q ),
    .RESET_B(_0015_),
    .Q(\mem_top_track_8.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1094_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_top_track_16.DFFR_6_.Q ),
    .RESET_B(_0016_),
    .Q(\mem_top_track_16.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1095_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_top_track_16.DFFR_5_.Q ),
    .RESET_B(_0017_),
    .Q(\mem_top_track_16.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1096_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_top_track_16.DFFR_4_.Q ),
    .RESET_B(_0018_),
    .Q(\mem_top_track_16.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1097_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_top_track_16.DFFR_3_.Q ),
    .RESET_B(_0019_),
    .Q(\mem_top_track_16.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1098_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_top_track_16.DFFR_2_.Q ),
    .RESET_B(_0020_),
    .Q(\mem_top_track_16.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1099_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_top_track_16.DFFR_1_.Q ),
    .RESET_B(_0021_),
    .Q(\mem_top_track_16.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1100_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_top_track_16.DFFR_0_.Q ),
    .RESET_B(_0022_),
    .Q(\mem_top_track_16.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1101_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_top_track_16.DFFR_0_.D ),
    .RESET_B(_0023_),
    .Q(\mem_top_track_16.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_top_track_24.DFFR_6_.Q ),
    .RESET_B(_0024_),
    .Q(\mem_top_track_24.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1103_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_top_track_24.DFFR_5_.Q ),
    .RESET_B(_0025_),
    .Q(\mem_top_track_24.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1104_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_top_track_24.DFFR_4_.Q ),
    .RESET_B(_0026_),
    .Q(\mem_top_track_24.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1105_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_top_track_24.DFFR_3_.Q ),
    .RESET_B(_0027_),
    .Q(\mem_top_track_24.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1106_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_top_track_24.DFFR_2_.Q ),
    .RESET_B(_0028_),
    .Q(\mem_top_track_24.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1107_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_top_track_24.DFFR_1_.Q ),
    .RESET_B(_0029_),
    .Q(\mem_top_track_24.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1108_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_top_track_24.DFFR_0_.Q ),
    .RESET_B(_0030_),
    .Q(\mem_top_track_24.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1109_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_top_track_16.DFFR_7_.Q ),
    .RESET_B(_0031_),
    .Q(\mem_top_track_24.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1110_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_right_track_0.DFFR_6_.Q ),
    .RESET_B(_0032_),
    .Q(\mem_right_track_0.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1111_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_right_track_0.DFFR_5_.Q ),
    .RESET_B(_0033_),
    .Q(\mem_right_track_0.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1112_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_right_track_0.DFFR_4_.Q ),
    .RESET_B(_0034_),
    .Q(\mem_right_track_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1113_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_0.DFFR_3_.Q ),
    .RESET_B(_0035_),
    .Q(\mem_right_track_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1114_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_0.DFFR_2_.Q ),
    .RESET_B(_0036_),
    .Q(\mem_right_track_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1115_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_right_track_0.DFFR_1_.Q ),
    .RESET_B(_0037_),
    .Q(\mem_right_track_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1116_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_right_track_0.DFFR_0_.Q ),
    .RESET_B(_0038_),
    .Q(\mem_right_track_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1117_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_right_track_0.DFFR_0_.D ),
    .RESET_B(_0039_),
    .Q(\mem_right_track_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1118_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_right_track_8.DFFR_6_.Q ),
    .RESET_B(_0040_),
    .Q(\mem_right_track_16.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_1 _1119_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_right_track_8.DFFR_5_.Q ),
    .RESET_B(_0041_),
    .Q(\mem_right_track_8.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_right_track_8.DFFR_4_.Q ),
    .RESET_B(_0042_),
    .Q(\mem_right_track_8.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1121_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_right_track_8.DFFR_3_.Q ),
    .RESET_B(_0043_),
    .Q(\mem_right_track_8.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1122_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_right_track_8.DFFR_2_.Q ),
    .RESET_B(_0044_),
    .Q(\mem_right_track_8.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1123_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_right_track_8.DFFR_1_.Q ),
    .RESET_B(_0045_),
    .Q(\mem_right_track_8.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1124_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_8.DFFR_0_.Q ),
    .RESET_B(_0046_),
    .Q(\mem_right_track_8.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1125_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_right_track_0.DFFR_7_.Q ),
    .RESET_B(_0047_),
    .Q(\mem_right_track_8.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1126_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_right_track_16.DFFR_6_.Q ),
    .RESET_B(_0048_),
    .Q(\mem_right_track_16.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1127_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_right_track_16.DFFR_5_.Q ),
    .RESET_B(_0049_),
    .Q(\mem_right_track_16.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_right_track_16.DFFR_4_.Q ),
    .RESET_B(_0050_),
    .Q(\mem_right_track_16.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1129_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_right_track_16.DFFR_3_.Q ),
    .RESET_B(_0051_),
    .Q(\mem_right_track_16.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1130_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_right_track_16.DFFR_2_.Q ),
    .RESET_B(_0052_),
    .Q(\mem_right_track_16.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1131_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_right_track_16.DFFR_1_.Q ),
    .RESET_B(_0053_),
    .Q(\mem_right_track_16.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1132_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_right_track_16.DFFR_0_.Q ),
    .RESET_B(_0054_),
    .Q(\mem_right_track_16.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1133_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_right_track_16.DFFR_0_.D ),
    .RESET_B(_0055_),
    .Q(\mem_right_track_16.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_right_track_24.DFFR_6_.Q ),
    .RESET_B(_0056_),
    .Q(\mem_right_track_24.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1135_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_right_track_24.DFFR_5_.Q ),
    .RESET_B(_0057_),
    .Q(\mem_right_track_24.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1136_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_24.DFFR_4_.Q ),
    .RESET_B(_0058_),
    .Q(\mem_right_track_24.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1137_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_24.DFFR_3_.Q ),
    .RESET_B(_0059_),
    .Q(\mem_right_track_24.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1138_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_right_track_24.DFFR_2_.Q ),
    .RESET_B(_0060_),
    .Q(\mem_right_track_24.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1139_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_right_track_24.DFFR_1_.Q ),
    .RESET_B(_0061_),
    .Q(\mem_right_track_24.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1140_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_right_track_24.DFFR_0_.Q ),
    .RESET_B(_0062_),
    .Q(\mem_right_track_24.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1141_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_right_track_16.DFFR_7_.Q ),
    .RESET_B(_0063_),
    .Q(\mem_right_track_24.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1142_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_6_.Q ),
    .RESET_B(_0064_),
    .Q(\mem_bottom_track_1.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1143_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_5_.Q ),
    .RESET_B(_0065_),
    .Q(\mem_bottom_track_1.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1144_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_4_.Q ),
    .RESET_B(_0066_),
    .Q(\mem_bottom_track_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1145_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_3_.Q ),
    .RESET_B(_0067_),
    .Q(\mem_bottom_track_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1146_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_2_.Q ),
    .RESET_B(_0068_),
    .Q(\mem_bottom_track_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1147_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_1_.Q ),
    .RESET_B(_0069_),
    .Q(\mem_bottom_track_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1148_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_0_.Q ),
    .RESET_B(_0070_),
    .Q(\mem_bottom_track_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1149_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_0_.D ),
    .RESET_B(_0071_),
    .Q(\mem_bottom_track_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1150_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_6_.Q ),
    .RESET_B(_0072_),
    .Q(\mem_bottom_track_17.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_1 _1151_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_5_.Q ),
    .RESET_B(_0073_),
    .Q(\mem_bottom_track_9.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1152_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_4_.Q ),
    .RESET_B(_0074_),
    .Q(\mem_bottom_track_9.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1153_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_3_.Q ),
    .RESET_B(_0075_),
    .Q(\mem_bottom_track_9.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1154_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_2_.Q ),
    .RESET_B(_0076_),
    .Q(\mem_bottom_track_9.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1155_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_1_.Q ),
    .RESET_B(_0077_),
    .Q(\mem_bottom_track_9.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1156_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_bottom_track_9.DFFR_0_.Q ),
    .RESET_B(_0078_),
    .Q(\mem_bottom_track_9.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1157_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_bottom_track_1.DFFR_7_.Q ),
    .RESET_B(_0079_),
    .Q(\mem_bottom_track_9.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1158_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_6_.Q ),
    .RESET_B(_0080_),
    .Q(\mem_bottom_track_17.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1159_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_5_.Q ),
    .RESET_B(_0081_),
    .Q(\mem_bottom_track_17.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1160_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_4_.Q ),
    .RESET_B(_0082_),
    .Q(\mem_bottom_track_17.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1161_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_3_.Q ),
    .RESET_B(_0083_),
    .Q(\mem_bottom_track_17.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1162_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_2_.Q ),
    .RESET_B(_0084_),
    .Q(\mem_bottom_track_17.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1163_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_1_.Q ),
    .RESET_B(_0085_),
    .Q(\mem_bottom_track_17.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1164_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_0_.Q ),
    .RESET_B(_0086_),
    .Q(\mem_bottom_track_17.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1165_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_0_.D ),
    .RESET_B(_0087_),
    .Q(\mem_bottom_track_17.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1166_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_6_.Q ),
    .RESET_B(_0088_),
    .Q(\mem_bottom_track_25.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1167_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_5_.Q ),
    .RESET_B(_0089_),
    .Q(\mem_bottom_track_25.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1168_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_4_.Q ),
    .RESET_B(_0090_),
    .Q(\mem_bottom_track_25.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1169_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_3_.Q ),
    .RESET_B(_0091_),
    .Q(\mem_bottom_track_25.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1170_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_2_.Q ),
    .RESET_B(_0092_),
    .Q(\mem_bottom_track_25.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1171_ (.CLK(clknet_4_13_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_1_.Q ),
    .RESET_B(_0093_),
    .Q(\mem_bottom_track_25.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1172_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_0_.Q ),
    .RESET_B(_0094_),
    .Q(\mem_bottom_track_25.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1173_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_bottom_track_17.DFFR_7_.Q ),
    .RESET_B(_0095_),
    .Q(\mem_bottom_track_25.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1174_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_left_track_1.DFFR_6_.Q ),
    .RESET_B(_0096_),
    .Q(\mem_left_track_1.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1175_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_left_track_1.DFFR_5_.Q ),
    .RESET_B(_0097_),
    .Q(\mem_left_track_1.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1176_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_left_track_1.DFFR_4_.Q ),
    .RESET_B(_0098_),
    .Q(\mem_left_track_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1177_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_left_track_1.DFFR_3_.Q ),
    .RESET_B(_0099_),
    .Q(\mem_left_track_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1178_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_left_track_1.DFFR_2_.Q ),
    .RESET_B(_0100_),
    .Q(\mem_left_track_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1179_ (.CLK(clknet_4_6_0_prog_clk),
    .D(\mem_left_track_1.DFFR_1_.Q ),
    .RESET_B(_0101_),
    .Q(\mem_left_track_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1180_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_left_track_1.DFFR_0_.Q ),
    .RESET_B(_0102_),
    .Q(\mem_left_track_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1181_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_5_.Q ),
    .RESET_B(_0103_),
    .Q(\mem_left_track_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1182_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_left_track_9.DFFR_6_.Q ),
    .RESET_B(_0104_),
    .Q(\mem_left_track_17.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_1 _1183_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_left_track_9.DFFR_5_.Q ),
    .RESET_B(_0105_),
    .Q(\mem_left_track_9.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1184_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_left_track_9.DFFR_4_.Q ),
    .RESET_B(_0106_),
    .Q(\mem_left_track_9.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1185_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_left_track_9.DFFR_3_.Q ),
    .RESET_B(_0107_),
    .Q(\mem_left_track_9.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _1186_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_left_track_9.DFFR_2_.Q ),
    .RESET_B(_0108_),
    .Q(\mem_left_track_9.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1187_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_left_track_9.DFFR_1_.Q ),
    .RESET_B(_0109_),
    .Q(\mem_left_track_9.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _1188_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_left_track_9.DFFR_0_.Q ),
    .RESET_B(_0110_),
    .Q(\mem_left_track_9.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1189_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_left_track_1.DFFR_7_.Q ),
    .RESET_B(_0111_),
    .Q(\mem_left_track_9.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1190_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_left_track_17.DFFR_6_.Q ),
    .RESET_B(_0112_),
    .Q(\mem_left_track_17.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1191_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_left_track_17.DFFR_5_.Q ),
    .RESET_B(_0113_),
    .Q(\mem_left_track_17.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1192_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_left_track_17.DFFR_4_.Q ),
    .RESET_B(_0114_),
    .Q(\mem_left_track_17.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1193_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_left_track_17.DFFR_3_.Q ),
    .RESET_B(_0115_),
    .Q(\mem_left_track_17.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1194_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_left_track_17.DFFR_2_.Q ),
    .RESET_B(_0116_),
    .Q(\mem_left_track_17.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1195_ (.CLK(clknet_4_15_0_prog_clk),
    .D(\mem_left_track_17.DFFR_1_.Q ),
    .RESET_B(_0117_),
    .Q(\mem_left_track_17.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1196_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_left_track_17.DFFR_0_.Q ),
    .RESET_B(_0118_),
    .Q(\mem_left_track_17.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1197_ (.CLK(clknet_4_14_0_prog_clk),
    .D(\mem_left_track_17.DFFR_0_.D ),
    .RESET_B(_0119_),
    .Q(\mem_left_track_17.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1198_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_left_track_25.DFFR_6_.Q ),
    .RESET_B(_0120_),
    .Q(\mem_left_track_25.DFFR_7_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1199_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_left_track_25.DFFR_5_.Q ),
    .RESET_B(_0121_),
    .Q(\mem_left_track_25.DFFR_6_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1200_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_left_track_25.DFFR_4_.Q ),
    .RESET_B(_0122_),
    .Q(\mem_left_track_25.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1201_ (.CLK(clknet_4_0_0_prog_clk),
    .D(\mem_left_track_25.DFFR_3_.Q ),
    .RESET_B(_0123_),
    .Q(\mem_left_track_25.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1202_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_left_track_25.DFFR_2_.Q ),
    .RESET_B(_0124_),
    .Q(\mem_left_track_25.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1203_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_left_track_25.DFFR_1_.Q ),
    .RESET_B(_0125_),
    .Q(\mem_left_track_25.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1204_ (.CLK(clknet_4_8_0_prog_clk),
    .D(\mem_left_track_25.DFFR_0_.Q ),
    .RESET_B(_0126_),
    .Q(\mem_left_track_25.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1205_ (.CLK(clknet_4_11_0_prog_clk),
    .D(\mem_left_track_17.DFFR_7_.Q ),
    .RESET_B(_0127_),
    .Q(\mem_left_track_25.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1206_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_top_track_32.DFFR_4_.Q ),
    .RESET_B(_0128_),
    .Q(\mem_right_track_0.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_1 _1207_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_top_track_32.DFFR_3_.Q ),
    .RESET_B(_0129_),
    .Q(\mem_top_track_32.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1208_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_top_track_32.DFFR_2_.Q ),
    .RESET_B(_0130_),
    .Q(\mem_top_track_32.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1209_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_top_track_32.DFFR_1_.Q ),
    .RESET_B(_0131_),
    .Q(\mem_top_track_32.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1210_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_top_track_32.DFFR_0_.Q ),
    .RESET_B(_0132_),
    .Q(\mem_top_track_32.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1211_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_top_track_24.DFFR_7_.Q ),
    .RESET_B(_0133_),
    .Q(\mem_top_track_32.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1212_ (.CLK(clknet_4_12_0_prog_clk),
    .D(\mem_right_track_32.DFFR_4_.Q ),
    .RESET_B(_0134_),
    .Q(\mem_bottom_track_1.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_1 _1213_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_right_track_32.DFFR_3_.Q ),
    .RESET_B(_0135_),
    .Q(\mem_right_track_32.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1214_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_right_track_32.DFFR_2_.Q ),
    .RESET_B(_0136_),
    .Q(\mem_right_track_32.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1215_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_right_track_32.DFFR_1_.Q ),
    .RESET_B(_0137_),
    .Q(\mem_right_track_32.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1216_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_32.DFFR_0_.Q ),
    .RESET_B(_0138_),
    .Q(\mem_right_track_32.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1217_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_right_track_24.DFFR_7_.Q ),
    .RESET_B(_0139_),
    .Q(\mem_right_track_32.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1218_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_4_.Q ),
    .RESET_B(_0140_),
    .Q(\mem_bottom_track_33.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1219_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_3_.Q ),
    .RESET_B(_0141_),
    .Q(\mem_bottom_track_33.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1220_ (.CLK(clknet_4_10_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_2_.Q ),
    .RESET_B(_0142_),
    .Q(\mem_bottom_track_33.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1221_ (.CLK(clknet_4_9_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_1_.Q ),
    .RESET_B(_0143_),
    .Q(\mem_bottom_track_33.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1222_ (.CLK(clknet_4_2_0_prog_clk),
    .D(\mem_bottom_track_33.DFFR_0_.Q ),
    .RESET_B(_0144_),
    .Q(\mem_bottom_track_33.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1223_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_bottom_track_25.DFFR_7_.Q ),
    .RESET_B(_0145_),
    .Q(\mem_bottom_track_33.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _1224_ (.CLK(clknet_4_7_0_prog_clk),
    .D(\mem_left_track_33.DFFR_4_.Q ),
    .RESET_B(_0146_),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _1225_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_left_track_33.DFFR_3_.Q ),
    .RESET_B(_0147_),
    .Q(\mem_left_track_33.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _1226_ (.CLK(clknet_4_5_0_prog_clk),
    .D(\mem_left_track_33.DFFR_2_.Q ),
    .RESET_B(_0148_),
    .Q(\mem_left_track_33.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1227_ (.CLK(clknet_4_4_0_prog_clk),
    .D(\mem_left_track_33.DFFR_1_.Q ),
    .RESET_B(_0149_),
    .Q(\mem_left_track_33.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1228_ (.CLK(clknet_4_3_0_prog_clk),
    .D(\mem_left_track_33.DFFR_0_.Q ),
    .RESET_B(_0150_),
    .Q(\mem_left_track_33.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _1229_ (.CLK(clknet_4_1_0_prog_clk),
    .D(\mem_left_track_25.DFFR_7_.Q ),
    .RESET_B(_0151_),
    .Q(\mem_left_track_33.DFFR_0_.Q ));
 sky130_fd_sc_hd__conb_1 _1344__173 (.HI(net173));
 sky130_fd_sc_hd__conb_1 _1360__174 (.HI(net174));
 sky130_fd_sc_hd__conb_1 _1376__175 (.HI(net175));
 sky130_fd_sc_hd__conb_1 _1392__176 (.HI(net176));
 sky130_fd_sc_hd__conb_1 _1408__177 (.HI(net177));
 sky130_fd_sc_hd__conb_1 _1424__178 (.HI(net178));
 sky130_fd_sc_hd__conb_1 _1440__179 (.HI(net179));
 sky130_fd_sc_hd__conb_1 _1456__180 (.HI(net180));
 sky130_fd_sc_hd__conb_1 _1472__181 (.HI(net181));
 sky130_fd_sc_hd__conb_1 _1488__182 (.HI(net182));
 sky130_fd_sc_hd__conb_1 _1504__183 (.HI(net183));
 sky130_fd_sc_hd__conb_1 _1520__184 (.HI(net184));
 sky130_fd_sc_hd__conb_1 _1536__185 (.HI(net185));
 sky130_fd_sc_hd__conb_1 _1552__186 (.HI(net186));
 sky130_fd_sc_hd__conb_1 _1568__187 (.HI(net187));
 sky130_fd_sc_hd__conb_1 _1585__188 (.HI(net188));
 sky130_fd_sc_hd__conb_1 _1597__189 (.HI(net189));
 sky130_fd_sc_hd__conb_1 _1609__190 (.HI(net190));
 sky130_fd_sc_hd__conb_1 _1621__191 (.HI(net191));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_prog_clk (.A(prog_clk),
    .X(clknet_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_2 _1250_ (.A(net33),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 _1251_ (.A(net32),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 _1252_ (.A(\mux_left_track_33.out ),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _1253_ (.A(net30),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _1254_ (.A(net29),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 _1255_ (.A(net28),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _1256_ (.A(\mux_left_track_25.out ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _1257_ (.A(net26),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _1258_ (.A(net43),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _1259_ (.A(net42),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 _1260_ (.A(\mux_left_track_17.out ),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 _1261_ (.A(net40),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 _1262_ (.A(net39),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 _1263_ (.A(net38),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 _1264_ (.A(\mux_left_track_9.out ),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 _1265_ (.A(net36),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 _1266_ (.A(net35),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 _1267_ (.A(net25),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 _1268_ (.A(\mux_left_track_1.out ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _1269_ (.A(net14),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _1270_ (.A(net13),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 _1271_ (.A(\mux_right_track_32.out ),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 _1272_ (.A(net11),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 _1273_ (.A(net10),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 _1274_ (.A(net9),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 _1275_ (.A(\mux_right_track_24.out ),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 _1276_ (.A(net7),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 _1277_ (.A(net24),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 _1278_ (.A(net23),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 _1279_ (.A(\mux_right_track_16.out ),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 _1280_ (.A(net21),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 _1281_ (.A(net20),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 _1282_ (.A(net19),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _1283_ (.A(\mux_right_track_8.out ),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 _1284_ (.A(net17),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 _1285_ (.A(net16),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 _1286_ (.A(net6),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 _1287_ (.A(\mux_right_track_0.out ),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 _1288_ (.A(net71),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 _1289_ (.A(net70),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _1290_ (.A(\mux_bottom_track_33.out ),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _1291_ (.A(net68),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 _1292_ (.A(net67),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 _1293_ (.A(net66),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 _1294_ (.A(\mux_bottom_track_25.out ),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 _1295_ (.A(net64),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 _1296_ (.A(net81),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 _1297_ (.A(net80),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _1298_ (.A(\mux_bottom_track_17.out ),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _1299_ (.A(net78),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _1300_ (.A(net77),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _1301_ (.A(net76),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _1302_ (.A(\mux_bottom_track_9.out ),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 _1303_ (.A(net74),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 _1304_ (.A(net73),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 _1305_ (.A(net63),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 _1306_ (.A(\mux_bottom_track_1.out ),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 _1307_ (.A(net52),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 _1308_ (.A(net51),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _1309_ (.A(\mux_top_track_32.out ),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _1310_ (.A(net49),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _1311_ (.A(net48),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 _1312_ (.A(net47),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 _1313_ (.A(\mux_top_track_24.out ),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 _1314_ (.A(net45),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 _1315_ (.A(net62),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _1316_ (.A(net61),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 _1317_ (.A(\mux_top_track_16.out ),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 _1318_ (.A(net59),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 _1319_ (.A(net58),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 _1320_ (.A(net57),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 _1321_ (.A(\mux_top_track_8.out ),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 _1322_ (.A(net55),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 _1323_ (.A(net54),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 _1324_ (.A(net44),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 _1325_ (.A(\mux_top_track_0.out ),
    .X(net153));
 sky130_fd_sc_hd__ebufn_4 _1326_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0169_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1327_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0170_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1328_ (.A(net172),
    .TE_B(_0171_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1329_ (.A(\mux_bottom_track_33.INVTX1_5_.out ),
    .TE_B(_0172_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1330_ (.A(\mux_bottom_track_1.INVTX1_9_.out ),
    .TE_B(_0173_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1331_ (.A(\mux_bottom_track_1.INVTX1_11_.out ),
    .TE_B(_0174_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1332_ (.A(\mux_left_track_1.INVTX1_7_.out ),
    .TE_B(_0175_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1333_ (.A(\mux_left_track_1.INVTX1_8_.out ),
    .TE_B(_0176_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1334_ (.A(\mux_left_track_1.INVTX1_9_.out ),
    .TE_B(_0177_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1335_ (.A(\mux_bottom_track_1.INVTX1_3_.out ),
    .TE_B(_0178_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1336_ (.A(\mux_bottom_track_1.INVTX1_4_.out ),
    .TE_B(_0179_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1337_ (.A(\mux_bottom_track_17.INVTX1_4_.out ),
    .TE_B(_0180_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1338_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0181_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1339_ (.A(\mux_bottom_track_1.INVTX1_8_.out ),
    .TE_B(_0182_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1340_ (.A(\mux_bottom_track_1.INVTX1_5_.out ),
    .TE_B(_0183_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1341_ (.A(\mux_top_track_0.INVTX1_0_.out ),
    .TE_B(_0184_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1342_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0185_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1343_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0186_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1344_ (.A(net173),
    .TE_B(_0187_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1345_ (.A(\mux_bottom_track_9.INVTX1_9_.out ),
    .TE_B(_0188_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1346_ (.A(\mux_bottom_track_9.INVTX1_11_.out ),
    .TE_B(_0189_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1347_ (.A(\mux_bottom_track_25.INVTX1_11_.out ),
    .TE_B(_0190_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1348_ (.A(\mux_left_track_9.INVTX1_7_.out ),
    .TE_B(_0191_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1349_ (.A(\mux_left_track_9.INVTX1_9_.out ),
    .TE_B(_0192_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1350_ (.A(\mux_left_track_9.INVTX1_10_.out ),
    .TE_B(_0193_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1351_ (.A(\mux_bottom_track_9.INVTX1_3_.out ),
    .TE_B(_0194_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1352_ (.A(\mux_bottom_track_9.INVTX1_4_.out ),
    .TE_B(_0195_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1353_ (.A(\mux_bottom_track_9.INVTX1_5_.out ),
    .TE_B(_0196_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1354_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0197_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1355_ (.A(\mux_bottom_track_9.INVTX1_8_.out ),
    .TE_B(_0198_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1356_ (.A(\mux_bottom_track_9.INVTX1_6_.out ),
    .TE_B(_0199_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1357_ (.A(\mux_top_track_8.INVTX1_0_.out ),
    .TE_B(_0200_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1358_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0201_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1359_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0202_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1360_ (.A(net174),
    .TE_B(_0203_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1361_ (.A(\mux_bottom_track_17.INVTX1_9_.out ),
    .TE_B(_0204_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1362_ (.A(\mux_bottom_track_17.INVTX1_10_.out ),
    .TE_B(_0205_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1363_ (.A(\mux_bottom_track_17.INVTX1_11_.out ),
    .TE_B(_0206_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1364_ (.A(\mux_left_track_17.INVTX1_7_.out ),
    .TE_B(_0207_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1365_ (.A(\mux_left_track_17.INVTX1_9_.out ),
    .TE_B(_0208_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1366_ (.A(\mux_left_track_17.INVTX1_10_.out ),
    .TE_B(_0209_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1367_ (.A(\mux_bottom_track_17.INVTX1_3_.out ),
    .TE_B(_0210_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1368_ (.A(\mux_bottom_track_17.INVTX1_5_.out ),
    .TE_B(_0211_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1369_ (.A(\mux_bottom_track_1.INVTX1_6_.out ),
    .TE_B(_0212_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1370_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0213_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1371_ (.A(\mux_bottom_track_17.INVTX1_8_.out ),
    .TE_B(_0214_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1372_ (.A(\mux_bottom_track_17.INVTX1_6_.out ),
    .TE_B(_0215_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1373_ (.A(\mux_top_track_16.INVTX1_0_.out ),
    .TE_B(_0216_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1374_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0217_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1375_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0218_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1376_ (.A(net175),
    .TE_B(_0219_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1377_ (.A(\mux_bottom_track_25.INVTX1_9_.out ),
    .TE_B(_0220_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1378_ (.A(\mux_bottom_track_9.INVTX1_10_.out ),
    .TE_B(_0221_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1379_ (.A(\mux_bottom_track_25.INVTX1_10_.out ),
    .TE_B(_0222_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1380_ (.A(\mux_left_track_25.INVTX1_7_.out ),
    .TE_B(_0223_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1381_ (.A(\mux_left_track_25.INVTX1_8_.out ),
    .TE_B(_0224_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1382_ (.A(\mux_left_track_25.INVTX1_10_.out ),
    .TE_B(_0225_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1383_ (.A(\mux_bottom_track_25.INVTX1_4_.out ),
    .TE_B(_0226_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1384_ (.A(\mux_bottom_track_25.INVTX1_5_.out ),
    .TE_B(_0227_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1385_ (.A(\mux_bottom_track_25.INVTX1_6_.out ),
    .TE_B(_0228_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1386_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0229_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1387_ (.A(\mux_bottom_track_25.INVTX1_8_.out ),
    .TE_B(_0230_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1388_ (.A(\mux_bottom_track_33.INVTX1_4_.out ),
    .TE_B(_0231_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1389_ (.A(\mux_top_track_24.INVTX1_0_.out ),
    .TE_B(_0232_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1390_ (.A(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0233_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1391_ (.A(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0234_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1392_ (.A(net176),
    .TE_B(_0235_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1393_ (.A(\mux_bottom_track_1.INVTX1_8_.out ),
    .TE_B(_0236_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1394_ (.A(\mux_bottom_track_1.INVTX1_9_.out ),
    .TE_B(_0237_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1395_ (.A(\mux_bottom_track_1.INVTX1_11_.out ),
    .TE_B(_0238_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1396_ (.A(\mux_left_track_1.INVTX1_7_.out ),
    .TE_B(_0239_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1397_ (.A(\mux_left_track_1.INVTX1_8_.out ),
    .TE_B(_0240_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1398_ (.A(\mux_left_track_1.INVTX1_9_.out ),
    .TE_B(_0241_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_8 _1399_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_0242_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_8 _1400_ (.A(\mux_bottom_track_1.INVTX1_2_.out ),
    .TE_B(_0243_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_8 _1401_ (.A(\mux_left_track_9.INVTX1_3_.out ),
    .TE_B(_0244_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1402_ (.A(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0245_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1403_ (.A(\mux_left_track_33.INVTX1_7_.out ),
    .TE_B(_0246_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1404_ (.A(\mux_right_track_0.INVTX1_4_.out ),
    .TE_B(_0247_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_8 _1405_ (.A(\mux_bottom_track_1.INVTX1_0_.out ),
    .TE_B(_0248_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1406_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0249_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1407_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0250_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1408_ (.A(net177),
    .TE_B(_0251_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1409_ (.A(\mux_bottom_track_9.INVTX1_8_.out ),
    .TE_B(_0252_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1410_ (.A(\mux_bottom_track_9.INVTX1_9_.out ),
    .TE_B(_0253_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1411_ (.A(\mux_bottom_track_9.INVTX1_11_.out ),
    .TE_B(_0254_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1412_ (.A(\mux_left_track_9.INVTX1_7_.out ),
    .TE_B(_0255_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1413_ (.A(\mux_left_track_9.INVTX1_9_.out ),
    .TE_B(_0256_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1414_ (.A(\mux_left_track_25.INVTX1_9_.out ),
    .TE_B(_0257_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1415_ (.A(\mux_left_track_1.INVTX1_1_.out ),
    .TE_B(_0258_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1416_ (.A(\mux_bottom_track_9.INVTX1_1_.out ),
    .TE_B(_0259_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1417_ (.A(\mux_bottom_track_9.INVTX1_2_.out ),
    .TE_B(_0260_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1418_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0261_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1419_ (.A(\mux_left_track_9.INVTX1_10_.out ),
    .TE_B(_0262_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1420_ (.A(\mux_right_track_8.INVTX1_4_.out ),
    .TE_B(_0263_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1421_ (.A(\mux_bottom_track_9.INVTX1_0_.out ),
    .TE_B(_0264_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1422_ (.A(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0265_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1423_ (.A(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0266_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1424_ (.A(net178),
    .TE_B(_0267_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1425_ (.A(\mux_bottom_track_17.INVTX1_8_.out ),
    .TE_B(_0268_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1426_ (.A(\mux_bottom_track_17.INVTX1_9_.out ),
    .TE_B(_0269_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1427_ (.A(\mux_bottom_track_17.INVTX1_11_.out ),
    .TE_B(_0270_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1428_ (.A(\mux_left_track_17.INVTX1_7_.out ),
    .TE_B(_0271_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1429_ (.A(\mux_left_track_17.INVTX1_8_.out ),
    .TE_B(_0272_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1430_ (.A(\mux_left_track_17.INVTX1_9_.out ),
    .TE_B(_0273_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1431_ (.A(\mux_left_track_33.INVTX1_1_.out ),
    .TE_B(_0274_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1432_ (.A(\mux_bottom_track_17.INVTX1_1_.out ),
    .TE_B(_0275_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1433_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_0276_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1434_ (.A(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0277_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1435_ (.A(\mux_left_track_17.INVTX1_10_.out ),
    .TE_B(_0278_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1436_ (.A(\mux_right_track_16.INVTX1_4_.out ),
    .TE_B(_0279_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1437_ (.A(\mux_bottom_track_17.INVTX1_0_.out ),
    .TE_B(_0280_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1438_ (.A(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0281_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1439_ (.A(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0282_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1440_ (.A(net179),
    .TE_B(_0283_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1441_ (.A(\mux_bottom_track_25.INVTX1_8_.out ),
    .TE_B(_0284_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1442_ (.A(\mux_bottom_track_25.INVTX1_9_.out ),
    .TE_B(_0285_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1443_ (.A(\mux_bottom_track_25.INVTX1_10_.out ),
    .TE_B(_0286_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1444_ (.A(\mux_left_track_9.INVTX1_8_.out ),
    .TE_B(_0287_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1445_ (.A(\mux_left_track_25.INVTX1_7_.out ),
    .TE_B(_0288_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1446_ (.A(\mux_left_track_25.INVTX1_8_.out ),
    .TE_B(_0289_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1447_ (.A(\mux_bottom_track_25.INVTX1_1_.out ),
    .TE_B(_0290_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1448_ (.A(\mux_left_track_25.INVTX1_2_.out ),
    .TE_B(_0291_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1449_ (.A(\mux_bottom_track_25.INVTX1_2_.out ),
    .TE_B(_0292_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1450_ (.A(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0293_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1451_ (.A(\mux_left_track_25.INVTX1_10_.out ),
    .TE_B(_0294_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1452_ (.A(\mux_right_track_24.INVTX1_4_.out ),
    .TE_B(_0295_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1453_ (.A(\mux_bottom_track_25.INVTX1_0_.out ),
    .TE_B(_0296_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1454_ (.A(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0297_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1455_ (.A(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0298_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1456_ (.A(net180),
    .TE_B(_0299_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1457_ (.A(\mux_bottom_track_1.INVTX1_9_.out ),
    .TE_B(_0300_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1458_ (.A(\mux_bottom_track_1.INVTX1_10_.out ),
    .TE_B(_0301_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1459_ (.A(\mux_bottom_track_1.INVTX1_11_.out ),
    .TE_B(_0302_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1460_ (.A(\mux_bottom_track_1.INVTX1_5_.out ),
    .TE_B(_0303_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1461_ (.A(\mux_bottom_track_1.INVTX1_6_.out ),
    .TE_B(_0304_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1462_ (.A(\mux_bottom_track_1.INVTX1_7_.out ),
    .TE_B(_0305_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1463_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_0306_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1464_ (.A(\mux_bottom_track_1.INVTX1_2_.out ),
    .TE_B(_0307_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1465_ (.A(\mux_bottom_track_1.INVTX1_3_.out ),
    .TE_B(_0308_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1466_ (.A(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0309_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1467_ (.A(\mux_bottom_track_1.INVTX1_8_.out ),
    .TE_B(_0310_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1468_ (.A(\mux_bottom_track_1.INVTX1_4_.out ),
    .TE_B(_0311_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1469_ (.A(\mux_bottom_track_1.INVTX1_0_.out ),
    .TE_B(_0312_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1470_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0313_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1471_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0314_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1472_ (.A(net181),
    .TE_B(_0315_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1473_ (.A(\mux_bottom_track_9.INVTX1_9_.out ),
    .TE_B(_0316_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1474_ (.A(\mux_bottom_track_9.INVTX1_10_.out ),
    .TE_B(_0317_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1475_ (.A(\mux_bottom_track_9.INVTX1_11_.out ),
    .TE_B(_0318_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1476_ (.A(\mux_bottom_track_9.INVTX1_5_.out ),
    .TE_B(_0319_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1477_ (.A(\mux_bottom_track_9.INVTX1_6_.out ),
    .TE_B(_0320_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1478_ (.A(\mux_bottom_track_9.INVTX1_7_.out ),
    .TE_B(_0321_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1479_ (.A(\mux_bottom_track_9.INVTX1_1_.out ),
    .TE_B(_0322_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1480_ (.A(\mux_bottom_track_9.INVTX1_2_.out ),
    .TE_B(_0323_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1481_ (.A(\mux_bottom_track_9.INVTX1_3_.out ),
    .TE_B(_0324_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1482_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0325_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1483_ (.A(\mux_bottom_track_9.INVTX1_8_.out ),
    .TE_B(_0326_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1484_ (.A(\mux_bottom_track_9.INVTX1_4_.out ),
    .TE_B(_0327_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1485_ (.A(\mux_bottom_track_9.INVTX1_0_.out ),
    .TE_B(_0328_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1486_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0329_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1487_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0330_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1488_ (.A(net182),
    .TE_B(_0331_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1489_ (.A(\mux_bottom_track_17.INVTX1_9_.out ),
    .TE_B(_0332_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1490_ (.A(\mux_bottom_track_17.INVTX1_10_.out ),
    .TE_B(_0333_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1491_ (.A(\mux_bottom_track_17.INVTX1_11_.out ),
    .TE_B(_0334_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1492_ (.A(\mux_bottom_track_17.INVTX1_5_.out ),
    .TE_B(_0335_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1493_ (.A(\mux_bottom_track_17.INVTX1_6_.out ),
    .TE_B(_0336_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1494_ (.A(\mux_bottom_track_17.INVTX1_7_.out ),
    .TE_B(_0337_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1495_ (.A(\mux_bottom_track_17.INVTX1_1_.out ),
    .TE_B(_0338_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1496_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_0339_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1497_ (.A(\mux_bottom_track_17.INVTX1_3_.out ),
    .TE_B(_0340_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1498_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0341_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1499_ (.A(\mux_bottom_track_17.INVTX1_8_.out ),
    .TE_B(_0342_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1500_ (.A(\mux_bottom_track_17.INVTX1_4_.out ),
    .TE_B(_0343_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1501_ (.A(\mux_bottom_track_17.INVTX1_0_.out ),
    .TE_B(_0344_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1502_ (.A(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0345_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1503_ (.A(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0346_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1504_ (.A(net183),
    .TE_B(_0347_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1505_ (.A(\mux_bottom_track_25.INVTX1_9_.out ),
    .TE_B(_0348_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1506_ (.A(\mux_bottom_track_25.INVTX1_10_.out ),
    .TE_B(_0349_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1507_ (.A(\mux_bottom_track_25.INVTX1_11_.out ),
    .TE_B(_0350_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1508_ (.A(\mux_bottom_track_25.INVTX1_5_.out ),
    .TE_B(_0351_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1509_ (.A(\mux_bottom_track_25.INVTX1_6_.out ),
    .TE_B(_0352_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1510_ (.A(\mux_bottom_track_25.INVTX1_7_.out ),
    .TE_B(_0353_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1511_ (.A(\mux_bottom_track_25.INVTX1_1_.out ),
    .TE_B(_0354_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1512_ (.A(\mux_bottom_track_25.INVTX1_2_.out ),
    .TE_B(_0355_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1513_ (.A(\mux_bottom_track_25.INVTX1_3_.out ),
    .TE_B(_0356_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1514_ (.A(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0357_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1515_ (.A(\mux_bottom_track_25.INVTX1_8_.out ),
    .TE_B(_0358_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1516_ (.A(\mux_bottom_track_25.INVTX1_4_.out ),
    .TE_B(_0359_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1517_ (.A(\mux_bottom_track_25.INVTX1_0_.out ),
    .TE_B(_0360_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1518_ (.A(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0361_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1519_ (.A(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0362_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1520_ (.A(net184),
    .TE_B(_0363_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1521_ (.A(\mux_left_track_1.INVTX1_9_.out ),
    .TE_B(_0364_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1522_ (.A(\mux_left_track_1.INVTX1_10_.out ),
    .TE_B(_0365_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1523_ (.A(\mux_left_track_1.INVTX1_11_.out ),
    .TE_B(_0366_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1524_ (.A(\mux_bottom_track_1.INVTX1_4_.out ),
    .TE_B(_0367_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1525_ (.A(\mux_bottom_track_1.INVTX1_5_.out ),
    .TE_B(_0368_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1526_ (.A(\mux_left_track_1.INVTX1_7_.out ),
    .TE_B(_0369_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1527_ (.A(\mux_left_track_1.INVTX1_1_.out ),
    .TE_B(_0370_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1528_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_0371_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1529_ (.A(\mux_bottom_track_1.INVTX1_2_.out ),
    .TE_B(_0372_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1530_ (.A(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0373_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1531_ (.A(\mux_left_track_1.INVTX1_8_.out ),
    .TE_B(_0374_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1532_ (.A(\mux_bottom_track_1.INVTX1_3_.out ),
    .TE_B(_0375_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1533_ (.A(\mux_bottom_track_1.INVTX1_0_.out ),
    .TE_B(_0376_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1534_ (.A(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0377_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1535_ (.A(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0378_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1536_ (.A(net185),
    .TE_B(_0379_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1537_ (.A(\mux_left_track_9.INVTX1_9_.out ),
    .TE_B(_0380_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1538_ (.A(\mux_left_track_9.INVTX1_10_.out ),
    .TE_B(_0381_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1539_ (.A(\mux_left_track_9.INVTX1_11_.out ),
    .TE_B(_0382_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1540_ (.A(\mux_bottom_track_9.INVTX1_4_.out ),
    .TE_B(_0383_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1541_ (.A(\mux_bottom_track_9.INVTX1_6_.out ),
    .TE_B(_0384_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1542_ (.A(\mux_left_track_9.INVTX1_7_.out ),
    .TE_B(_0385_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1543_ (.A(\mux_bottom_track_9.INVTX1_1_.out ),
    .TE_B(_0386_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1544_ (.A(\mux_bottom_track_9.INVTX1_2_.out ),
    .TE_B(_0387_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1545_ (.A(\mux_left_track_9.INVTX1_3_.out ),
    .TE_B(_0388_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1546_ (.A(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0389_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1547_ (.A(\mux_left_track_9.INVTX1_8_.out ),
    .TE_B(_0390_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1548_ (.A(\mux_bottom_track_9.INVTX1_3_.out ),
    .TE_B(_0391_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1549_ (.A(\mux_bottom_track_9.INVTX1_0_.out ),
    .TE_B(_0392_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1550_ (.A(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0393_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1551_ (.A(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0394_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1552_ (.A(net186),
    .TE_B(_0395_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1553_ (.A(\mux_left_track_17.INVTX1_9_.out ),
    .TE_B(_0396_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1554_ (.A(\mux_left_track_17.INVTX1_10_.out ),
    .TE_B(_0397_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1555_ (.A(\mux_left_track_17.INVTX1_11_.out ),
    .TE_B(_0398_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1556_ (.A(\mux_bottom_track_17.INVTX1_5_.out ),
    .TE_B(_0399_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1557_ (.A(\mux_bottom_track_17.INVTX1_6_.out ),
    .TE_B(_0400_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1558_ (.A(\mux_left_track_17.INVTX1_7_.out ),
    .TE_B(_0401_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1559_ (.A(\mux_bottom_track_17.INVTX1_1_.out ),
    .TE_B(_0402_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1560_ (.A(\mux_left_track_17.INVTX1_2_.out ),
    .TE_B(_0403_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1561_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_0404_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1562_ (.A(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0405_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1563_ (.A(\mux_left_track_17.INVTX1_8_.out ),
    .TE_B(_0406_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1564_ (.A(\mux_bottom_track_17.INVTX1_3_.out ),
    .TE_B(_0407_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1565_ (.A(\mux_bottom_track_17.INVTX1_0_.out ),
    .TE_B(_0408_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1566_ (.A(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ),
    .TE_B(_0409_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1567_ (.A(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ),
    .TE_B(_0410_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1568_ (.A(net187),
    .TE_B(_0411_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_8 _1569_ (.A(\mux_left_track_25.INVTX1_9_.out ),
    .TE_B(_0412_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_8 _1570_ (.A(\mux_left_track_25.INVTX1_10_.out ),
    .TE_B(_0413_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_8 _1571_ (.A(\mux_left_track_25.INVTX1_11_.out ),
    .TE_B(_0414_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1572_ (.A(\mux_bottom_track_25.INVTX1_5_.out ),
    .TE_B(_0415_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1573_ (.A(\mux_bottom_track_25.INVTX1_6_.out ),
    .TE_B(_0416_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1574_ (.A(\mux_left_track_25.INVTX1_7_.out ),
    .TE_B(_0417_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1575_ (.A(\mux_bottom_track_25.INVTX1_1_.out ),
    .TE_B(_0418_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1576_ (.A(\mux_left_track_25.INVTX1_2_.out ),
    .TE_B(_0419_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1577_ (.A(\mux_bottom_track_25.INVTX1_2_.out ),
    .TE_B(_0420_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1578_ (.A(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ),
    .TE_B(_0421_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out ));
 sky130_fd_sc_hd__ebufn_8 _1579_ (.A(\mux_left_track_25.INVTX1_8_.out ),
    .TE_B(_0422_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1580_ (.A(\mux_bottom_track_25.INVTX1_4_.out ),
    .TE_B(_0423_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1581_ (.A(\mux_bottom_track_25.INVTX1_0_.out ),
    .TE_B(_0424_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1582_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_0425_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1583_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_0426_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1584_ (.A(\mux_bottom_track_33.INVTX1_7_.out ),
    .TE_B(_0427_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1585_ (.A(net188),
    .TE_B(_0428_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1586_ (.A(\mux_left_track_33.INVTX1_6_.out ),
    .TE_B(_0429_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1587_ (.A(\mux_bottom_track_33.INVTX1_6_.out ),
    .TE_B(_0430_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1588_ (.A(\mux_bottom_track_33.INVTX1_2_.out ),
    .TE_B(_0431_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1589_ (.A(\mux_bottom_track_33.INVTX1_3_.out ),
    .TE_B(_0432_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1590_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0433_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1591_ (.A(\mux_bottom_track_1.INVTX1_10_.out ),
    .TE_B(_0434_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1592_ (.A(\mux_left_track_33.INVTX1_5_.out ),
    .TE_B(_0435_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1593_ (.A(\mux_bottom_track_25.INVTX1_3_.out ),
    .TE_B(_0436_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1594_ (.A(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_0437_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1595_ (.A(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_0438_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1596_ (.A(\mux_bottom_track_33.INVTX1_7_.out ),
    .TE_B(_0439_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1597_ (.A(net189),
    .TE_B(_0440_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1598_ (.A(\mux_left_track_33.INVTX1_6_.out ),
    .TE_B(_0441_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1599_ (.A(\mux_left_track_1.INVTX1_10_.out ),
    .TE_B(_0442_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1600_ (.A(\mux_bottom_track_33.INVTX1_1_.out ),
    .TE_B(_0443_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1601_ (.A(\mux_left_track_17.INVTX1_2_.out ),
    .TE_B(_0444_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1602_ (.A(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0445_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1603_ (.A(\mux_bottom_track_33.INVTX1_6_.out ),
    .TE_B(_0446_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1604_ (.A(\mux_left_track_33.INVTX1_5_.out ),
    .TE_B(_0447_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1605_ (.A(\mux_bottom_track_33.INVTX1_0_.out ),
    .TE_B(_0448_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1606_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_0449_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _1607_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_0450_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1608_ (.A(\mux_bottom_track_33.INVTX1_7_.out ),
    .TE_B(_0451_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1609_ (.A(net190),
    .TE_B(_0452_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1610_ (.A(\mux_bottom_track_33.INVTX1_4_.out ),
    .TE_B(_0453_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_4 _1611_ (.A(\mux_bottom_track_33.INVTX1_5_.out ),
    .TE_B(_0454_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1612_ (.A(\mux_bottom_track_33.INVTX1_1_.out ),
    .TE_B(_0455_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1613_ (.A(\mux_bottom_track_33.INVTX1_2_.out ),
    .TE_B(_0456_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1614_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0457_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1615_ (.A(\mux_bottom_track_33.INVTX1_6_.out ),
    .TE_B(_0458_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _1616_ (.A(\mux_bottom_track_33.INVTX1_3_.out ),
    .TE_B(_0459_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1617_ (.A(\mux_bottom_track_33.INVTX1_0_.out ),
    .TE_B(_0460_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1618_ (.A(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_0461_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _1619_ (.A(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_0462_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_1 _1620_ (.A(\mux_left_track_33.INVTX1_7_.out ),
    .TE_B(_0463_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1621_ (.A(net191),
    .TE_B(_0464_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1622_ (.A(\mux_bottom_track_33.INVTX1_3_.out ),
    .TE_B(_0465_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1623_ (.A(\mux_left_track_33.INVTX1_5_.out ),
    .TE_B(_0466_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1624_ (.A(\mux_left_track_33.INVTX1_1_.out ),
    .TE_B(_0467_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1625_ (.A(\mux_bottom_track_33.INVTX1_1_.out ),
    .TE_B(_0468_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1626_ (.A(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_0469_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_1 _1627_ (.A(\mux_left_track_33.INVTX1_6_.out ),
    .TE_B(_0470_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1628_ (.A(\mux_bottom_track_33.INVTX1_2_.out ),
    .TE_B(_0471_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1629_ (.A(\mux_bottom_track_33.INVTX1_0_.out ),
    .TE_B(_0472_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ccff_head),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(chanx_left_in[0]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(chanx_left_in[10]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(chanx_left_in[11]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(chanx_left_in[12]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(chanx_left_in[13]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(chanx_left_in[14]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(chanx_left_in[15]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(chanx_left_in[16]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(chanx_left_in[17]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(chanx_left_in[18]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(chanx_left_in[1]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(chanx_left_in[2]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(chanx_left_in[3]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(chanx_left_in[4]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(chanx_left_in[5]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(chanx_left_in[6]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(chanx_left_in[7]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(chanx_left_in[8]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(chanx_left_in[9]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(chanx_right_in[0]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(chanx_right_in[10]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(chanx_right_in[11]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(chanx_right_in[12]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(chanx_right_in[13]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(chanx_right_in[14]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(chanx_right_in[15]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(chanx_right_in[16]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(chanx_right_in[17]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(chanx_right_in[18]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(chanx_right_in[1]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(chanx_right_in[2]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(chanx_right_in[3]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(chanx_right_in[4]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(chanx_right_in[5]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(chanx_right_in[6]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(chanx_right_in[7]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(chanx_right_in[8]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(chanx_right_in[9]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(chany_bottom_in[0]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(chany_bottom_in[10]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(chany_bottom_in[11]),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(chany_bottom_in[12]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(chany_bottom_in[13]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(chany_bottom_in[14]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(chany_bottom_in[15]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(chany_bottom_in[16]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(chany_bottom_in[17]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(chany_bottom_in[18]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(chany_bottom_in[1]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(chany_bottom_in[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(chany_bottom_in[3]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(chany_bottom_in[4]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(chany_bottom_in[5]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(chany_bottom_in[6]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(chany_bottom_in[7]),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(chany_bottom_in[8]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(chany_bottom_in[9]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(chany_top_in[0]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(chany_top_in[10]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(chany_top_in[11]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(chany_top_in[12]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(chany_top_in[13]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(chany_top_in[14]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(chany_top_in[15]),
    .X(net69));
 sky130_fd_sc_hd__dlymetal6s2s_1 input70 (.A(chany_top_in[16]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input71 (.A(chany_top_in[17]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(chany_top_in[18]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(chany_top_in[1]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(chany_top_in[2]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(chany_top_in[3]),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 input76 (.A(chany_top_in[4]),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 input77 (.A(chany_top_in[5]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(chany_top_in[6]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(chany_top_in[7]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(chany_top_in[8]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(chany_top_in[9]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(pReset),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_),
    .X(net94));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(ccff_tail));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(chanx_left_out[0]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(chanx_left_out[10]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(chanx_left_out[11]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(chanx_left_out[12]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(chanx_left_out[13]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(chanx_left_out[14]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(chanx_left_out[15]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(chanx_left_out[16]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(chanx_left_out[17]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(chanx_left_out[18]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(chanx_left_out[1]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(chanx_left_out[2]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(chanx_left_out[3]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(chanx_left_out[4]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(chanx_left_out[5]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(chanx_left_out[6]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(chanx_left_out[7]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(chanx_left_out[8]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(chanx_left_out[9]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(chanx_right_out[0]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(chanx_right_out[10]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(chanx_right_out[11]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(chanx_right_out[12]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(chanx_right_out[13]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(chanx_right_out[14]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(chanx_right_out[15]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(chanx_right_out[16]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(chanx_right_out[17]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(chanx_right_out[18]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(chanx_right_out[1]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(chanx_right_out[2]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(chanx_right_out[3]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(chanx_right_out[4]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(chanx_right_out[5]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(chanx_right_out[6]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(chanx_right_out[7]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(chanx_right_out[8]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(chanx_right_out[9]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(chany_bottom_out[0]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(chany_bottom_out[10]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(chany_bottom_out[11]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(chany_bottom_out[12]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(chany_bottom_out[13]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(chany_bottom_out[14]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(chany_bottom_out[15]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(chany_bottom_out[16]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(chany_bottom_out[17]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(chany_bottom_out[18]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(chany_bottom_out[1]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(chany_bottom_out[2]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(chany_bottom_out[3]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(chany_bottom_out[4]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(chany_bottom_out[5]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(chany_bottom_out[6]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(chany_bottom_out[7]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(chany_bottom_out[8]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(chany_bottom_out[9]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(chany_top_out[0]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(chany_top_out[10]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(chany_top_out[11]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(chany_top_out[12]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(chany_top_out[13]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(chany_top_out[14]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(chany_top_out[15]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(chany_top_out[16]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(chany_top_out[17]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(chany_top_out[18]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(chany_top_out[1]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(chany_top_out[2]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(chany_top_out[3]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(chany_top_out[4]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(chany_top_out[5]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(chany_top_out[6]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(chany_top_out[7]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(chany_top_out[8]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(chany_top_out[9]));
 sky130_fd_sc_hd__conb_1 _1328__172 (.HI(net172));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_0_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_1_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_2_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_3_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_4_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_5_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_6_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_7_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_8_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_9_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_10_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_11_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_12_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_13_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_14_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_15_0_prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\mux_bottom_track_17.INVTX1_4_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\mux_bottom_track_17.INVTX1_4_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\mux_bottom_track_33.INVTX1_4_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\mux_bottom_track_33.INVTX1_4_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\mem_bottom_track_17.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\mem_top_track_0.DFFR_7_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net30));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
endmodule

