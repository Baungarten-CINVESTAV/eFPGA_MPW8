magic
tech sky130A
magscale 1 2
timestamp 1672417827
<< viali >>
rect 1869 37213 1903 37247
rect 2329 37213 2363 37247
rect 2973 37213 3007 37247
rect 4261 37213 4295 37247
rect 5549 37213 5583 37247
rect 7389 37213 7423 37247
rect 9321 37213 9355 37247
rect 10609 37213 10643 37247
rect 11897 37213 11931 37247
rect 13001 37213 13035 37247
rect 15209 37213 15243 37247
rect 16865 37213 16899 37247
rect 18153 37213 18187 37247
rect 19441 37213 19475 37247
rect 20913 37213 20947 37247
rect 22845 37213 22879 37247
rect 24593 37213 24627 37247
rect 25881 37213 25915 37247
rect 27353 37213 27387 37247
rect 29745 37213 29779 37247
rect 30665 37213 30699 37247
rect 32505 37213 32539 37247
rect 33793 37213 33827 37247
rect 35081 37213 35115 37247
rect 36921 37213 36955 37247
rect 38025 37213 38059 37247
rect 1685 37077 1719 37111
rect 2513 37077 2547 37111
rect 3157 37077 3191 37111
rect 4077 37077 4111 37111
rect 5365 37077 5399 37111
rect 7205 37077 7239 37111
rect 9137 37077 9171 37111
rect 10425 37077 10459 37111
rect 11713 37077 11747 37111
rect 13185 37077 13219 37111
rect 15025 37077 15059 37111
rect 17049 37077 17083 37111
rect 18337 37077 18371 37111
rect 19625 37077 19659 37111
rect 20729 37077 20763 37111
rect 22661 37077 22695 37111
rect 24777 37077 24811 37111
rect 26065 37077 26099 37111
rect 27169 37077 27203 37111
rect 29929 37077 29963 37111
rect 30481 37077 30515 37111
rect 32321 37077 32355 37111
rect 33609 37077 33643 37111
rect 34897 37077 34931 37111
rect 36737 37077 36771 37111
rect 38209 37077 38243 37111
rect 1685 36873 1719 36907
rect 1869 36737 1903 36771
rect 36921 36737 36955 36771
rect 37565 36737 37599 36771
rect 36737 36533 36771 36567
rect 37565 36533 37599 36567
rect 38209 36329 38243 36363
rect 1593 36125 1627 36159
rect 37381 36125 37415 36159
rect 38025 36125 38059 36159
rect 1777 35989 1811 36023
rect 37565 35989 37599 36023
rect 5733 35785 5767 35819
rect 16865 35785 16899 35819
rect 5917 35649 5951 35683
rect 17049 35649 17083 35683
rect 38301 35649 38335 35683
rect 38117 35445 38151 35479
rect 6469 35241 6503 35275
rect 17693 35241 17727 35275
rect 17049 35173 17083 35207
rect 6653 35037 6687 35071
rect 16865 35037 16899 35071
rect 17509 35037 17543 35071
rect 38025 35037 38059 35071
rect 38209 34901 38243 34935
rect 6745 34697 6779 34731
rect 15485 34697 15519 34731
rect 21373 34697 21407 34731
rect 22845 34697 22879 34731
rect 25789 34697 25823 34731
rect 1869 34561 1903 34595
rect 6929 34561 6963 34595
rect 14841 34561 14875 34595
rect 15669 34561 15703 34595
rect 20729 34561 20763 34595
rect 21189 34561 21223 34595
rect 22661 34561 22695 34595
rect 25605 34561 25639 34595
rect 33241 34561 33275 34595
rect 14933 34493 14967 34527
rect 20637 34493 20671 34527
rect 33149 34493 33183 34527
rect 1685 34357 1719 34391
rect 9873 33949 9907 33983
rect 10333 33949 10367 33983
rect 30297 33949 30331 33983
rect 9781 33813 9815 33847
rect 10425 33813 10459 33847
rect 30205 33813 30239 33847
rect 14289 33609 14323 33643
rect 14197 33473 14231 33507
rect 19993 33473 20027 33507
rect 29377 33473 29411 33507
rect 38025 33473 38059 33507
rect 29285 33337 29319 33371
rect 38209 33337 38243 33371
rect 19901 33269 19935 33303
rect 1593 32861 1627 32895
rect 1777 32725 1811 32759
rect 33977 32521 34011 32555
rect 5273 32385 5307 32419
rect 33793 32385 33827 32419
rect 5365 32181 5399 32215
rect 38117 31909 38151 31943
rect 23213 31773 23247 31807
rect 23305 31773 23339 31807
rect 38301 31773 38335 31807
rect 16957 31433 16991 31467
rect 16865 31297 16899 31331
rect 3985 30889 4019 30923
rect 6193 30889 6227 30923
rect 35081 30889 35115 30923
rect 1777 30821 1811 30855
rect 1593 30685 1627 30719
rect 4169 30685 4203 30719
rect 6285 30685 6319 30719
rect 8309 30685 8343 30719
rect 34897 30685 34931 30719
rect 8217 30549 8251 30583
rect 11805 30277 11839 30311
rect 20913 30277 20947 30311
rect 2697 30209 2731 30243
rect 6561 30209 6595 30243
rect 11897 30209 11931 30243
rect 20821 30209 20855 30243
rect 27353 30209 27387 30243
rect 29285 30209 29319 30243
rect 33333 30209 33367 30243
rect 38301 30209 38335 30243
rect 2421 30141 2455 30175
rect 33517 30073 33551 30107
rect 6653 30005 6687 30039
rect 27261 30005 27295 30039
rect 29193 30005 29227 30039
rect 38117 30005 38151 30039
rect 12081 29801 12115 29835
rect 16497 29801 16531 29835
rect 17141 29801 17175 29835
rect 24685 29801 24719 29835
rect 2605 29665 2639 29699
rect 5181 29665 5215 29699
rect 1869 29597 1903 29631
rect 2789 29597 2823 29631
rect 5089 29597 5123 29631
rect 5733 29597 5767 29631
rect 6377 29597 6411 29631
rect 12173 29597 12207 29631
rect 16405 29597 16439 29631
rect 17049 29597 17083 29631
rect 24593 29597 24627 29631
rect 25513 29597 25547 29631
rect 30573 29597 30607 29631
rect 5825 29529 5859 29563
rect 1685 29461 1719 29495
rect 6469 29461 6503 29495
rect 25421 29461 25455 29495
rect 30481 29461 30515 29495
rect 1593 29121 1627 29155
rect 2789 29121 2823 29155
rect 4353 29121 4387 29155
rect 4997 29121 5031 29155
rect 38025 29121 38059 29155
rect 2513 29053 2547 29087
rect 5089 29053 5123 29087
rect 1777 28985 1811 29019
rect 4445 28985 4479 29019
rect 38209 28985 38243 29019
rect 4077 28713 4111 28747
rect 19717 28713 19751 28747
rect 33425 28713 33459 28747
rect 2605 28509 2639 28543
rect 4169 28509 4203 28543
rect 16313 28509 16347 28543
rect 19625 28509 19659 28543
rect 33333 28509 33367 28543
rect 34161 28509 34195 28543
rect 2329 28441 2363 28475
rect 16497 28373 16531 28407
rect 34069 28373 34103 28407
rect 1961 28033 1995 28067
rect 2605 28033 2639 28067
rect 3525 28033 3559 28067
rect 4169 28033 4203 28067
rect 6745 28033 6779 28067
rect 15853 28033 15887 28067
rect 16865 28033 16899 28067
rect 33793 28033 33827 28067
rect 2053 27829 2087 27863
rect 2697 27829 2731 27863
rect 3617 27829 3651 27863
rect 4261 27829 4295 27863
rect 6837 27829 6871 27863
rect 16037 27829 16071 27863
rect 16957 27829 16991 27863
rect 33701 27829 33735 27863
rect 16681 27557 16715 27591
rect 17509 27557 17543 27591
rect 2329 27489 2363 27523
rect 16865 27489 16899 27523
rect 1777 27421 1811 27455
rect 2421 27421 2455 27455
rect 3065 27421 3099 27455
rect 4169 27421 4203 27455
rect 4629 27421 4663 27455
rect 6745 27421 6779 27455
rect 7389 27421 7423 27455
rect 9137 27421 9171 27455
rect 13277 27421 13311 27455
rect 15945 27421 15979 27455
rect 17049 27421 17083 27455
rect 17693 27421 17727 27455
rect 18153 27353 18187 27387
rect 1685 27285 1719 27319
rect 2881 27285 2915 27319
rect 4077 27285 4111 27319
rect 4721 27285 4755 27319
rect 5917 27285 5951 27319
rect 6561 27285 6595 27319
rect 7205 27285 7239 27319
rect 9229 27285 9263 27319
rect 13093 27285 13127 27319
rect 15761 27285 15795 27319
rect 3617 27081 3651 27115
rect 6929 27081 6963 27115
rect 16865 27081 16899 27115
rect 29837 27081 29871 27115
rect 1593 26945 1627 26979
rect 2513 26945 2547 26979
rect 2973 26945 3007 26979
rect 3801 26945 3835 26979
rect 4445 26945 4479 26979
rect 4905 26945 4939 26979
rect 8033 26945 8067 26979
rect 8677 26945 8711 26979
rect 11713 26945 11747 26979
rect 12633 26945 12667 26979
rect 13369 26945 13403 26979
rect 14013 26945 14047 26979
rect 14841 26945 14875 26979
rect 16313 26945 16347 26979
rect 17325 26945 17359 26979
rect 18429 26945 18463 26979
rect 19073 26945 19107 26979
rect 29745 26945 29779 26979
rect 38025 26945 38059 26979
rect 7389 26877 7423 26911
rect 7573 26877 7607 26911
rect 15485 26877 15519 26911
rect 17509 26877 17543 26911
rect 8125 26809 8159 26843
rect 11897 26809 11931 26843
rect 1777 26741 1811 26775
rect 2421 26741 2455 26775
rect 3065 26741 3099 26775
rect 4261 26741 4295 26775
rect 4997 26741 5031 26775
rect 8861 26741 8895 26775
rect 12725 26741 12759 26775
rect 13553 26741 13587 26775
rect 14197 26741 14231 26775
rect 14933 26741 14967 26775
rect 16129 26741 16163 26775
rect 18245 26741 18279 26775
rect 18889 26741 18923 26775
rect 38209 26741 38243 26775
rect 4997 26537 5031 26571
rect 6285 26537 6319 26571
rect 17049 26537 17083 26571
rect 18153 26537 18187 26571
rect 36277 26537 36311 26571
rect 12449 26469 12483 26503
rect 17509 26469 17543 26503
rect 5917 26401 5951 26435
rect 6101 26401 6135 26435
rect 8033 26401 8067 26435
rect 9229 26401 9263 26435
rect 18797 26401 18831 26435
rect 2329 26333 2363 26367
rect 2789 26333 2823 26367
rect 4537 26333 4571 26367
rect 5181 26333 5215 26367
rect 8217 26333 8251 26367
rect 9137 26333 9171 26367
rect 9965 26333 9999 26367
rect 10977 26333 11011 26367
rect 11621 26333 11655 26367
rect 12265 26333 12299 26367
rect 13093 26333 13127 26367
rect 13553 26333 13587 26367
rect 14381 26333 14415 26367
rect 15577 26333 15611 26367
rect 16865 26333 16899 26367
rect 17693 26333 17727 26367
rect 18613 26333 18647 26367
rect 19441 26333 19475 26367
rect 36093 26333 36127 26367
rect 2237 26265 2271 26299
rect 2881 26265 2915 26299
rect 11069 26265 11103 26299
rect 11713 26265 11747 26299
rect 14473 26265 14507 26299
rect 4353 26197 4387 26231
rect 7573 26197 7607 26231
rect 9781 26197 9815 26231
rect 13001 26197 13035 26231
rect 13737 26197 13771 26231
rect 15761 26197 15795 26231
rect 16221 26197 16255 26231
rect 19533 26197 19567 26231
rect 3801 25993 3835 26027
rect 7665 25993 7699 26027
rect 11897 25993 11931 26027
rect 20085 25993 20119 26027
rect 20821 25993 20855 26027
rect 29653 25993 29687 26027
rect 9045 25925 9079 25959
rect 1593 25857 1627 25891
rect 2421 25857 2455 25891
rect 3249 25857 3283 25891
rect 3893 25857 3927 25891
rect 4537 25857 4571 25891
rect 5181 25857 5215 25891
rect 6009 25857 6043 25891
rect 7205 25857 7239 25891
rect 8309 25857 8343 25891
rect 9137 25857 9171 25891
rect 10241 25857 10275 25891
rect 11161 25857 11195 25891
rect 11713 25857 11747 25891
rect 12541 25857 12575 25891
rect 13185 25857 13219 25891
rect 14105 25857 14139 25891
rect 14565 25857 14599 25891
rect 15485 25857 15519 25891
rect 16129 25857 16163 25891
rect 17509 25857 17543 25891
rect 18521 25857 18555 25891
rect 19441 25855 19475 25889
rect 20269 25857 20303 25891
rect 20729 25857 20763 25891
rect 29561 25857 29595 25891
rect 8125 25789 8159 25823
rect 10057 25789 10091 25823
rect 15577 25789 15611 25823
rect 17325 25789 17359 25823
rect 18705 25789 18739 25823
rect 2513 25721 2547 25755
rect 5825 25721 5859 25755
rect 13001 25721 13035 25755
rect 1777 25653 1811 25687
rect 3065 25653 3099 25687
rect 4445 25653 4479 25687
rect 5365 25653 5399 25687
rect 7021 25653 7055 25687
rect 9597 25653 9631 25687
rect 10977 25653 11011 25687
rect 12357 25653 12391 25687
rect 13921 25653 13955 25687
rect 14749 25653 14783 25687
rect 16221 25653 16255 25687
rect 16865 25653 16899 25687
rect 18337 25653 18371 25687
rect 19533 25653 19567 25687
rect 8493 25449 8527 25483
rect 18153 25449 18187 25483
rect 35725 25449 35759 25483
rect 3249 25381 3283 25415
rect 15393 25381 15427 25415
rect 16497 25381 16531 25415
rect 2605 25313 2639 25347
rect 9965 25313 9999 25347
rect 13001 25313 13035 25347
rect 13645 25313 13679 25347
rect 15209 25313 15243 25347
rect 16129 25313 16163 25347
rect 18521 25313 18555 25347
rect 1869 25245 1903 25279
rect 2513 25245 2547 25279
rect 3157 25245 3191 25279
rect 4721 25245 4755 25279
rect 5181 25245 5215 25279
rect 5825 25245 5859 25279
rect 6469 25245 6503 25279
rect 7297 25245 7331 25279
rect 7757 25245 7791 25279
rect 8585 25245 8619 25279
rect 9229 25245 9263 25279
rect 10057 25245 10091 25279
rect 10517 25245 10551 25279
rect 11897 25245 11931 25279
rect 15025 25245 15059 25279
rect 16313 25245 16347 25279
rect 17417 25245 17451 25279
rect 18705 25245 18739 25279
rect 19717 25245 19751 25279
rect 20361 25245 20395 25279
rect 35633 25245 35667 25279
rect 38301 25245 38335 25279
rect 1961 25177 1995 25211
rect 13553 25177 13587 25211
rect 4537 25109 4571 25143
rect 5273 25109 5307 25143
rect 6009 25109 6043 25143
rect 6653 25109 6687 25143
rect 7205 25109 7239 25143
rect 7849 25109 7883 25143
rect 9321 25109 9355 25143
rect 10609 25109 10643 25143
rect 11713 25109 11747 25143
rect 12541 25109 12575 25143
rect 14289 25109 14323 25143
rect 17601 25109 17635 25143
rect 19901 25109 19935 25143
rect 20545 25109 20579 25143
rect 38117 25109 38151 25143
rect 6009 24905 6043 24939
rect 12817 24837 12851 24871
rect 13369 24837 13403 24871
rect 18705 24837 18739 24871
rect 1869 24769 1903 24803
rect 2421 24769 2455 24803
rect 3065 24769 3099 24803
rect 3249 24769 3283 24803
rect 4445 24769 4479 24803
rect 4905 24769 4939 24803
rect 5825 24769 5859 24803
rect 6653 24769 6687 24803
rect 7297 24769 7331 24803
rect 8125 24769 8159 24803
rect 9045 24769 9079 24803
rect 9689 24769 9723 24803
rect 10333 24769 10367 24803
rect 11897 24769 11931 24803
rect 14657 24769 14691 24803
rect 15577 24769 15611 24803
rect 15761 24769 15795 24803
rect 17601 24769 17635 24803
rect 20545 24769 20579 24803
rect 20729 24769 20763 24803
rect 3709 24701 3743 24735
rect 4261 24701 4295 24735
rect 7941 24701 7975 24735
rect 11161 24701 11195 24735
rect 11713 24701 11747 24735
rect 13461 24701 13495 24735
rect 14841 24701 14875 24735
rect 16221 24701 16255 24735
rect 17417 24701 17451 24735
rect 18613 24701 18647 24735
rect 19625 24701 19659 24735
rect 21189 24701 21223 24735
rect 6745 24633 6779 24667
rect 14197 24633 14231 24667
rect 1685 24565 1719 24599
rect 2513 24565 2547 24599
rect 7389 24565 7423 24599
rect 8585 24565 8619 24599
rect 9137 24565 9171 24599
rect 9873 24565 9907 24599
rect 10425 24565 10459 24599
rect 12081 24565 12115 24599
rect 17969 24565 18003 24599
rect 20085 24565 20119 24599
rect 4629 24361 4663 24395
rect 16957 24361 16991 24395
rect 35357 24361 35391 24395
rect 6009 24293 6043 24327
rect 14657 24293 14691 24327
rect 2789 24225 2823 24259
rect 3985 24225 4019 24259
rect 4169 24225 4203 24259
rect 5365 24225 5399 24259
rect 5549 24225 5583 24259
rect 6561 24225 6595 24259
rect 7205 24225 7239 24259
rect 8033 24225 8067 24259
rect 11437 24225 11471 24259
rect 17509 24225 17543 24259
rect 17693 24225 17727 24259
rect 20913 24225 20947 24259
rect 21097 24225 21131 24259
rect 1961 24157 1995 24191
rect 3433 24157 3467 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 10609 24157 10643 24191
rect 11253 24157 11287 24191
rect 13553 24157 13587 24191
rect 16405 24157 16439 24191
rect 16865 24157 16899 24191
rect 18705 24157 18739 24191
rect 35173 24157 35207 24191
rect 2053 24089 2087 24123
rect 6653 24089 6687 24123
rect 7757 24089 7791 24123
rect 7849 24089 7883 24123
rect 15117 24089 15151 24123
rect 15209 24089 15243 24123
rect 20453 24089 20487 24123
rect 3341 24021 3375 24055
rect 9413 24021 9447 24055
rect 10149 24021 10183 24055
rect 10793 24021 10827 24055
rect 11897 24021 11931 24055
rect 13093 24021 13127 24055
rect 13645 24021 13679 24055
rect 16221 24021 16255 24055
rect 18153 24021 18187 24055
rect 18889 24021 18923 24055
rect 19441 24021 19475 24055
rect 1777 23817 1811 23851
rect 4353 23749 4387 23783
rect 7113 23749 7147 23783
rect 7665 23749 7699 23783
rect 7757 23749 7791 23783
rect 12081 23749 12115 23783
rect 18981 23749 19015 23783
rect 19901 23749 19935 23783
rect 1593 23681 1627 23715
rect 2513 23681 2547 23715
rect 2973 23681 3007 23715
rect 3617 23681 3651 23715
rect 4261 23681 4295 23715
rect 5089 23681 5123 23715
rect 5825 23681 5859 23715
rect 8769 23681 8803 23715
rect 9873 23681 9907 23715
rect 10977 23681 11011 23715
rect 13277 23681 13311 23715
rect 13921 23681 13955 23715
rect 14565 23681 14599 23715
rect 15025 23681 15059 23715
rect 16129 23681 16163 23715
rect 17509 23681 17543 23715
rect 18153 23681 18187 23715
rect 20545 23681 20579 23715
rect 33977 23681 34011 23715
rect 38301 23681 38335 23715
rect 8953 23613 8987 23647
rect 9689 23613 9723 23647
rect 11989 23613 12023 23647
rect 15209 23613 15243 23647
rect 16313 23613 16347 23647
rect 17325 23613 17359 23647
rect 18889 23613 18923 23647
rect 3065 23545 3099 23579
rect 3709 23545 3743 23579
rect 8401 23545 8435 23579
rect 12541 23545 12575 23579
rect 20361 23545 20395 23579
rect 2421 23477 2455 23511
rect 4997 23477 5031 23511
rect 5917 23477 5951 23511
rect 10333 23477 10367 23511
rect 11161 23477 11195 23511
rect 13461 23477 13495 23511
rect 14105 23477 14139 23511
rect 15945 23477 15979 23511
rect 16865 23477 16899 23511
rect 18337 23477 18371 23511
rect 33885 23477 33919 23511
rect 38117 23477 38151 23511
rect 7775 23273 7809 23307
rect 12541 23273 12575 23307
rect 14657 23273 14691 23307
rect 20545 23273 20579 23307
rect 4077 23205 4111 23239
rect 1593 23137 1627 23171
rect 10885 23137 10919 23171
rect 11897 23137 11931 23171
rect 12081 23137 12115 23171
rect 13093 23137 13127 23171
rect 13553 23137 13587 23171
rect 16129 23137 16163 23171
rect 18245 23137 18279 23171
rect 18429 23137 18463 23171
rect 20085 23137 20119 23171
rect 3985 23069 4019 23103
rect 4629 23069 4663 23103
rect 8033 23069 8067 23103
rect 10701 23069 10735 23103
rect 15117 23069 15151 23103
rect 15301 23069 15335 23103
rect 17325 23069 17359 23103
rect 19901 23069 19935 23103
rect 20729 23069 20763 23103
rect 1869 23001 1903 23035
rect 9230 23001 9264 23035
rect 9330 23001 9364 23035
rect 9873 23001 9907 23035
rect 13185 23001 13219 23035
rect 16221 23001 16255 23035
rect 16773 23001 16807 23035
rect 3341 22933 3375 22967
rect 4721 22933 4755 22967
rect 5825 22933 5859 22967
rect 6285 22933 6319 22967
rect 11345 22933 11379 22967
rect 17417 22933 17451 22967
rect 18889 22933 18923 22967
rect 19441 22933 19475 22967
rect 1777 22729 1811 22763
rect 7757 22729 7791 22763
rect 19257 22729 19291 22763
rect 5273 22661 5307 22695
rect 6653 22661 6687 22695
rect 6745 22661 6779 22695
rect 7297 22661 7331 22695
rect 9229 22661 9263 22695
rect 11161 22661 11195 22695
rect 13829 22661 13863 22695
rect 15485 22661 15519 22695
rect 15577 22661 15611 22695
rect 17417 22661 17451 22695
rect 1593 22593 1627 22627
rect 2237 22593 2271 22627
rect 4629 22593 4663 22627
rect 5365 22593 5399 22627
rect 5825 22593 5859 22627
rect 9505 22593 9539 22627
rect 10701 22593 10735 22627
rect 13001 22593 13035 22627
rect 18245 22593 18279 22627
rect 18705 22593 18739 22627
rect 19165 22593 19199 22627
rect 21465 22593 21499 22627
rect 2513 22525 2547 22559
rect 10517 22525 10551 22559
rect 11713 22525 11747 22559
rect 11897 22525 11931 22559
rect 13737 22525 13771 22559
rect 17233 22525 17267 22559
rect 17509 22525 17543 22559
rect 18061 22525 18095 22559
rect 20637 22525 20671 22559
rect 20821 22525 20855 22559
rect 4537 22457 4571 22491
rect 12081 22457 12115 22491
rect 14289 22457 14323 22491
rect 16037 22457 16071 22491
rect 21281 22457 21315 22491
rect 3985 22389 4019 22423
rect 5917 22389 5951 22423
rect 13185 22389 13219 22423
rect 20453 22389 20487 22423
rect 3169 22185 3203 22219
rect 8327 22185 8361 22219
rect 12909 22185 12943 22219
rect 6837 22117 6871 22151
rect 3433 22049 3467 22083
rect 4629 22049 4663 22083
rect 11437 22049 11471 22083
rect 12725 22049 12759 22083
rect 14381 22049 14415 22083
rect 14657 22049 14691 22083
rect 16129 22049 16163 22083
rect 16773 22049 16807 22083
rect 18889 22049 18923 22083
rect 21925 22049 21959 22083
rect 3985 21981 4019 22015
rect 8585 21981 8619 22015
rect 12541 21981 12575 22015
rect 15669 21981 15703 22015
rect 16313 21981 16347 22015
rect 17509 21981 17543 22015
rect 19625 21981 19659 22015
rect 20269 21981 20303 22015
rect 38301 21981 38335 22015
rect 4905 21913 4939 21947
rect 9137 21913 9171 21947
rect 10885 21913 10919 21947
rect 11529 21913 11563 21947
rect 12081 21913 12115 21947
rect 14473 21913 14507 21947
rect 18234 21913 18268 21947
rect 18330 21913 18364 21947
rect 21281 21913 21315 21947
rect 21833 21913 21867 21947
rect 1685 21845 1719 21879
rect 4077 21845 4111 21879
rect 6377 21845 6411 21879
rect 15485 21845 15519 21879
rect 17693 21845 17727 21879
rect 19533 21845 19567 21879
rect 20085 21845 20119 21879
rect 38117 21845 38151 21879
rect 4261 21641 4295 21675
rect 7297 21641 7331 21675
rect 10793 21641 10827 21675
rect 12909 21641 12943 21675
rect 18153 21641 18187 21675
rect 20177 21641 20211 21675
rect 21281 21641 21315 21675
rect 29469 21641 29503 21675
rect 3341 21573 3375 21607
rect 5733 21573 5767 21607
rect 10149 21573 10183 21607
rect 14565 21573 14599 21607
rect 14657 21573 14691 21607
rect 18981 21573 19015 21607
rect 7113 21505 7147 21539
rect 10057 21505 10091 21539
rect 10701 21505 10735 21539
rect 13369 21505 13403 21539
rect 14013 21505 14047 21539
rect 15853 21505 15887 21539
rect 16865 21505 16899 21539
rect 17049 21505 17083 21539
rect 18337 21505 18371 21539
rect 19993 21505 20027 21539
rect 21189 21505 21223 21539
rect 22845 21505 22879 21539
rect 29377 21505 29411 21539
rect 30757 21505 30791 21539
rect 1593 21437 1627 21471
rect 3617 21437 3651 21471
rect 6009 21437 6043 21471
rect 9229 21437 9263 21471
rect 9505 21437 9539 21471
rect 12265 21437 12299 21471
rect 15669 21437 15703 21471
rect 18889 21437 18923 21471
rect 22017 21437 22051 21471
rect 13461 21369 13495 21403
rect 19441 21369 19475 21403
rect 7757 21301 7791 21335
rect 16313 21301 16347 21335
rect 17233 21301 17267 21335
rect 23029 21301 23063 21335
rect 30665 21301 30699 21335
rect 2145 21097 2179 21131
rect 5181 21097 5215 21131
rect 7941 21097 7975 21131
rect 13737 21097 13771 21131
rect 18521 21029 18555 21063
rect 20085 21029 20119 21063
rect 21373 21029 21407 21063
rect 4537 20961 4571 20995
rect 11897 20961 11931 20995
rect 14473 20961 14507 20995
rect 16037 20961 16071 20995
rect 16865 20961 16899 20995
rect 18705 20961 18739 20995
rect 19533 20961 19567 20995
rect 21925 20961 21959 20995
rect 23121 20961 23155 20995
rect 4445 20893 4479 20927
rect 6929 20893 6963 20927
rect 7757 20893 7791 20927
rect 8585 20893 8619 20927
rect 9137 20893 9171 20927
rect 12081 20893 12115 20927
rect 13553 20893 13587 20927
rect 14289 20893 14323 20927
rect 15853 20893 15887 20927
rect 18889 20893 18923 20927
rect 20637 20893 20671 20927
rect 32229 20893 32263 20927
rect 3433 20825 3467 20859
rect 6653 20825 6687 20859
rect 9413 20825 9447 20859
rect 16957 20825 16991 20859
rect 17509 20825 17543 20859
rect 19625 20825 19659 20859
rect 21833 20825 21867 20859
rect 22845 20825 22879 20859
rect 22937 20825 22971 20859
rect 8401 20757 8435 20791
rect 10885 20757 10919 20791
rect 12541 20757 12575 20791
rect 14933 20757 14967 20791
rect 15393 20757 15427 20791
rect 20821 20757 20855 20791
rect 32137 20757 32171 20791
rect 1685 20553 1719 20587
rect 7021 20553 7055 20587
rect 10241 20553 10275 20587
rect 12357 20553 12391 20587
rect 14105 20553 14139 20587
rect 14841 20553 14875 20587
rect 15945 20553 15979 20587
rect 18429 20553 18463 20587
rect 19533 20553 19567 20587
rect 20177 20553 20211 20587
rect 21281 20553 21315 20587
rect 22845 20553 22879 20587
rect 23489 20553 23523 20587
rect 4169 20485 4203 20519
rect 10885 20485 10919 20519
rect 1869 20417 1903 20451
rect 5181 20417 5215 20451
rect 5825 20417 5859 20451
rect 6837 20417 6871 20451
rect 10057 20417 10091 20451
rect 11897 20417 11931 20451
rect 13369 20417 13403 20451
rect 14013 20417 14047 20451
rect 14657 20417 14691 20451
rect 15301 20417 15335 20451
rect 15485 20417 15519 20451
rect 17325 20417 17359 20451
rect 17969 20417 18003 20451
rect 18889 20417 18923 20451
rect 19717 20417 19751 20451
rect 21465 20417 21499 20451
rect 22017 20417 22051 20451
rect 23673 20417 23707 20451
rect 24133 20417 24167 20451
rect 2421 20349 2455 20383
rect 4445 20349 4479 20383
rect 7481 20349 7515 20383
rect 7757 20349 7791 20383
rect 9505 20349 9539 20383
rect 11713 20349 11747 20383
rect 17785 20349 17819 20383
rect 17141 20281 17175 20315
rect 19073 20281 19107 20315
rect 5365 20213 5399 20247
rect 5917 20213 5951 20247
rect 13553 20213 13587 20247
rect 22109 20213 22143 20247
rect 24317 20213 24351 20247
rect 3433 20009 3467 20043
rect 4445 20009 4479 20043
rect 9137 20009 9171 20043
rect 15209 20009 15243 20043
rect 18061 20009 18095 20043
rect 5089 19941 5123 19975
rect 13737 19941 13771 19975
rect 21649 19941 21683 19975
rect 1685 19873 1719 19907
rect 10885 19873 10919 19907
rect 11897 19873 11931 19907
rect 12541 19873 12575 19907
rect 16957 19873 16991 19907
rect 18705 19873 18739 19907
rect 24041 19873 24075 19907
rect 4261 19805 4295 19839
rect 4905 19805 4939 19839
rect 5549 19805 5583 19839
rect 7573 19805 7607 19839
rect 8401 19805 8435 19839
rect 12081 19805 12115 19839
rect 13553 19805 13587 19839
rect 14565 19805 14599 19839
rect 14749 19805 14783 19839
rect 18521 19805 18555 19839
rect 19533 19805 19567 19839
rect 20361 19805 20395 19839
rect 21005 19805 21039 19839
rect 21465 19805 21499 19839
rect 22293 19805 22327 19839
rect 24593 19805 24627 19839
rect 25421 19805 25455 19839
rect 38301 19805 38335 19839
rect 1961 19737 1995 19771
rect 5825 19737 5859 19771
rect 10609 19737 10643 19771
rect 15761 19737 15795 19771
rect 15853 19737 15887 19771
rect 16405 19737 16439 19771
rect 17049 19737 17083 19771
rect 17601 19737 17635 19771
rect 23397 19737 23431 19771
rect 23489 19737 23523 19771
rect 24685 19737 24719 19771
rect 8493 19669 8527 19703
rect 19717 19669 19751 19703
rect 20269 19669 20303 19703
rect 20821 19669 20855 19703
rect 22109 19669 22143 19703
rect 25237 19669 25271 19703
rect 38117 19669 38151 19703
rect 1869 19465 1903 19499
rect 3065 19465 3099 19499
rect 9965 19465 9999 19499
rect 12541 19465 12575 19499
rect 14289 19465 14323 19499
rect 19073 19465 19107 19499
rect 19717 19465 19751 19499
rect 9137 19397 9171 19431
rect 16129 19397 16163 19431
rect 16221 19397 16255 19431
rect 1685 19329 1719 19363
rect 2329 19329 2363 19363
rect 3157 19329 3191 19363
rect 3617 19329 3651 19363
rect 6929 19329 6963 19363
rect 9413 19329 9447 19363
rect 9873 19329 9907 19363
rect 10517 19329 10551 19363
rect 11897 19329 11931 19363
rect 14473 19329 14507 19363
rect 14933 19329 14967 19363
rect 17325 19329 17359 19363
rect 17969 19329 18003 19363
rect 20177 19329 20211 19363
rect 20361 19329 20395 19363
rect 20821 19329 20855 19363
rect 21465 19329 21499 19363
rect 22201 19329 22235 19363
rect 23121 19329 23155 19363
rect 23765 19329 23799 19363
rect 24869 19329 24903 19363
rect 25513 19329 25547 19363
rect 5365 19261 5399 19295
rect 5641 19261 5675 19295
rect 10701 19261 10735 19295
rect 12081 19261 12115 19295
rect 13461 19261 13495 19295
rect 13645 19261 13679 19295
rect 15577 19261 15611 19295
rect 17785 19261 17819 19295
rect 18429 19261 18463 19295
rect 18613 19261 18647 19295
rect 21281 19261 21315 19295
rect 23581 19261 23615 19295
rect 24685 19261 24719 19295
rect 15117 19193 15151 19227
rect 2513 19125 2547 19159
rect 7113 19125 7147 19159
rect 7665 19125 7699 19159
rect 11069 19125 11103 19159
rect 13001 19125 13035 19159
rect 22017 19125 22051 19159
rect 24501 19125 24535 19159
rect 25329 19125 25363 19159
rect 5076 18921 5110 18955
rect 8585 18921 8619 18955
rect 13001 18921 13035 18955
rect 14657 18921 14691 18955
rect 19441 18921 19475 18955
rect 20913 18921 20947 18955
rect 21373 18921 21407 18955
rect 25789 18921 25823 18955
rect 31033 18921 31067 18955
rect 6561 18853 6595 18887
rect 9137 18853 9171 18887
rect 18245 18853 18279 18887
rect 26433 18853 26467 18887
rect 3433 18785 3467 18819
rect 4813 18785 4847 18819
rect 8125 18785 8159 18819
rect 13185 18785 13219 18819
rect 15577 18785 15611 18819
rect 17233 18785 17267 18819
rect 18705 18785 18739 18819
rect 19901 18785 19935 18819
rect 22109 18785 22143 18819
rect 24041 18785 24075 18819
rect 24685 18785 24719 18819
rect 25329 18785 25363 18819
rect 4353 18717 4387 18751
rect 7113 18717 7147 18751
rect 7941 18717 7975 18751
rect 10885 18717 10919 18751
rect 11621 18717 11655 18751
rect 11805 18717 11839 18751
rect 13369 18717 13403 18751
rect 14841 18717 14875 18751
rect 18889 18717 18923 18751
rect 20085 18717 20119 18751
rect 20729 18717 20763 18751
rect 21557 18717 21591 18751
rect 22017 18717 22051 18751
rect 25973 18717 26007 18751
rect 26617 18717 26651 18751
rect 31125 18717 31159 18751
rect 38301 18717 38335 18751
rect 3157 18649 3191 18683
rect 10609 18649 10643 18683
rect 15853 18649 15887 18683
rect 15945 18649 15979 18683
rect 16589 18649 16623 18683
rect 16681 18649 16715 18683
rect 23397 18649 23431 18683
rect 23489 18649 23523 18683
rect 24777 18649 24811 18683
rect 1685 18581 1719 18615
rect 4261 18581 4295 18615
rect 7205 18581 7239 18615
rect 12265 18581 12299 18615
rect 22661 18581 22695 18615
rect 38117 18581 38151 18615
rect 3985 18377 4019 18411
rect 8861 18377 8895 18411
rect 12357 18377 12391 18411
rect 14565 18377 14599 18411
rect 16313 18377 16347 18411
rect 17509 18377 17543 18411
rect 19533 18377 19567 18411
rect 22661 18377 22695 18411
rect 24317 18377 24351 18411
rect 26157 18377 26191 18411
rect 13369 18309 13403 18343
rect 13461 18309 13495 18343
rect 18337 18309 18371 18343
rect 5733 18241 5767 18275
rect 8401 18241 8435 18275
rect 10609 18241 10643 18275
rect 11897 18241 11931 18275
rect 15025 18241 15059 18275
rect 19993 18241 20027 18275
rect 21281 18241 21315 18275
rect 21465 18241 21499 18275
rect 23673 18241 23707 18275
rect 24961 18241 24995 18275
rect 25605 18241 25639 18275
rect 26249 18241 26283 18275
rect 34345 18241 34379 18275
rect 1685 18173 1719 18207
rect 1961 18173 1995 18207
rect 5457 18173 5491 18207
rect 6653 18173 6687 18207
rect 8125 18173 8159 18207
rect 10333 18173 10367 18207
rect 11713 18173 11747 18207
rect 15669 18173 15703 18207
rect 15853 18173 15887 18207
rect 16865 18173 16899 18207
rect 17049 18173 17083 18207
rect 18245 18173 18279 18207
rect 18521 18173 18555 18207
rect 20177 18173 20211 18207
rect 22017 18173 22051 18207
rect 22201 18173 22235 18207
rect 23857 18173 23891 18207
rect 25513 18173 25547 18207
rect 12909 18105 12943 18139
rect 3433 18037 3467 18071
rect 15117 18037 15151 18071
rect 20821 18037 20855 18071
rect 24777 18037 24811 18071
rect 34253 18037 34287 18071
rect 1593 17833 1627 17867
rect 4077 17833 4111 17867
rect 8585 17833 8619 17867
rect 17509 17833 17543 17867
rect 22293 17833 22327 17867
rect 23121 17833 23155 17867
rect 24777 17833 24811 17867
rect 25421 17833 25455 17867
rect 9137 17765 9171 17799
rect 14289 17765 14323 17799
rect 16037 17765 16071 17799
rect 3341 17697 3375 17731
rect 6653 17697 6687 17731
rect 11437 17697 11471 17731
rect 15485 17697 15519 17731
rect 16773 17697 16807 17731
rect 18429 17697 18463 17731
rect 18613 17697 18647 17731
rect 21189 17697 21223 17731
rect 22477 17697 22511 17731
rect 3985 17629 4019 17663
rect 7297 17629 7331 17663
rect 7941 17629 7975 17663
rect 8409 17629 8443 17663
rect 10885 17629 10919 17663
rect 14749 17629 14783 17663
rect 14933 17629 14967 17663
rect 16681 17629 16715 17663
rect 17325 17629 17359 17663
rect 19809 17629 19843 17663
rect 22661 17629 22695 17663
rect 23581 17629 23615 17663
rect 23765 17629 23799 17663
rect 24593 17629 24627 17663
rect 25237 17629 25271 17663
rect 29745 17629 29779 17663
rect 3065 17561 3099 17595
rect 4629 17561 4663 17595
rect 6377 17561 6411 17595
rect 10609 17561 10643 17595
rect 11529 17561 11563 17595
rect 12081 17561 12115 17595
rect 13001 17561 13035 17595
rect 13553 17561 13587 17595
rect 13645 17561 13679 17595
rect 15577 17561 15611 17595
rect 20545 17561 20579 17595
rect 20637 17561 20671 17595
rect 7113 17493 7147 17527
rect 7757 17493 7791 17527
rect 17969 17493 18003 17527
rect 19901 17493 19935 17527
rect 25881 17493 25915 17527
rect 29837 17493 29871 17527
rect 22201 17289 22235 17323
rect 22661 17289 22695 17323
rect 33977 17289 34011 17323
rect 2145 17221 2179 17255
rect 9965 17221 9999 17255
rect 10057 17221 10091 17255
rect 11989 17221 12023 17255
rect 20821 17221 20855 17255
rect 25145 17221 25179 17255
rect 4169 17153 4203 17187
rect 5181 17153 5215 17187
rect 5825 17153 5859 17187
rect 6745 17153 6779 17187
rect 11713 17153 11747 17187
rect 14105 17153 14139 17187
rect 15485 17153 15519 17187
rect 16129 17153 16163 17187
rect 17233 17153 17267 17187
rect 17877 17153 17911 17187
rect 18061 17153 18095 17187
rect 20269 17153 20303 17187
rect 21281 17153 21315 17187
rect 22017 17153 22051 17187
rect 26157 17153 26191 17187
rect 27353 17153 27387 17187
rect 33793 17153 33827 17187
rect 38025 17153 38059 17187
rect 3893 17085 3927 17119
rect 7389 17085 7423 17119
rect 7665 17085 7699 17119
rect 13461 17085 13495 17119
rect 13921 17085 13955 17119
rect 18981 17085 19015 17119
rect 19165 17085 19199 17119
rect 21465 17085 21499 17119
rect 24317 17085 24351 17119
rect 24501 17085 24535 17119
rect 25053 17085 25087 17119
rect 25329 17085 25363 17119
rect 10517 17017 10551 17051
rect 14289 17017 14323 17051
rect 16313 17017 16347 17051
rect 17417 17017 17451 17051
rect 18245 17017 18279 17051
rect 19349 17017 19383 17051
rect 20085 17017 20119 17051
rect 38209 17017 38243 17051
rect 5365 16949 5399 16983
rect 6009 16949 6043 16983
rect 6929 16949 6963 16983
rect 9137 16949 9171 16983
rect 15669 16949 15703 16983
rect 24133 16949 24167 16983
rect 26249 16949 26283 16983
rect 27169 16949 27203 16983
rect 4432 16745 4466 16779
rect 16313 16745 16347 16779
rect 17141 16745 17175 16779
rect 23489 16745 23523 16779
rect 24593 16745 24627 16779
rect 25697 16745 25731 16779
rect 1685 16609 1719 16643
rect 1961 16609 1995 16643
rect 4169 16609 4203 16643
rect 9137 16609 9171 16643
rect 10609 16609 10643 16643
rect 10885 16609 10919 16643
rect 11345 16609 11379 16643
rect 18061 16609 18095 16643
rect 18245 16609 18279 16643
rect 19993 16609 20027 16643
rect 20177 16609 20211 16643
rect 22753 16609 22787 16643
rect 22937 16609 22971 16643
rect 25237 16609 25271 16643
rect 6837 16541 6871 16575
rect 13553 16541 13587 16575
rect 14473 16541 14507 16575
rect 14565 16541 14599 16575
rect 15853 16541 15887 16575
rect 16497 16541 16531 16575
rect 16957 16541 16991 16575
rect 18797 16541 18831 16575
rect 18889 16541 18923 16575
rect 21465 16541 21499 16575
rect 21557 16541 21591 16575
rect 23397 16541 23431 16575
rect 25053 16541 25087 16575
rect 25881 16541 25915 16575
rect 34989 16541 35023 16575
rect 35081 16541 35115 16575
rect 6193 16473 6227 16507
rect 11621 16473 11655 16507
rect 15209 16473 15243 16507
rect 15301 16473 15335 16507
rect 17601 16473 17635 16507
rect 3433 16405 3467 16439
rect 8125 16405 8159 16439
rect 13093 16405 13127 16439
rect 13737 16405 13771 16439
rect 20637 16405 20671 16439
rect 22293 16405 22327 16439
rect 1685 16201 1719 16235
rect 13001 16201 13035 16235
rect 22661 16201 22695 16235
rect 23121 16201 23155 16235
rect 23765 16201 23799 16235
rect 25053 16201 25087 16235
rect 10149 16133 10183 16167
rect 10241 16133 10275 16167
rect 11161 16133 11195 16167
rect 16129 16133 16163 16167
rect 19993 16133 20027 16167
rect 20821 16133 20855 16167
rect 20913 16133 20947 16167
rect 1869 16065 1903 16099
rect 6009 16065 6043 16099
rect 6745 16065 6779 16099
rect 11713 16065 11747 16099
rect 17141 16065 17175 16099
rect 17233 16065 17267 16099
rect 19533 16065 19567 16099
rect 23305 16065 23339 16099
rect 23949 16065 23983 16099
rect 24593 16065 24627 16099
rect 25237 16065 25271 16099
rect 25881 16065 25915 16099
rect 2881 15997 2915 16031
rect 3157 15997 3191 16031
rect 4905 15997 4939 16031
rect 7481 15997 7515 16031
rect 7757 15997 7791 16031
rect 13921 15997 13955 16031
rect 14105 15997 14139 16031
rect 15945 15997 15979 16031
rect 16221 15997 16255 16031
rect 17785 15997 17819 16031
rect 17969 15997 18003 16031
rect 19349 15997 19383 16031
rect 22017 15997 22051 16031
rect 22201 15997 22235 16031
rect 6929 15929 6963 15963
rect 18153 15929 18187 15963
rect 21373 15929 21407 15963
rect 24409 15929 24443 15963
rect 25697 15929 25731 15963
rect 5825 15861 5859 15895
rect 9229 15861 9263 15895
rect 14289 15861 14323 15895
rect 3341 15657 3375 15691
rect 8585 15657 8619 15691
rect 13645 15657 13679 15691
rect 14565 15657 14599 15691
rect 16957 15657 16991 15691
rect 20085 15657 20119 15691
rect 24685 15657 24719 15691
rect 38117 15657 38151 15691
rect 4077 15589 4111 15623
rect 1593 15521 1627 15555
rect 5273 15521 5307 15555
rect 12357 15521 12391 15555
rect 13001 15521 13035 15555
rect 15761 15521 15795 15555
rect 18889 15521 18923 15555
rect 21189 15521 21223 15555
rect 21465 15521 21499 15555
rect 23121 15521 23155 15555
rect 4169 15453 4203 15487
rect 4629 15453 4663 15487
rect 7941 15453 7975 15487
rect 8125 15453 8159 15487
rect 9137 15453 9171 15487
rect 13185 15453 13219 15487
rect 14381 15453 14415 15487
rect 16773 15453 16807 15487
rect 20269 15453 20303 15487
rect 20453 15453 20487 15487
rect 24041 15453 24075 15487
rect 24593 15453 24627 15487
rect 38301 15453 38335 15487
rect 1869 15385 1903 15419
rect 5549 15385 5583 15419
rect 7297 15385 7331 15419
rect 9413 15385 9447 15419
rect 11713 15385 11747 15419
rect 12265 15385 12299 15419
rect 15117 15385 15151 15419
rect 15209 15385 15243 15419
rect 17417 15385 17451 15419
rect 17969 15385 18003 15419
rect 18061 15385 18095 15419
rect 21281 15385 21315 15419
rect 22753 15385 22787 15419
rect 22845 15385 22879 15419
rect 4813 15317 4847 15351
rect 10885 15317 10919 15351
rect 23857 15317 23891 15351
rect 1777 15113 1811 15147
rect 17233 15113 17267 15147
rect 19717 15113 19751 15147
rect 22017 15113 22051 15147
rect 3893 15045 3927 15079
rect 9137 15045 9171 15079
rect 12265 15045 12299 15079
rect 12357 15045 12391 15079
rect 15669 15045 15703 15079
rect 15761 15045 15795 15079
rect 17969 15045 18003 15079
rect 23305 15045 23339 15079
rect 1685 14977 1719 15011
rect 2329 14977 2363 15011
rect 2973 14977 3007 15011
rect 3617 14977 3651 15011
rect 6561 14977 6595 15011
rect 17141 14977 17175 15011
rect 20637 14977 20671 15011
rect 21281 14977 21315 15011
rect 22201 14977 22235 15011
rect 24133 14977 24167 15011
rect 24777 14977 24811 15011
rect 29193 14977 29227 15011
rect 5641 14909 5675 14943
rect 6837 14909 6871 14943
rect 8861 14909 8895 14943
rect 12909 14909 12943 14943
rect 13093 14909 13127 14943
rect 14473 14909 14507 14943
rect 14657 14909 14691 14943
rect 17877 14909 17911 14943
rect 19073 14909 19107 14943
rect 19257 14909 19291 14943
rect 20821 14909 20855 14943
rect 23121 14909 23155 14943
rect 23397 14909 23431 14943
rect 24685 14909 24719 14943
rect 3157 14841 3191 14875
rect 11805 14841 11839 14875
rect 16221 14841 16255 14875
rect 18429 14841 18463 14875
rect 2421 14773 2455 14807
rect 8309 14773 8343 14807
rect 10609 14773 10643 14807
rect 13553 14773 13587 14807
rect 15117 14773 15151 14807
rect 20177 14773 20211 14807
rect 21465 14773 21499 14807
rect 23949 14773 23983 14807
rect 29285 14773 29319 14807
rect 4721 14569 4755 14603
rect 10885 14569 10919 14603
rect 16129 14569 16163 14603
rect 18705 14569 18739 14603
rect 19533 14569 19567 14603
rect 20361 14569 20395 14603
rect 21373 14569 21407 14603
rect 24593 14569 24627 14603
rect 25237 14569 25271 14603
rect 13737 14501 13771 14535
rect 15485 14501 15519 14535
rect 1685 14433 1719 14467
rect 4077 14433 4111 14467
rect 7665 14433 7699 14467
rect 9137 14433 9171 14467
rect 11805 14433 11839 14467
rect 12173 14433 12207 14467
rect 33609 14433 33643 14467
rect 4169 14365 4203 14399
rect 4813 14365 4847 14399
rect 8401 14365 8435 14399
rect 13093 14365 13127 14399
rect 13277 14365 13311 14399
rect 15669 14365 15703 14399
rect 16589 14365 16623 14399
rect 16773 14365 16807 14399
rect 18889 14365 18923 14399
rect 19441 14365 19475 14399
rect 20545 14365 20579 14399
rect 20729 14365 20763 14399
rect 21465 14365 21499 14399
rect 22477 14365 22511 14399
rect 22661 14365 22695 14399
rect 23305 14365 23339 14399
rect 23765 14365 23799 14399
rect 24777 14365 24811 14399
rect 25421 14365 25455 14399
rect 33701 14365 33735 14399
rect 3433 14297 3467 14331
rect 5641 14297 5675 14331
rect 7389 14297 7423 14331
rect 9413 14297 9447 14331
rect 11897 14297 11931 14331
rect 14381 14297 14415 14331
rect 14473 14297 14507 14331
rect 15025 14297 15059 14331
rect 17509 14297 17543 14331
rect 18061 14297 18095 14331
rect 18153 14297 18187 14331
rect 23857 14297 23891 14331
rect 8585 14229 8619 14263
rect 22017 14229 22051 14263
rect 6837 14025 6871 14059
rect 13645 14025 13679 14059
rect 16037 14025 16071 14059
rect 16865 14025 16899 14059
rect 17969 14025 18003 14059
rect 18613 14025 18647 14059
rect 19993 14025 20027 14059
rect 21465 14025 21499 14059
rect 35081 14025 35115 14059
rect 3617 13957 3651 13991
rect 4353 13957 4387 13991
rect 9321 13957 9355 13991
rect 11897 13957 11931 13991
rect 14933 13957 14967 13991
rect 15485 13957 15519 13991
rect 22661 13957 22695 13991
rect 4077 13889 4111 13923
rect 8585 13889 8619 13923
rect 9045 13889 9079 13923
rect 13001 13889 13035 13923
rect 15945 13889 15979 13923
rect 18429 13889 18463 13923
rect 19349 13889 19383 13923
rect 20821 13889 20855 13923
rect 23489 13889 23523 13923
rect 34897 13889 34931 13923
rect 38025 13889 38059 13923
rect 1593 13821 1627 13855
rect 11805 13821 11839 13855
rect 12081 13821 12115 13855
rect 14105 13821 14139 13855
rect 14289 13821 14323 13855
rect 14841 13821 14875 13855
rect 19533 13821 19567 13855
rect 21005 13821 21039 13855
rect 22477 13821 22511 13855
rect 22753 13821 22787 13855
rect 23949 13821 23983 13855
rect 5825 13753 5859 13787
rect 10793 13753 10827 13787
rect 1850 13685 1884 13719
rect 8327 13685 8361 13719
rect 13185 13685 13219 13719
rect 23305 13685 23339 13719
rect 38209 13685 38243 13719
rect 7941 13481 7975 13515
rect 10885 13481 10919 13515
rect 21189 13481 21223 13515
rect 23489 13481 23523 13515
rect 30665 13481 30699 13515
rect 8493 13413 8527 13447
rect 13645 13413 13679 13447
rect 1593 13345 1627 13379
rect 3341 13345 3375 13379
rect 4997 13345 5031 13379
rect 9137 13345 9171 13379
rect 11345 13345 11379 13379
rect 11989 13345 12023 13379
rect 14565 13345 14599 13379
rect 16313 13345 16347 13379
rect 16773 13345 16807 13379
rect 17693 13345 17727 13379
rect 21649 13345 21683 13379
rect 22385 13345 22419 13379
rect 22661 13345 22695 13379
rect 4261 13277 4295 13311
rect 7297 13277 7331 13311
rect 7757 13277 7791 13311
rect 8401 13277 8435 13311
rect 11529 13277 11563 13311
rect 16129 13277 16163 13311
rect 17877 13277 17911 13311
rect 19901 13277 19935 13311
rect 20085 13277 20119 13311
rect 21005 13277 21039 13311
rect 23673 13277 23707 13311
rect 30757 13277 30791 13311
rect 1869 13209 1903 13243
rect 7021 13209 7055 13243
rect 9413 13209 9447 13243
rect 13093 13209 13127 13243
rect 13185 13209 13219 13243
rect 14657 13209 14691 13243
rect 15209 13209 15243 13243
rect 22477 13209 22511 13243
rect 4077 13141 4111 13175
rect 5549 13141 5583 13175
rect 18337 13141 18371 13175
rect 20545 13141 20579 13175
rect 7297 12937 7331 12971
rect 9137 12937 9171 12971
rect 10701 12937 10735 12971
rect 14841 12937 14875 12971
rect 22017 12937 22051 12971
rect 22661 12937 22695 12971
rect 24041 12937 24075 12971
rect 3341 12869 3375 12903
rect 5641 12869 5675 12903
rect 7849 12869 7883 12903
rect 15577 12869 15611 12903
rect 16129 12869 16163 12903
rect 18337 12869 18371 12903
rect 19533 12869 19567 12903
rect 20913 12869 20947 12903
rect 3617 12801 3651 12835
rect 6561 12801 6595 12835
rect 7205 12801 7239 12835
rect 10057 12801 10091 12835
rect 12081 12801 12115 12835
rect 14105 12801 14139 12835
rect 14749 12801 14783 12835
rect 22201 12801 22235 12835
rect 22845 12801 22879 12835
rect 23489 12801 23523 12835
rect 23949 12801 23983 12835
rect 29653 12801 29687 12835
rect 1593 12733 1627 12767
rect 5917 12733 5951 12767
rect 10241 12733 10275 12767
rect 12541 12733 12575 12767
rect 12725 12733 12759 12767
rect 15485 12733 15519 12767
rect 17509 12733 17543 12767
rect 17693 12733 17727 12767
rect 18245 12733 18279 12767
rect 19441 12733 19475 12767
rect 20821 12733 20855 12767
rect 21465 12733 21499 12767
rect 6745 12665 6779 12699
rect 11897 12665 11931 12699
rect 12909 12665 12943 12699
rect 14289 12665 14323 12699
rect 17325 12665 17359 12699
rect 18797 12665 18831 12699
rect 19993 12665 20027 12699
rect 23305 12665 23339 12699
rect 4169 12597 4203 12631
rect 29745 12597 29779 12631
rect 3175 12393 3209 12427
rect 6561 12393 6595 12427
rect 13553 12393 13587 12427
rect 15485 12393 15519 12427
rect 16313 12393 16347 12427
rect 17509 12393 17543 12427
rect 18337 12393 18371 12427
rect 19625 12393 19659 12427
rect 20729 12393 20763 12427
rect 21557 12393 21591 12427
rect 12817 12325 12851 12359
rect 14473 12325 14507 12359
rect 23489 12325 23523 12359
rect 3433 12257 3467 12291
rect 3985 12257 4019 12291
rect 8033 12257 8067 12291
rect 10885 12257 10919 12291
rect 11345 12257 11379 12291
rect 11989 12257 12023 12291
rect 14933 12257 14967 12291
rect 8309 12189 8343 12223
rect 11529 12189 11563 12223
rect 12449 12189 12483 12223
rect 12633 12189 12667 12223
rect 13737 12189 13771 12223
rect 14289 12189 14323 12223
rect 15117 12189 15151 12223
rect 16497 12189 16531 12223
rect 16681 12189 16715 12223
rect 17141 12189 17175 12223
rect 17325 12189 17359 12223
rect 18705 12189 18739 12223
rect 18889 12189 18923 12223
rect 19717 12189 19751 12223
rect 20361 12189 20395 12223
rect 20545 12189 20579 12223
rect 21649 12189 21683 12223
rect 4261 12121 4295 12155
rect 6009 12121 6043 12155
rect 10609 12121 10643 12155
rect 22385 12121 22419 12155
rect 22937 12121 22971 12155
rect 23029 12121 23063 12155
rect 1685 12053 1719 12087
rect 9137 12053 9171 12087
rect 5917 11849 5951 11883
rect 6837 11849 6871 11883
rect 12357 11849 12391 11883
rect 14473 11849 14507 11883
rect 15669 11849 15703 11883
rect 16313 11849 16347 11883
rect 17969 11849 18003 11883
rect 18613 11849 18647 11883
rect 19717 11849 19751 11883
rect 20453 11849 20487 11883
rect 21097 11849 21131 11883
rect 23397 11849 23431 11883
rect 38117 11849 38151 11883
rect 2329 11781 2363 11815
rect 8861 11781 8895 11815
rect 17417 11781 17451 11815
rect 4813 11713 4847 11747
rect 5825 11713 5859 11747
rect 6745 11713 6779 11747
rect 9137 11713 9171 11747
rect 10609 11713 10643 11747
rect 11897 11713 11931 11747
rect 12817 11713 12851 11747
rect 13645 11713 13679 11747
rect 17325 11713 17359 11747
rect 18797 11713 18831 11747
rect 19625 11713 19659 11747
rect 20269 11713 20303 11747
rect 21189 11713 21223 11747
rect 22109 11713 22143 11747
rect 22753 11713 22787 11747
rect 23581 11713 23615 11747
rect 27445 11713 27479 11747
rect 34161 11713 34195 11747
rect 38301 11713 38335 11747
rect 2053 11645 2087 11679
rect 4077 11645 4111 11679
rect 10425 11645 10459 11679
rect 11713 11645 11747 11679
rect 15025 11645 15059 11679
rect 15209 11645 15243 11679
rect 4905 11577 4939 11611
rect 12909 11577 12943 11611
rect 22293 11577 22327 11611
rect 22937 11577 22971 11611
rect 7389 11509 7423 11543
rect 10793 11509 10827 11543
rect 13829 11509 13863 11543
rect 27537 11509 27571 11543
rect 34345 11509 34379 11543
rect 1685 11305 1719 11339
rect 4261 11305 4295 11339
rect 9781 11305 9815 11339
rect 10977 11305 11011 11339
rect 11805 11305 11839 11339
rect 13185 11305 13219 11339
rect 14565 11305 14599 11339
rect 15485 11305 15519 11339
rect 16681 11305 16715 11339
rect 17877 11305 17911 11339
rect 18705 11305 18739 11339
rect 19625 11305 19659 11339
rect 20453 11305 20487 11339
rect 12449 11237 12483 11271
rect 17325 11237 17359 11271
rect 6009 11169 6043 11203
rect 6837 11169 6871 11203
rect 8309 11169 8343 11203
rect 3433 11101 3467 11135
rect 8585 11101 8619 11135
rect 9689 11101 9723 11135
rect 10333 11101 10367 11135
rect 10517 11101 10551 11135
rect 11897 11101 11931 11135
rect 12357 11101 12391 11135
rect 13001 11101 13035 11135
rect 14381 11101 14415 11135
rect 15393 11101 15427 11135
rect 16773 11101 16807 11135
rect 17233 11101 17267 11135
rect 18061 11101 18095 11135
rect 18521 11101 18555 11135
rect 19809 11101 19843 11135
rect 20269 11101 20303 11135
rect 3157 11033 3191 11067
rect 5733 11033 5767 11067
rect 3433 10761 3467 10795
rect 6653 10761 6687 10795
rect 7665 10761 7699 10795
rect 10149 10761 10183 10795
rect 12817 10761 12851 10795
rect 13553 10761 13587 10795
rect 14841 10761 14875 10795
rect 15669 10761 15703 10795
rect 16313 10761 16347 10795
rect 17325 10761 17359 10795
rect 18061 10761 18095 10795
rect 18889 10761 18923 10795
rect 19717 10761 19751 10795
rect 1961 10693 1995 10727
rect 5733 10693 5767 10727
rect 9137 10693 9171 10727
rect 10701 10693 10735 10727
rect 1685 10625 1719 10659
rect 6009 10625 6043 10659
rect 6561 10625 6595 10659
rect 9413 10625 9447 10659
rect 9965 10625 9999 10659
rect 10609 10625 10643 10659
rect 11989 10625 12023 10659
rect 12633 10625 12667 10659
rect 13461 10625 13495 10659
rect 14289 10625 14323 10659
rect 14933 10625 14967 10659
rect 16129 10625 16163 10659
rect 17233 10625 17267 10659
rect 17877 10625 17911 10659
rect 19533 10625 19567 10659
rect 20361 10625 20395 10659
rect 30021 10625 30055 10659
rect 38025 10625 38059 10659
rect 14105 10489 14139 10523
rect 4261 10421 4295 10455
rect 12173 10421 12207 10455
rect 20177 10421 20211 10455
rect 30113 10421 30147 10455
rect 38209 10421 38243 10455
rect 6837 10217 6871 10251
rect 8321 10217 8355 10251
rect 10517 10217 10551 10251
rect 11345 10217 11379 10251
rect 11989 10217 12023 10251
rect 13093 10217 13127 10251
rect 14749 10217 14783 10251
rect 15761 10217 15795 10251
rect 16405 10217 16439 10251
rect 17233 10217 17267 10251
rect 17969 10217 18003 10251
rect 18705 10217 18739 10251
rect 19533 10217 19567 10251
rect 25329 10217 25363 10251
rect 4077 10149 4111 10183
rect 6377 10149 6411 10183
rect 9321 10149 9355 10183
rect 20177 10149 20211 10183
rect 4629 10081 4663 10115
rect 8585 10081 8619 10115
rect 12541 10081 12575 10115
rect 3985 10013 4019 10047
rect 9229 10013 9263 10047
rect 10057 10013 10091 10047
rect 10701 10013 10735 10047
rect 11161 10013 11195 10047
rect 11805 10013 11839 10047
rect 12633 10013 12667 10047
rect 13277 10013 13311 10047
rect 14933 10013 14967 10047
rect 15577 10013 15611 10047
rect 16221 10013 16255 10047
rect 17417 10013 17451 10047
rect 18061 10013 18095 10047
rect 18889 10013 18923 10047
rect 19441 10013 19475 10047
rect 20269 10013 20303 10047
rect 24593 10013 24627 10047
rect 25421 10013 25455 10047
rect 34897 10013 34931 10047
rect 3433 9945 3467 9979
rect 4905 9945 4939 9979
rect 24685 9945 24719 9979
rect 2145 9877 2179 9911
rect 9873 9877 9907 9911
rect 35081 9877 35115 9911
rect 8309 9673 8343 9707
rect 12449 9673 12483 9707
rect 14841 9673 14875 9707
rect 16865 9673 16899 9707
rect 17693 9673 17727 9707
rect 2789 9605 2823 9639
rect 4353 9605 4387 9639
rect 7297 9605 7331 9639
rect 9597 9605 9631 9639
rect 10609 9605 10643 9639
rect 11161 9605 11195 9639
rect 13645 9605 13679 9639
rect 16221 9605 16255 9639
rect 1685 9537 1719 9571
rect 4813 9537 4847 9571
rect 5825 9537 5859 9571
rect 6561 9537 6595 9571
rect 7389 9537 7423 9571
rect 12909 9537 12943 9571
rect 13553 9537 13587 9571
rect 14197 9537 14231 9571
rect 14289 9537 14323 9571
rect 15025 9537 15059 9571
rect 15669 9537 15703 9571
rect 16313 9537 16347 9571
rect 17049 9537 17083 9571
rect 17877 9537 17911 9571
rect 34713 9537 34747 9571
rect 1777 9469 1811 9503
rect 5917 9469 5951 9503
rect 6653 9469 6687 9503
rect 10517 9469 10551 9503
rect 13093 9401 13127 9435
rect 15485 9401 15519 9435
rect 4905 9333 4939 9367
rect 34621 9333 34655 9367
rect 1685 9129 1719 9163
rect 3175 9129 3209 9163
rect 5089 9129 5123 9163
rect 5733 9129 5767 9163
rect 8493 9129 8527 9163
rect 9781 9129 9815 9163
rect 11345 9129 11379 9163
rect 12081 9129 12115 9163
rect 12817 9129 12851 9163
rect 13553 9129 13587 9163
rect 14473 9129 14507 9163
rect 15669 9129 15703 9163
rect 4077 9061 4111 9095
rect 3433 8993 3467 9027
rect 7481 8993 7515 9027
rect 15025 8993 15059 9027
rect 3985 8925 4019 8959
rect 5181 8925 5215 8959
rect 8401 8925 8435 8959
rect 9689 8925 9723 8959
rect 11253 8925 11287 8959
rect 11897 8925 11931 8959
rect 12633 8925 12667 8959
rect 13737 8925 13771 8959
rect 14381 8925 14415 8959
rect 15853 8925 15887 8959
rect 16497 8925 16531 8959
rect 18613 8925 18647 8959
rect 25145 8925 25179 8959
rect 30849 8925 30883 8959
rect 38025 8925 38059 8959
rect 7205 8857 7239 8891
rect 10333 8789 10367 8823
rect 16313 8789 16347 8823
rect 18705 8789 18739 8823
rect 25237 8789 25271 8823
rect 30941 8789 30975 8823
rect 38209 8789 38243 8823
rect 6653 8585 6687 8619
rect 7205 8585 7239 8619
rect 7941 8585 7975 8619
rect 8677 8585 8711 8619
rect 9413 8585 9447 8619
rect 10425 8585 10459 8619
rect 11805 8585 11839 8619
rect 12633 8585 12667 8619
rect 14749 8585 14783 8619
rect 15301 8585 15335 8619
rect 1961 8517 1995 8551
rect 6009 8449 6043 8483
rect 6745 8449 6779 8483
rect 7389 8449 7423 8483
rect 7849 8449 7883 8483
rect 8585 8449 8619 8483
rect 9229 8449 9263 8483
rect 10333 8449 10367 8483
rect 11161 8449 11195 8483
rect 11713 8449 11747 8483
rect 12817 8449 12851 8483
rect 14657 8449 14691 8483
rect 15485 8449 15519 8483
rect 16037 8449 16071 8483
rect 16865 8449 16899 8483
rect 1685 8381 1719 8415
rect 3433 8381 3467 8415
rect 5733 8381 5767 8415
rect 10977 8313 11011 8347
rect 16129 8313 16163 8347
rect 16957 8313 16991 8347
rect 4261 8245 4295 8279
rect 6837 8041 6871 8075
rect 9873 8041 9907 8075
rect 3433 7973 3467 8007
rect 1685 7905 1719 7939
rect 5089 7905 5123 7939
rect 5365 7905 5399 7939
rect 7389 7905 7423 7939
rect 4353 7837 4387 7871
rect 7297 7837 7331 7871
rect 8585 7837 8619 7871
rect 9689 7837 9723 7871
rect 11621 7837 11655 7871
rect 35357 7837 35391 7871
rect 1961 7769 1995 7803
rect 4445 7769 4479 7803
rect 8493 7701 8527 7735
rect 11437 7701 11471 7735
rect 35541 7701 35575 7735
rect 1685 7497 1719 7531
rect 3065 7497 3099 7531
rect 3709 7497 3743 7531
rect 6653 7497 6687 7531
rect 9229 7497 9263 7531
rect 24593 7497 24627 7531
rect 38117 7497 38151 7531
rect 1869 7361 1903 7395
rect 2329 7361 2363 7395
rect 3157 7361 3191 7395
rect 3617 7361 3651 7395
rect 4261 7361 4295 7395
rect 6561 7361 6595 7395
rect 9137 7361 9171 7395
rect 24685 7361 24719 7395
rect 34437 7361 34471 7395
rect 38301 7361 38335 7395
rect 2421 7293 2455 7327
rect 4537 7293 4571 7327
rect 6009 7225 6043 7259
rect 34345 7225 34379 7259
rect 5917 6953 5951 6987
rect 4629 6885 4663 6919
rect 2697 6817 2731 6851
rect 5273 6817 5307 6851
rect 9689 6817 9723 6851
rect 14381 6817 14415 6851
rect 21281 6817 21315 6851
rect 35173 6817 35207 6851
rect 1961 6749 1995 6783
rect 2605 6749 2639 6783
rect 3249 6749 3283 6783
rect 3341 6749 3375 6783
rect 4545 6751 4579 6785
rect 5181 6749 5215 6783
rect 6009 6749 6043 6783
rect 6469 6749 6503 6783
rect 14289 6749 14323 6783
rect 21373 6749 21407 6783
rect 29929 6749 29963 6783
rect 30757 6749 30791 6783
rect 35265 6749 35299 6783
rect 2053 6681 2087 6715
rect 9229 6681 9263 6715
rect 9321 6681 9355 6715
rect 30665 6681 30699 6715
rect 6561 6613 6595 6647
rect 29837 6613 29871 6647
rect 2697 6409 2731 6443
rect 3341 6409 3375 6443
rect 4077 6409 4111 6443
rect 4721 6409 4755 6443
rect 5365 6409 5399 6443
rect 8861 6409 8895 6443
rect 1593 6273 1627 6307
rect 2605 6273 2639 6307
rect 3433 6273 3467 6307
rect 4169 6273 4203 6307
rect 4629 6273 4663 6307
rect 5273 6273 5307 6307
rect 6745 6273 6779 6307
rect 8033 6273 8067 6307
rect 8677 6273 8711 6307
rect 28181 6273 28215 6307
rect 8125 6205 8159 6239
rect 1777 6137 1811 6171
rect 6653 6069 6687 6103
rect 28089 6069 28123 6103
rect 2697 5865 2731 5899
rect 4445 5865 4479 5899
rect 8585 5865 8619 5899
rect 9965 5865 9999 5899
rect 15577 5865 15611 5899
rect 3341 5797 3375 5831
rect 6837 5797 6871 5831
rect 6285 5729 6319 5763
rect 1593 5661 1627 5695
rect 2605 5661 2639 5695
rect 3249 5661 3283 5695
rect 4353 5661 4387 5695
rect 5733 5661 5767 5695
rect 7941 5661 7975 5695
rect 8401 5661 8435 5695
rect 10057 5661 10091 5695
rect 15485 5661 15519 5695
rect 32873 5661 32907 5695
rect 36829 5661 36863 5695
rect 38025 5661 38059 5695
rect 6377 5593 6411 5627
rect 7665 5593 7699 5627
rect 1777 5525 1811 5559
rect 5641 5525 5675 5559
rect 33057 5525 33091 5559
rect 36921 5525 36955 5559
rect 38209 5525 38243 5559
rect 4261 5321 4295 5355
rect 4997 5321 5031 5355
rect 1869 5185 1903 5219
rect 2697 5185 2731 5219
rect 3341 5185 3375 5219
rect 4445 5185 4479 5219
rect 4905 5185 4939 5219
rect 7665 5185 7699 5219
rect 7941 5185 7975 5219
rect 16865 5185 16899 5219
rect 20177 5185 20211 5219
rect 25513 5185 25547 5219
rect 27169 5185 27203 5219
rect 37473 5185 37507 5219
rect 2789 5117 2823 5151
rect 25697 5049 25731 5083
rect 1685 4981 1719 5015
rect 3433 4981 3467 5015
rect 17049 4981 17083 5015
rect 20361 4981 20395 5015
rect 27353 4981 27387 5015
rect 37657 4981 37691 5015
rect 1685 4777 1719 4811
rect 2973 4777 3007 4811
rect 4077 4777 4111 4811
rect 2329 4709 2363 4743
rect 9321 4641 9355 4675
rect 1777 4573 1811 4607
rect 2237 4573 2271 4607
rect 2881 4573 2915 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 7941 4573 7975 4607
rect 9597 4573 9631 4607
rect 16957 4573 16991 4607
rect 7665 4505 7699 4539
rect 4629 4437 4663 4471
rect 17141 4437 17175 4471
rect 1685 4097 1719 4131
rect 2789 4097 2823 4131
rect 3433 4097 3467 4131
rect 9781 4097 9815 4131
rect 1777 4029 1811 4063
rect 2881 4029 2915 4063
rect 3525 3961 3559 3995
rect 9689 3893 9723 3927
rect 2237 3689 2271 3723
rect 4169 3689 4203 3723
rect 38117 3689 38151 3723
rect 2881 3621 2915 3655
rect 2329 3485 2363 3519
rect 2789 3485 2823 3519
rect 3985 3485 4019 3519
rect 38301 3485 38335 3519
rect 2329 3145 2363 3179
rect 3065 3145 3099 3179
rect 36737 3145 36771 3179
rect 1593 3009 1627 3043
rect 2237 3009 2271 3043
rect 2881 3009 2915 3043
rect 3525 3009 3559 3043
rect 9597 3009 9631 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 3709 2873 3743 2907
rect 1777 2805 1811 2839
rect 9413 2805 9447 2839
rect 38209 2805 38243 2839
rect 2881 2601 2915 2635
rect 4813 2601 4847 2635
rect 6745 2601 6779 2635
rect 8033 2601 8067 2635
rect 10425 2601 10459 2635
rect 14473 2601 14507 2635
rect 15577 2601 15611 2635
rect 17049 2601 17083 2635
rect 22017 2601 22051 2635
rect 24593 2601 24627 2635
rect 27169 2601 27203 2635
rect 29745 2601 29779 2635
rect 32321 2601 32355 2635
rect 36737 2601 36771 2635
rect 34897 2533 34931 2567
rect 12633 2465 12667 2499
rect 1869 2397 1903 2431
rect 2697 2397 2731 2431
rect 4629 2397 4663 2431
rect 6561 2397 6595 2431
rect 7849 2397 7883 2431
rect 9413 2397 9447 2431
rect 10609 2397 10643 2431
rect 12357 2397 12391 2431
rect 14289 2397 14323 2431
rect 15761 2397 15795 2431
rect 16865 2397 16899 2431
rect 18613 2397 18647 2431
rect 20085 2397 20119 2431
rect 22201 2397 22235 2431
rect 23305 2397 23339 2431
rect 24777 2397 24811 2431
rect 27353 2397 27387 2431
rect 27813 2397 27847 2431
rect 29929 2397 29963 2431
rect 31033 2397 31067 2431
rect 32505 2397 32539 2431
rect 35081 2397 35115 2431
rect 35725 2397 35759 2431
rect 36921 2397 36955 2431
rect 37473 2397 37507 2431
rect 1685 2261 1719 2295
rect 9229 2261 9263 2295
rect 18797 2261 18831 2295
rect 20269 2261 20303 2295
rect 23489 2261 23523 2295
rect 27997 2261 28031 2295
rect 31217 2261 31251 2295
rect 35541 2261 35575 2295
rect 37657 2261 37691 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1854 37244 1860 37256
rect 1815 37216 1860 37244
rect 1854 37204 1860 37216
rect 1912 37204 1918 37256
rect 1946 37204 1952 37256
rect 2004 37244 2010 37256
rect 2317 37247 2375 37253
rect 2317 37244 2329 37247
rect 2004 37216 2329 37244
rect 2004 37204 2010 37216
rect 2317 37213 2329 37216
rect 2363 37213 2375 37247
rect 2958 37244 2964 37256
rect 2919 37216 2964 37244
rect 2317 37207 2375 37213
rect 2958 37204 2964 37216
rect 3016 37204 3022 37256
rect 4246 37244 4252 37256
rect 4207 37216 4252 37244
rect 4246 37204 4252 37216
rect 4304 37204 4310 37256
rect 5534 37244 5540 37256
rect 5495 37216 5540 37244
rect 5534 37204 5540 37216
rect 5592 37204 5598 37256
rect 7098 37204 7104 37256
rect 7156 37244 7162 37256
rect 7377 37247 7435 37253
rect 7377 37244 7389 37247
rect 7156 37216 7389 37244
rect 7156 37204 7162 37216
rect 7377 37213 7389 37216
rect 7423 37213 7435 37247
rect 7377 37207 7435 37213
rect 8386 37204 8392 37256
rect 8444 37244 8450 37256
rect 9309 37247 9367 37253
rect 9309 37244 9321 37247
rect 8444 37216 9321 37244
rect 8444 37204 8450 37216
rect 9309 37213 9321 37216
rect 9355 37213 9367 37247
rect 9309 37207 9367 37213
rect 10318 37204 10324 37256
rect 10376 37244 10382 37256
rect 10597 37247 10655 37253
rect 10597 37244 10609 37247
rect 10376 37216 10609 37244
rect 10376 37204 10382 37216
rect 10597 37213 10609 37216
rect 10643 37213 10655 37247
rect 10597 37207 10655 37213
rect 11606 37204 11612 37256
rect 11664 37244 11670 37256
rect 11885 37247 11943 37253
rect 11885 37244 11897 37247
rect 11664 37216 11897 37244
rect 11664 37204 11670 37216
rect 11885 37213 11897 37216
rect 11931 37213 11943 37247
rect 11885 37207 11943 37213
rect 12894 37204 12900 37256
rect 12952 37244 12958 37256
rect 12989 37247 13047 37253
rect 12989 37244 13001 37247
rect 12952 37216 13001 37244
rect 12952 37204 12958 37216
rect 12989 37213 13001 37216
rect 13035 37213 13047 37247
rect 15194 37244 15200 37256
rect 15155 37216 15200 37244
rect 12989 37207 13047 37213
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 16850 37244 16856 37256
rect 16811 37216 16856 37244
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 18138 37244 18144 37256
rect 18099 37216 18144 37244
rect 18138 37204 18144 37216
rect 18196 37204 18202 37256
rect 18230 37204 18236 37256
rect 18288 37244 18294 37256
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 18288 37216 19441 37244
rect 18288 37204 18294 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 19429 37207 19487 37213
rect 20714 37204 20720 37256
rect 20772 37244 20778 37256
rect 20901 37247 20959 37253
rect 20901 37244 20913 37247
rect 20772 37216 20913 37244
rect 20772 37204 20778 37216
rect 20901 37213 20913 37216
rect 20947 37213 20959 37247
rect 20901 37207 20959 37213
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 22612 37216 22845 37244
rect 22612 37204 22618 37216
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 22833 37207 22891 37213
rect 22922 37204 22928 37256
rect 22980 37244 22986 37256
rect 24581 37247 24639 37253
rect 24581 37244 24593 37247
rect 22980 37216 24593 37244
rect 22980 37204 22986 37216
rect 24581 37213 24593 37216
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 24762 37204 24768 37256
rect 24820 37244 24826 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 24820 37216 25881 37244
rect 24820 37204 24826 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 27062 37204 27068 37256
rect 27120 37244 27126 37256
rect 27341 37247 27399 37253
rect 27341 37244 27353 37247
rect 27120 37216 27353 37244
rect 27120 37204 27126 37216
rect 27341 37213 27353 37216
rect 27387 37213 27399 37247
rect 27341 37207 27399 37213
rect 27430 37204 27436 37256
rect 27488 37244 27494 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 27488 37216 29745 37244
rect 27488 37204 27494 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30653 37247 30711 37253
rect 30653 37244 30665 37247
rect 30432 37216 30665 37244
rect 30432 37204 30438 37216
rect 30653 37213 30665 37216
rect 30699 37213 30711 37247
rect 30653 37207 30711 37213
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 31812 37216 32505 37244
rect 31812 37204 31818 37216
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33560 37216 33793 37244
rect 33560 37204 33566 37216
rect 33781 37213 33793 37216
rect 33827 37213 33839 37247
rect 33781 37207 33839 37213
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34848 37216 35081 37244
rect 34848 37204 34854 37216
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 36722 37204 36728 37256
rect 36780 37244 36786 37256
rect 36909 37247 36967 37253
rect 36909 37244 36921 37247
rect 36780 37216 36921 37244
rect 36780 37204 36786 37216
rect 36909 37213 36921 37216
rect 36955 37213 36967 37247
rect 36909 37207 36967 37213
rect 38013 37247 38071 37253
rect 38013 37213 38025 37247
rect 38059 37213 38071 37247
rect 38013 37207 38071 37213
rect 2774 37176 2780 37188
rect 1688 37148 2780 37176
rect 1688 37117 1716 37148
rect 2774 37136 2780 37148
rect 2832 37136 2838 37188
rect 6546 37176 6552 37188
rect 2976 37148 6552 37176
rect 1673 37111 1731 37117
rect 1673 37077 1685 37111
rect 1719 37077 1731 37111
rect 1673 37071 1731 37077
rect 2501 37111 2559 37117
rect 2501 37077 2513 37111
rect 2547 37108 2559 37111
rect 2976 37108 3004 37148
rect 6546 37136 6552 37148
rect 6604 37136 6610 37188
rect 19978 37136 19984 37188
rect 20036 37176 20042 37188
rect 20036 37148 22692 37176
rect 20036 37136 20042 37148
rect 3142 37108 3148 37120
rect 2547 37080 3004 37108
rect 3103 37080 3148 37108
rect 2547 37077 2559 37080
rect 2501 37071 2559 37077
rect 3142 37068 3148 37080
rect 3200 37068 3206 37120
rect 3878 37068 3884 37120
rect 3936 37108 3942 37120
rect 4065 37111 4123 37117
rect 4065 37108 4077 37111
rect 3936 37080 4077 37108
rect 3936 37068 3942 37080
rect 4065 37077 4077 37080
rect 4111 37077 4123 37111
rect 4065 37071 4123 37077
rect 5166 37068 5172 37120
rect 5224 37108 5230 37120
rect 5353 37111 5411 37117
rect 5353 37108 5365 37111
rect 5224 37080 5365 37108
rect 5224 37068 5230 37080
rect 5353 37077 5365 37080
rect 5399 37077 5411 37111
rect 7190 37108 7196 37120
rect 7151 37080 7196 37108
rect 5353 37071 5411 37077
rect 7190 37068 7196 37080
rect 7248 37068 7254 37120
rect 8294 37068 8300 37120
rect 8352 37108 8358 37120
rect 9125 37111 9183 37117
rect 9125 37108 9137 37111
rect 8352 37080 9137 37108
rect 8352 37068 8358 37080
rect 9125 37077 9137 37080
rect 9171 37077 9183 37111
rect 9125 37071 9183 37077
rect 10318 37068 10324 37120
rect 10376 37108 10382 37120
rect 10413 37111 10471 37117
rect 10413 37108 10425 37111
rect 10376 37080 10425 37108
rect 10376 37068 10382 37080
rect 10413 37077 10425 37080
rect 10459 37077 10471 37111
rect 10413 37071 10471 37077
rect 10870 37068 10876 37120
rect 10928 37108 10934 37120
rect 11701 37111 11759 37117
rect 11701 37108 11713 37111
rect 10928 37080 11713 37108
rect 10928 37068 10934 37080
rect 11701 37077 11713 37080
rect 11747 37077 11759 37111
rect 11701 37071 11759 37077
rect 13173 37111 13231 37117
rect 13173 37077 13185 37111
rect 13219 37108 13231 37111
rect 14734 37108 14740 37120
rect 13219 37080 14740 37108
rect 13219 37077 13231 37080
rect 13173 37071 13231 37077
rect 14734 37068 14740 37080
rect 14792 37068 14798 37120
rect 14826 37068 14832 37120
rect 14884 37108 14890 37120
rect 15013 37111 15071 37117
rect 15013 37108 15025 37111
rect 14884 37080 15025 37108
rect 14884 37068 14890 37080
rect 15013 37077 15025 37080
rect 15059 37077 15071 37111
rect 15013 37071 15071 37077
rect 16574 37068 16580 37120
rect 16632 37108 16638 37120
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 16632 37080 17049 37108
rect 16632 37068 16638 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 17037 37071 17095 37077
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18325 37111 18383 37117
rect 18325 37108 18337 37111
rect 18104 37080 18337 37108
rect 18104 37068 18110 37080
rect 18325 37077 18337 37080
rect 18371 37077 18383 37111
rect 18325 37071 18383 37077
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 19613 37111 19671 37117
rect 19613 37108 19625 37111
rect 19392 37080 19625 37108
rect 19392 37068 19398 37080
rect 19613 37077 19625 37080
rect 19659 37077 19671 37111
rect 20714 37108 20720 37120
rect 20675 37080 20720 37108
rect 19613 37071 19671 37077
rect 20714 37068 20720 37080
rect 20772 37068 20778 37120
rect 22664 37117 22692 37148
rect 29362 37136 29368 37188
rect 29420 37176 29426 37188
rect 29420 37148 33640 37176
rect 29420 37136 29426 37148
rect 22649 37111 22707 37117
rect 22649 37077 22661 37111
rect 22695 37077 22707 37111
rect 22649 37071 22707 37077
rect 23842 37068 23848 37120
rect 23900 37108 23906 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 23900 37080 24777 37108
rect 23900 37068 23906 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25774 37068 25780 37120
rect 25832 37108 25838 37120
rect 26053 37111 26111 37117
rect 26053 37108 26065 37111
rect 25832 37080 26065 37108
rect 25832 37068 25838 37080
rect 26053 37077 26065 37080
rect 26099 37077 26111 37111
rect 27154 37108 27160 37120
rect 27115 37080 27160 37108
rect 26053 37071 26111 37077
rect 27154 37068 27160 37080
rect 27212 37068 27218 37120
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29052 37080 29929 37108
rect 29052 37068 29058 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 30466 37108 30472 37120
rect 30427 37080 30472 37108
rect 29917 37071 29975 37077
rect 30466 37068 30472 37080
rect 30524 37068 30530 37120
rect 32306 37108 32312 37120
rect 32267 37080 32312 37108
rect 32306 37068 32312 37080
rect 32364 37068 32370 37120
rect 33612 37117 33640 37148
rect 33962 37136 33968 37188
rect 34020 37176 34026 37188
rect 38028 37176 38056 37207
rect 34020 37148 38056 37176
rect 34020 37136 34026 37148
rect 33597 37111 33655 37117
rect 33597 37077 33609 37111
rect 33643 37077 33655 37111
rect 34882 37108 34888 37120
rect 34843 37080 34888 37108
rect 33597 37071 33655 37077
rect 34882 37068 34888 37080
rect 34940 37068 34946 37120
rect 35894 37068 35900 37120
rect 35952 37108 35958 37120
rect 36725 37111 36783 37117
rect 36725 37108 36737 37111
rect 35952 37080 36737 37108
rect 35952 37068 35958 37080
rect 36725 37077 36737 37080
rect 36771 37077 36783 37111
rect 38194 37108 38200 37120
rect 38155 37080 38200 37108
rect 36725 37071 36783 37077
rect 38194 37068 38200 37080
rect 38252 37068 38258 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 658 36864 664 36916
rect 716 36904 722 36916
rect 1673 36907 1731 36913
rect 1673 36904 1685 36907
rect 716 36876 1685 36904
rect 716 36864 722 36876
rect 1673 36873 1685 36876
rect 1719 36873 1731 36907
rect 1673 36867 1731 36873
rect 1854 36864 1860 36916
rect 1912 36904 1918 36916
rect 3970 36904 3976 36916
rect 1912 36876 3976 36904
rect 1912 36864 1918 36876
rect 3970 36864 3976 36876
rect 4028 36864 4034 36916
rect 30282 36864 30288 36916
rect 30340 36904 30346 36916
rect 34882 36904 34888 36916
rect 30340 36876 34888 36904
rect 30340 36864 30346 36876
rect 34882 36864 34888 36876
rect 34940 36864 34946 36916
rect 39298 36836 39304 36848
rect 36924 36808 39304 36836
rect 1857 36771 1915 36777
rect 1857 36737 1869 36771
rect 1903 36768 1915 36771
rect 4062 36768 4068 36780
rect 1903 36740 4068 36768
rect 1903 36737 1915 36740
rect 1857 36731 1915 36737
rect 4062 36728 4068 36740
rect 4120 36728 4126 36780
rect 36924 36777 36952 36808
rect 39298 36796 39304 36808
rect 39356 36796 39362 36848
rect 36909 36771 36967 36777
rect 36909 36737 36921 36771
rect 36955 36737 36967 36771
rect 37550 36768 37556 36780
rect 37511 36740 37556 36768
rect 36909 36731 36967 36737
rect 37550 36728 37556 36740
rect 37608 36728 37614 36780
rect 36722 36564 36728 36576
rect 36683 36536 36728 36564
rect 36722 36524 36728 36536
rect 36780 36524 36786 36576
rect 37366 36524 37372 36576
rect 37424 36564 37430 36576
rect 37553 36567 37611 36573
rect 37553 36564 37565 36567
rect 37424 36536 37565 36564
rect 37424 36524 37430 36536
rect 37553 36533 37565 36536
rect 37599 36533 37611 36567
rect 37553 36527 37611 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 37182 36320 37188 36372
rect 37240 36360 37246 36372
rect 38197 36363 38255 36369
rect 38197 36360 38209 36363
rect 37240 36332 38209 36360
rect 37240 36320 37246 36332
rect 38197 36329 38209 36332
rect 38243 36329 38255 36363
rect 38197 36323 38255 36329
rect 1578 36156 1584 36168
rect 1539 36128 1584 36156
rect 1578 36116 1584 36128
rect 1636 36116 1642 36168
rect 37366 36156 37372 36168
rect 37327 36128 37372 36156
rect 37366 36116 37372 36128
rect 37424 36116 37430 36168
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 37568 36128 38025 36156
rect 1765 36023 1823 36029
rect 1765 35989 1777 36023
rect 1811 36020 1823 36023
rect 6638 36020 6644 36032
rect 1811 35992 6644 36020
rect 1811 35989 1823 35992
rect 1765 35983 1823 35989
rect 6638 35980 6644 35992
rect 6696 35980 6702 36032
rect 37568 36029 37596 36128
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 37553 36023 37611 36029
rect 37553 35989 37565 36023
rect 37599 35989 37611 36023
rect 37553 35983 37611 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 5534 35776 5540 35828
rect 5592 35816 5598 35828
rect 5721 35819 5779 35825
rect 5721 35816 5733 35819
rect 5592 35788 5733 35816
rect 5592 35776 5598 35788
rect 5721 35785 5733 35788
rect 5767 35785 5779 35819
rect 16850 35816 16856 35828
rect 16811 35788 16856 35816
rect 5721 35779 5779 35785
rect 16850 35776 16856 35788
rect 16908 35776 16914 35828
rect 5902 35680 5908 35692
rect 5863 35652 5908 35680
rect 5902 35640 5908 35652
rect 5960 35640 5966 35692
rect 17034 35680 17040 35692
rect 16995 35652 17040 35680
rect 17034 35640 17040 35652
rect 17092 35640 17098 35692
rect 38010 35640 38016 35692
rect 38068 35680 38074 35692
rect 38289 35683 38347 35689
rect 38289 35680 38301 35683
rect 38068 35652 38301 35680
rect 38068 35640 38074 35652
rect 38289 35649 38301 35652
rect 38335 35649 38347 35683
rect 38289 35643 38347 35649
rect 33226 35436 33232 35488
rect 33284 35476 33290 35488
rect 38105 35479 38163 35485
rect 38105 35476 38117 35479
rect 33284 35448 38117 35476
rect 33284 35436 33290 35448
rect 38105 35445 38117 35448
rect 38151 35445 38163 35479
rect 38105 35439 38163 35445
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 3970 35232 3976 35284
rect 4028 35272 4034 35284
rect 6457 35275 6515 35281
rect 6457 35272 6469 35275
rect 4028 35244 6469 35272
rect 4028 35232 4034 35244
rect 6457 35241 6469 35244
rect 6503 35241 6515 35275
rect 6457 35235 6515 35241
rect 17681 35275 17739 35281
rect 17681 35241 17693 35275
rect 17727 35272 17739 35275
rect 18138 35272 18144 35284
rect 17727 35244 18144 35272
rect 17727 35241 17739 35244
rect 17681 35235 17739 35241
rect 18138 35232 18144 35244
rect 18196 35232 18202 35284
rect 17037 35207 17095 35213
rect 17037 35173 17049 35207
rect 17083 35204 17095 35207
rect 18230 35204 18236 35216
rect 17083 35176 18236 35204
rect 17083 35173 17095 35176
rect 17037 35167 17095 35173
rect 18230 35164 18236 35176
rect 18288 35164 18294 35216
rect 6641 35071 6699 35077
rect 6641 35037 6653 35071
rect 6687 35068 6699 35071
rect 6730 35068 6736 35080
rect 6687 35040 6736 35068
rect 6687 35037 6699 35040
rect 6641 35031 6699 35037
rect 6730 35028 6736 35040
rect 6788 35028 6794 35080
rect 16482 35028 16488 35080
rect 16540 35068 16546 35080
rect 16853 35071 16911 35077
rect 16853 35068 16865 35071
rect 16540 35040 16865 35068
rect 16540 35028 16546 35040
rect 16853 35037 16865 35040
rect 16899 35037 16911 35071
rect 17494 35068 17500 35080
rect 17455 35040 17500 35068
rect 16853 35031 16911 35037
rect 17494 35028 17500 35040
rect 17552 35028 17558 35080
rect 35342 35028 35348 35080
rect 35400 35068 35406 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 35400 35040 38025 35068
rect 35400 35028 35406 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 38194 34932 38200 34944
rect 38155 34904 38200 34932
rect 38194 34892 38200 34904
rect 38252 34892 38258 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 4062 34688 4068 34740
rect 4120 34728 4126 34740
rect 6733 34731 6791 34737
rect 6733 34728 6745 34731
rect 4120 34700 6745 34728
rect 4120 34688 4126 34700
rect 6733 34697 6745 34700
rect 6779 34697 6791 34731
rect 6733 34691 6791 34697
rect 15194 34688 15200 34740
rect 15252 34728 15258 34740
rect 15473 34731 15531 34737
rect 15473 34728 15485 34731
rect 15252 34700 15485 34728
rect 15252 34688 15258 34700
rect 15473 34697 15485 34700
rect 15519 34697 15531 34731
rect 15473 34691 15531 34697
rect 21361 34731 21419 34737
rect 21361 34697 21373 34731
rect 21407 34697 21419 34731
rect 21361 34691 21419 34697
rect 22833 34731 22891 34737
rect 22833 34697 22845 34731
rect 22879 34728 22891 34731
rect 24762 34728 24768 34740
rect 22879 34700 24768 34728
rect 22879 34697 22891 34700
rect 22833 34691 22891 34697
rect 20070 34620 20076 34672
rect 20128 34660 20134 34672
rect 21376 34660 21404 34691
rect 24762 34688 24768 34700
rect 24820 34688 24826 34740
rect 25777 34731 25835 34737
rect 25777 34697 25789 34731
rect 25823 34728 25835 34731
rect 27430 34728 27436 34740
rect 25823 34700 27436 34728
rect 25823 34697 25835 34700
rect 25777 34691 25835 34697
rect 27430 34688 27436 34700
rect 27488 34688 27494 34740
rect 22922 34660 22928 34672
rect 20128 34632 21220 34660
rect 21376 34632 22928 34660
rect 20128 34620 20134 34632
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34592 1915 34595
rect 3970 34592 3976 34604
rect 1903 34564 3976 34592
rect 1903 34561 1915 34564
rect 1857 34555 1915 34561
rect 3970 34552 3976 34564
rect 4028 34552 4034 34604
rect 6917 34595 6975 34601
rect 6917 34561 6929 34595
rect 6963 34592 6975 34595
rect 12066 34592 12072 34604
rect 6963 34564 12072 34592
rect 6963 34561 6975 34564
rect 6917 34555 6975 34561
rect 12066 34552 12072 34564
rect 12124 34552 12130 34604
rect 14734 34552 14740 34604
rect 14792 34592 14798 34604
rect 14829 34595 14887 34601
rect 14829 34592 14841 34595
rect 14792 34564 14841 34592
rect 14792 34552 14798 34564
rect 14829 34561 14841 34564
rect 14875 34561 14887 34595
rect 15654 34592 15660 34604
rect 15615 34564 15660 34592
rect 14829 34555 14887 34561
rect 15654 34552 15660 34564
rect 15712 34552 15718 34604
rect 20714 34592 20720 34604
rect 20675 34564 20720 34592
rect 20714 34552 20720 34564
rect 20772 34552 20778 34604
rect 21192 34601 21220 34632
rect 22922 34620 22928 34632
rect 22980 34620 22986 34672
rect 21177 34595 21235 34601
rect 21177 34561 21189 34595
rect 21223 34561 21235 34595
rect 21177 34555 21235 34561
rect 21266 34552 21272 34604
rect 21324 34592 21330 34604
rect 22649 34595 22707 34601
rect 22649 34592 22661 34595
rect 21324 34564 22661 34592
rect 21324 34552 21330 34564
rect 22649 34561 22661 34564
rect 22695 34561 22707 34595
rect 22649 34555 22707 34561
rect 24670 34552 24676 34604
rect 24728 34592 24734 34604
rect 25593 34595 25651 34601
rect 25593 34592 25605 34595
rect 24728 34564 25605 34592
rect 24728 34552 24734 34564
rect 25593 34561 25605 34564
rect 25639 34561 25651 34595
rect 33226 34592 33232 34604
rect 33187 34564 33232 34592
rect 25593 34555 25651 34561
rect 33226 34552 33232 34564
rect 33284 34552 33290 34604
rect 14921 34527 14979 34533
rect 14921 34493 14933 34527
rect 14967 34524 14979 34527
rect 16114 34524 16120 34536
rect 14967 34496 16120 34524
rect 14967 34493 14979 34496
rect 14921 34487 14979 34493
rect 16114 34484 16120 34496
rect 16172 34484 16178 34536
rect 20346 34484 20352 34536
rect 20404 34524 20410 34536
rect 20625 34527 20683 34533
rect 20625 34524 20637 34527
rect 20404 34496 20637 34524
rect 20404 34484 20410 34496
rect 20625 34493 20637 34496
rect 20671 34493 20683 34527
rect 33134 34524 33140 34536
rect 33095 34496 33140 34524
rect 20625 34487 20683 34493
rect 33134 34484 33140 34496
rect 33192 34484 33198 34536
rect 1670 34388 1676 34400
rect 1631 34360 1676 34388
rect 1670 34348 1676 34360
rect 1728 34348 1734 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 10870 34048 10876 34060
rect 9876 34020 10876 34048
rect 9876 33989 9904 34020
rect 10870 34008 10876 34020
rect 10928 34008 10934 34060
rect 9861 33983 9919 33989
rect 9861 33949 9873 33983
rect 9907 33949 9919 33983
rect 10318 33980 10324 33992
rect 10279 33952 10324 33980
rect 9861 33943 9919 33949
rect 10318 33940 10324 33952
rect 10376 33940 10382 33992
rect 30282 33980 30288 33992
rect 30243 33952 30288 33980
rect 30282 33940 30288 33952
rect 30340 33940 30346 33992
rect 8386 33804 8392 33856
rect 8444 33844 8450 33856
rect 9769 33847 9827 33853
rect 9769 33844 9781 33847
rect 8444 33816 9781 33844
rect 8444 33804 8450 33816
rect 9769 33813 9781 33816
rect 9815 33813 9827 33847
rect 9769 33807 9827 33813
rect 10226 33804 10232 33856
rect 10284 33844 10290 33856
rect 10413 33847 10471 33853
rect 10413 33844 10425 33847
rect 10284 33816 10425 33844
rect 10284 33804 10290 33816
rect 10413 33813 10425 33816
rect 10459 33813 10471 33847
rect 10413 33807 10471 33813
rect 18782 33804 18788 33856
rect 18840 33844 18846 33856
rect 30193 33847 30251 33853
rect 30193 33844 30205 33847
rect 18840 33816 30205 33844
rect 18840 33804 18846 33816
rect 30193 33813 30205 33816
rect 30239 33813 30251 33847
rect 30193 33807 30251 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 14277 33643 14335 33649
rect 14277 33609 14289 33643
rect 14323 33640 14335 33643
rect 15654 33640 15660 33652
rect 14323 33612 15660 33640
rect 14323 33609 14335 33612
rect 14277 33603 14335 33609
rect 15654 33600 15660 33612
rect 15712 33600 15718 33652
rect 13538 33464 13544 33516
rect 13596 33504 13602 33516
rect 14185 33507 14243 33513
rect 14185 33504 14197 33507
rect 13596 33476 14197 33504
rect 13596 33464 13602 33476
rect 14185 33473 14197 33476
rect 14231 33473 14243 33507
rect 19978 33504 19984 33516
rect 19939 33476 19984 33504
rect 14185 33467 14243 33473
rect 19978 33464 19984 33476
rect 20036 33464 20042 33516
rect 29362 33504 29368 33516
rect 29323 33476 29368 33504
rect 29362 33464 29368 33476
rect 29420 33464 29426 33516
rect 33502 33464 33508 33516
rect 33560 33504 33566 33516
rect 38013 33507 38071 33513
rect 38013 33504 38025 33507
rect 33560 33476 38025 33504
rect 33560 33464 33566 33476
rect 38013 33473 38025 33476
rect 38059 33473 38071 33507
rect 38013 33467 38071 33473
rect 12158 33328 12164 33380
rect 12216 33368 12222 33380
rect 29273 33371 29331 33377
rect 29273 33368 29285 33371
rect 12216 33340 29285 33368
rect 12216 33328 12222 33340
rect 29273 33337 29285 33340
rect 29319 33337 29331 33371
rect 38194 33368 38200 33380
rect 38155 33340 38200 33368
rect 29273 33331 29331 33337
rect 38194 33328 38200 33340
rect 38252 33328 38258 33380
rect 17586 33260 17592 33312
rect 17644 33300 17650 33312
rect 19889 33303 19947 33309
rect 19889 33300 19901 33303
rect 17644 33272 19901 33300
rect 17644 33260 17650 33272
rect 19889 33269 19901 33272
rect 19935 33269 19947 33303
rect 19889 33263 19947 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1578 32892 1584 32904
rect 1539 32864 1584 32892
rect 1578 32852 1584 32864
rect 1636 32852 1642 32904
rect 1765 32759 1823 32765
rect 1765 32725 1777 32759
rect 1811 32756 1823 32759
rect 4614 32756 4620 32768
rect 1811 32728 4620 32756
rect 1811 32725 1823 32728
rect 1765 32719 1823 32725
rect 4614 32716 4620 32728
rect 4672 32716 4678 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 33962 32552 33968 32564
rect 33923 32524 33968 32552
rect 33962 32512 33968 32524
rect 34020 32512 34026 32564
rect 3142 32376 3148 32428
rect 3200 32416 3206 32428
rect 5261 32419 5319 32425
rect 5261 32416 5273 32419
rect 3200 32388 5273 32416
rect 3200 32376 3206 32388
rect 5261 32385 5273 32388
rect 5307 32385 5319 32419
rect 5261 32379 5319 32385
rect 33226 32376 33232 32428
rect 33284 32416 33290 32428
rect 33781 32419 33839 32425
rect 33781 32416 33793 32419
rect 33284 32388 33793 32416
rect 33284 32376 33290 32388
rect 33781 32385 33793 32388
rect 33827 32385 33839 32419
rect 33781 32379 33839 32385
rect 5353 32215 5411 32221
rect 5353 32181 5365 32215
rect 5399 32212 5411 32215
rect 6178 32212 6184 32224
rect 5399 32184 6184 32212
rect 5399 32181 5411 32184
rect 5353 32175 5411 32181
rect 6178 32172 6184 32184
rect 6236 32172 6242 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 33778 31900 33784 31952
rect 33836 31940 33842 31952
rect 38105 31943 38163 31949
rect 38105 31940 38117 31943
rect 33836 31912 38117 31940
rect 33836 31900 33842 31912
rect 38105 31909 38117 31912
rect 38151 31909 38163 31943
rect 38105 31903 38163 31909
rect 18966 31764 18972 31816
rect 19024 31804 19030 31816
rect 23201 31807 23259 31813
rect 23201 31804 23213 31807
rect 19024 31776 23213 31804
rect 19024 31764 19030 31776
rect 23201 31773 23213 31776
rect 23247 31773 23259 31807
rect 23201 31767 23259 31773
rect 23293 31807 23351 31813
rect 23293 31773 23305 31807
rect 23339 31804 23351 31807
rect 27154 31804 27160 31816
rect 23339 31776 27160 31804
rect 23339 31773 23351 31776
rect 23293 31767 23351 31773
rect 27154 31764 27160 31776
rect 27212 31764 27218 31816
rect 38286 31804 38292 31816
rect 38247 31776 38292 31804
rect 38286 31764 38292 31776
rect 38344 31764 38350 31816
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 16945 31467 17003 31473
rect 16945 31433 16957 31467
rect 16991 31464 17003 31467
rect 17034 31464 17040 31476
rect 16991 31436 17040 31464
rect 16991 31433 17003 31436
rect 16945 31427 17003 31433
rect 17034 31424 17040 31436
rect 17092 31424 17098 31476
rect 16666 31288 16672 31340
rect 16724 31328 16730 31340
rect 16853 31331 16911 31337
rect 16853 31328 16865 31331
rect 16724 31300 16865 31328
rect 16724 31288 16730 31300
rect 16853 31297 16865 31300
rect 16899 31297 16911 31331
rect 16853 31291 16911 31297
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 3970 30920 3976 30932
rect 3931 30892 3976 30920
rect 3970 30880 3976 30892
rect 4028 30880 4034 30932
rect 5902 30880 5908 30932
rect 5960 30920 5966 30932
rect 6181 30923 6239 30929
rect 6181 30920 6193 30923
rect 5960 30892 6193 30920
rect 5960 30880 5966 30892
rect 6181 30889 6193 30892
rect 6227 30889 6239 30923
rect 6181 30883 6239 30889
rect 35069 30923 35127 30929
rect 35069 30889 35081 30923
rect 35115 30920 35127 30923
rect 35342 30920 35348 30932
rect 35115 30892 35348 30920
rect 35115 30889 35127 30892
rect 35069 30883 35127 30889
rect 35342 30880 35348 30892
rect 35400 30880 35406 30932
rect 1765 30855 1823 30861
rect 1765 30821 1777 30855
rect 1811 30852 1823 30855
rect 9122 30852 9128 30864
rect 1811 30824 9128 30852
rect 1811 30821 1823 30824
rect 1765 30815 1823 30821
rect 9122 30812 9128 30824
rect 9180 30812 9186 30864
rect 1578 30716 1584 30728
rect 1539 30688 1584 30716
rect 1578 30676 1584 30688
rect 1636 30676 1642 30728
rect 4062 30676 4068 30728
rect 4120 30716 4126 30728
rect 4157 30719 4215 30725
rect 4157 30716 4169 30719
rect 4120 30688 4169 30716
rect 4120 30676 4126 30688
rect 4157 30685 4169 30688
rect 4203 30685 4215 30719
rect 6270 30716 6276 30728
rect 6231 30688 6276 30716
rect 4157 30679 4215 30685
rect 6270 30676 6276 30688
rect 6328 30676 6334 30728
rect 8294 30716 8300 30728
rect 8255 30688 8300 30716
rect 8294 30676 8300 30688
rect 8352 30676 8358 30728
rect 33870 30676 33876 30728
rect 33928 30716 33934 30728
rect 34885 30719 34943 30725
rect 34885 30716 34897 30719
rect 33928 30688 34897 30716
rect 33928 30676 33934 30688
rect 34885 30685 34897 30688
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 8202 30580 8208 30592
rect 8163 30552 8208 30580
rect 8202 30540 8208 30552
rect 8260 30540 8266 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 6730 30268 6736 30320
rect 6788 30308 6794 30320
rect 11793 30311 11851 30317
rect 11793 30308 11805 30311
rect 6788 30280 11805 30308
rect 6788 30268 6794 30280
rect 11793 30277 11805 30280
rect 11839 30277 11851 30311
rect 11793 30271 11851 30277
rect 20901 30311 20959 30317
rect 20901 30277 20913 30311
rect 20947 30308 20959 30311
rect 21266 30308 21272 30320
rect 20947 30280 21272 30308
rect 20947 30277 20959 30280
rect 20901 30271 20959 30277
rect 21266 30268 21272 30280
rect 21324 30268 21330 30320
rect 35894 30308 35900 30320
rect 29288 30280 35900 30308
rect 2685 30243 2743 30249
rect 2685 30209 2697 30243
rect 2731 30240 2743 30243
rect 2958 30240 2964 30252
rect 2731 30212 2964 30240
rect 2731 30209 2743 30212
rect 2685 30203 2743 30209
rect 2958 30200 2964 30212
rect 3016 30200 3022 30252
rect 6546 30240 6552 30252
rect 6507 30212 6552 30240
rect 6546 30200 6552 30212
rect 6604 30200 6610 30252
rect 11885 30243 11943 30249
rect 11885 30209 11897 30243
rect 11931 30240 11943 30243
rect 12986 30240 12992 30252
rect 11931 30212 12992 30240
rect 11931 30209 11943 30212
rect 11885 30203 11943 30209
rect 12986 30200 12992 30212
rect 13044 30200 13050 30252
rect 17126 30200 17132 30252
rect 17184 30240 17190 30252
rect 29288 30249 29316 30280
rect 35894 30268 35900 30280
rect 35952 30268 35958 30320
rect 20809 30243 20867 30249
rect 20809 30240 20821 30243
rect 17184 30212 20821 30240
rect 17184 30200 17190 30212
rect 20809 30209 20821 30212
rect 20855 30209 20867 30243
rect 20809 30203 20867 30209
rect 27341 30243 27399 30249
rect 27341 30209 27353 30243
rect 27387 30209 27399 30243
rect 27341 30203 27399 30209
rect 29273 30243 29331 30249
rect 29273 30209 29285 30243
rect 29319 30209 29331 30243
rect 33318 30240 33324 30252
rect 33279 30212 33324 30240
rect 29273 30203 29331 30209
rect 2222 30132 2228 30184
rect 2280 30172 2286 30184
rect 2409 30175 2467 30181
rect 2409 30172 2421 30175
rect 2280 30144 2421 30172
rect 2280 30132 2286 30144
rect 2409 30141 2421 30144
rect 2455 30141 2467 30175
rect 27356 30172 27384 30203
rect 33318 30200 33324 30212
rect 33376 30200 33382 30252
rect 38286 30240 38292 30252
rect 38247 30212 38292 30240
rect 38286 30200 38292 30212
rect 38344 30200 38350 30252
rect 32306 30172 32312 30184
rect 27356 30144 32312 30172
rect 2409 30135 2467 30141
rect 32306 30132 32312 30144
rect 32364 30132 32370 30184
rect 33502 30104 33508 30116
rect 33463 30076 33508 30104
rect 33502 30064 33508 30076
rect 33560 30064 33566 30116
rect 6641 30039 6699 30045
rect 6641 30005 6653 30039
rect 6687 30036 6699 30039
rect 7742 30036 7748 30048
rect 6687 30008 7748 30036
rect 6687 30005 6699 30008
rect 6641 29999 6699 30005
rect 7742 29996 7748 30008
rect 7800 29996 7806 30048
rect 27246 30036 27252 30048
rect 27207 30008 27252 30036
rect 27246 29996 27252 30008
rect 27304 29996 27310 30048
rect 29178 30036 29184 30048
rect 29139 30008 29184 30036
rect 29178 29996 29184 30008
rect 29236 29996 29242 30048
rect 35434 29996 35440 30048
rect 35492 30036 35498 30048
rect 38105 30039 38163 30045
rect 38105 30036 38117 30039
rect 35492 30008 38117 30036
rect 35492 29996 35498 30008
rect 38105 30005 38117 30008
rect 38151 30005 38163 30039
rect 38105 29999 38163 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 12066 29832 12072 29844
rect 12027 29804 12072 29832
rect 12066 29792 12072 29804
rect 12124 29792 12130 29844
rect 16482 29832 16488 29844
rect 16443 29804 16488 29832
rect 16482 29792 16488 29804
rect 16540 29792 16546 29844
rect 17129 29835 17187 29841
rect 17129 29801 17141 29835
rect 17175 29832 17187 29835
rect 17494 29832 17500 29844
rect 17175 29804 17500 29832
rect 17175 29801 17187 29804
rect 17129 29795 17187 29801
rect 17494 29792 17500 29804
rect 17552 29792 17558 29844
rect 24670 29832 24676 29844
rect 24631 29804 24676 29832
rect 24670 29792 24676 29804
rect 24728 29792 24734 29844
rect 2590 29696 2596 29708
rect 2551 29668 2596 29696
rect 2590 29656 2596 29668
rect 2648 29656 2654 29708
rect 5169 29699 5227 29705
rect 5169 29665 5181 29699
rect 5215 29696 5227 29699
rect 9858 29696 9864 29708
rect 5215 29668 9864 29696
rect 5215 29665 5227 29668
rect 5169 29659 5227 29665
rect 9858 29656 9864 29668
rect 9916 29656 9922 29708
rect 1857 29631 1915 29637
rect 1857 29597 1869 29631
rect 1903 29628 1915 29631
rect 2777 29631 2835 29637
rect 1903 29600 2636 29628
rect 1903 29597 1915 29600
rect 1857 29591 1915 29597
rect 2608 29560 2636 29600
rect 2777 29597 2789 29631
rect 2823 29628 2835 29631
rect 2958 29628 2964 29640
rect 2823 29600 2964 29628
rect 2823 29597 2835 29600
rect 2777 29591 2835 29597
rect 2958 29588 2964 29600
rect 3016 29588 3022 29640
rect 4982 29588 4988 29640
rect 5040 29628 5046 29640
rect 5077 29631 5135 29637
rect 5077 29628 5089 29631
rect 5040 29600 5089 29628
rect 5040 29588 5046 29600
rect 5077 29597 5089 29600
rect 5123 29628 5135 29631
rect 5721 29631 5779 29637
rect 5721 29628 5733 29631
rect 5123 29600 5733 29628
rect 5123 29597 5135 29600
rect 5077 29591 5135 29597
rect 5721 29597 5733 29600
rect 5767 29628 5779 29631
rect 6365 29631 6423 29637
rect 6365 29628 6377 29631
rect 5767 29600 6377 29628
rect 5767 29597 5779 29600
rect 5721 29591 5779 29597
rect 6365 29597 6377 29600
rect 6411 29597 6423 29631
rect 6365 29591 6423 29597
rect 12161 29631 12219 29637
rect 12161 29597 12173 29631
rect 12207 29628 12219 29631
rect 12207 29600 12434 29628
rect 12207 29597 12219 29600
rect 12161 29591 12219 29597
rect 3602 29560 3608 29572
rect 2608 29532 3608 29560
rect 3602 29520 3608 29532
rect 3660 29520 3666 29572
rect 5813 29563 5871 29569
rect 5813 29529 5825 29563
rect 5859 29560 5871 29563
rect 7466 29560 7472 29572
rect 5859 29532 7472 29560
rect 5859 29529 5871 29532
rect 5813 29523 5871 29529
rect 7466 29520 7472 29532
rect 7524 29520 7530 29572
rect 12406 29560 12434 29600
rect 14642 29588 14648 29640
rect 14700 29628 14706 29640
rect 16393 29631 16451 29637
rect 16393 29628 16405 29631
rect 14700 29600 16405 29628
rect 14700 29588 14706 29600
rect 16393 29597 16405 29600
rect 16439 29597 16451 29631
rect 17034 29628 17040 29640
rect 16995 29600 17040 29628
rect 16393 29591 16451 29597
rect 17034 29588 17040 29600
rect 17092 29588 17098 29640
rect 23382 29588 23388 29640
rect 23440 29628 23446 29640
rect 24581 29631 24639 29637
rect 24581 29628 24593 29631
rect 23440 29600 24593 29628
rect 23440 29588 23446 29600
rect 24581 29597 24593 29600
rect 24627 29597 24639 29631
rect 24581 29591 24639 29597
rect 25501 29631 25559 29637
rect 25501 29597 25513 29631
rect 25547 29628 25559 29631
rect 30466 29628 30472 29640
rect 25547 29600 30472 29628
rect 25547 29597 25559 29600
rect 25501 29591 25559 29597
rect 30466 29588 30472 29600
rect 30524 29588 30530 29640
rect 30561 29631 30619 29637
rect 30561 29597 30573 29631
rect 30607 29628 30619 29631
rect 36722 29628 36728 29640
rect 30607 29600 36728 29628
rect 30607 29597 30619 29600
rect 30561 29591 30619 29597
rect 36722 29588 36728 29600
rect 36780 29588 36786 29640
rect 15378 29560 15384 29572
rect 12406 29532 15384 29560
rect 15378 29520 15384 29532
rect 15436 29520 15442 29572
rect 1670 29492 1676 29504
rect 1631 29464 1676 29492
rect 1670 29452 1676 29464
rect 1728 29452 1734 29504
rect 6457 29495 6515 29501
rect 6457 29461 6469 29495
rect 6503 29492 6515 29495
rect 8018 29492 8024 29504
rect 6503 29464 8024 29492
rect 6503 29461 6515 29464
rect 6457 29455 6515 29461
rect 8018 29452 8024 29464
rect 8076 29452 8082 29504
rect 25406 29492 25412 29504
rect 25367 29464 25412 29492
rect 25406 29452 25412 29464
rect 25464 29452 25470 29504
rect 30466 29492 30472 29504
rect 30427 29464 30472 29492
rect 30466 29452 30472 29464
rect 30524 29452 30530 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1578 29152 1584 29164
rect 1539 29124 1584 29152
rect 1578 29112 1584 29124
rect 1636 29112 1642 29164
rect 2777 29155 2835 29161
rect 2777 29121 2789 29155
rect 2823 29152 2835 29155
rect 4341 29155 4399 29161
rect 2823 29124 3004 29152
rect 2823 29121 2835 29124
rect 2777 29115 2835 29121
rect 2976 29096 3004 29124
rect 4341 29121 4353 29155
rect 4387 29152 4399 29155
rect 4614 29152 4620 29164
rect 4387 29124 4620 29152
rect 4387 29121 4399 29124
rect 4341 29115 4399 29121
rect 4614 29112 4620 29124
rect 4672 29112 4678 29164
rect 4982 29152 4988 29164
rect 4724 29124 4988 29152
rect 2314 29044 2320 29096
rect 2372 29084 2378 29096
rect 2501 29087 2559 29093
rect 2501 29084 2513 29087
rect 2372 29056 2513 29084
rect 2372 29044 2378 29056
rect 2501 29053 2513 29056
rect 2547 29053 2559 29087
rect 2501 29047 2559 29053
rect 2958 29044 2964 29096
rect 3016 29084 3022 29096
rect 4724 29084 4752 29124
rect 4982 29112 4988 29124
rect 5040 29112 5046 29164
rect 38010 29152 38016 29164
rect 37971 29124 38016 29152
rect 38010 29112 38016 29124
rect 38068 29112 38074 29164
rect 5074 29084 5080 29096
rect 3016 29056 4752 29084
rect 5035 29056 5080 29084
rect 3016 29044 3022 29056
rect 5074 29044 5080 29056
rect 5132 29044 5138 29096
rect 1765 29019 1823 29025
rect 1765 28985 1777 29019
rect 1811 29016 1823 29019
rect 3878 29016 3884 29028
rect 1811 28988 3884 29016
rect 1811 28985 1823 28988
rect 1765 28979 1823 28985
rect 3878 28976 3884 28988
rect 3936 28976 3942 29028
rect 4433 29019 4491 29025
rect 4433 28985 4445 29019
rect 4479 29016 4491 29019
rect 5350 29016 5356 29028
rect 4479 28988 5356 29016
rect 4479 28985 4491 28988
rect 4433 28979 4491 28985
rect 5350 28976 5356 28988
rect 5408 28976 5414 29028
rect 38194 29016 38200 29028
rect 38155 28988 38200 29016
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 4062 28744 4068 28756
rect 4023 28716 4068 28744
rect 4062 28704 4068 28716
rect 4120 28704 4126 28756
rect 19705 28747 19763 28753
rect 19705 28713 19717 28747
rect 19751 28744 19763 28747
rect 20070 28744 20076 28756
rect 19751 28716 20076 28744
rect 19751 28713 19763 28716
rect 19705 28707 19763 28713
rect 20070 28704 20076 28716
rect 20128 28704 20134 28756
rect 33318 28704 33324 28756
rect 33376 28744 33382 28756
rect 33413 28747 33471 28753
rect 33413 28744 33425 28747
rect 33376 28716 33425 28744
rect 33376 28704 33382 28716
rect 33413 28713 33425 28716
rect 33459 28713 33471 28747
rect 33413 28707 33471 28713
rect 2593 28543 2651 28549
rect 2593 28509 2605 28543
rect 2639 28540 2651 28543
rect 2958 28540 2964 28552
rect 2639 28512 2964 28540
rect 2639 28509 2651 28512
rect 2593 28503 2651 28509
rect 2958 28500 2964 28512
rect 3016 28500 3022 28552
rect 4157 28543 4215 28549
rect 4157 28509 4169 28543
rect 4203 28540 4215 28543
rect 4890 28540 4896 28552
rect 4203 28512 4896 28540
rect 4203 28509 4215 28512
rect 4157 28503 4215 28509
rect 4890 28500 4896 28512
rect 4948 28500 4954 28552
rect 15654 28500 15660 28552
rect 15712 28540 15718 28552
rect 16298 28540 16304 28552
rect 15712 28512 16304 28540
rect 15712 28500 15718 28512
rect 16298 28500 16304 28512
rect 16356 28500 16362 28552
rect 19058 28500 19064 28552
rect 19116 28540 19122 28552
rect 19613 28543 19671 28549
rect 19613 28540 19625 28543
rect 19116 28512 19625 28540
rect 19116 28500 19122 28512
rect 19613 28509 19625 28512
rect 19659 28509 19671 28543
rect 33318 28540 33324 28552
rect 33279 28512 33324 28540
rect 19613 28503 19671 28509
rect 33318 28500 33324 28512
rect 33376 28500 33382 28552
rect 34149 28543 34207 28549
rect 34149 28509 34161 28543
rect 34195 28540 34207 28543
rect 35434 28540 35440 28552
rect 34195 28512 35440 28540
rect 34195 28509 34207 28512
rect 34149 28503 34207 28509
rect 35434 28500 35440 28512
rect 35492 28500 35498 28552
rect 2317 28475 2375 28481
rect 2317 28441 2329 28475
rect 2363 28472 2375 28475
rect 2498 28472 2504 28484
rect 2363 28444 2504 28472
rect 2363 28441 2375 28444
rect 2317 28435 2375 28441
rect 2498 28432 2504 28444
rect 2556 28432 2562 28484
rect 16485 28407 16543 28413
rect 16485 28373 16497 28407
rect 16531 28404 16543 28407
rect 17678 28404 17684 28416
rect 16531 28376 17684 28404
rect 16531 28373 16543 28376
rect 16485 28367 16543 28373
rect 17678 28364 17684 28376
rect 17736 28364 17742 28416
rect 34054 28404 34060 28416
rect 34015 28376 34060 28404
rect 34054 28364 34060 28376
rect 34112 28364 34118 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 18690 28160 18696 28212
rect 18748 28200 18754 28212
rect 34054 28200 34060 28212
rect 18748 28172 34060 28200
rect 18748 28160 18754 28172
rect 34054 28160 34060 28172
rect 34112 28160 34118 28212
rect 1949 28067 2007 28073
rect 1949 28033 1961 28067
rect 1995 28064 2007 28067
rect 2222 28064 2228 28076
rect 1995 28036 2228 28064
rect 1995 28033 2007 28036
rect 1949 28027 2007 28033
rect 2222 28024 2228 28036
rect 2280 28064 2286 28076
rect 2593 28067 2651 28073
rect 2593 28064 2605 28067
rect 2280 28036 2605 28064
rect 2280 28024 2286 28036
rect 2593 28033 2605 28036
rect 2639 28064 2651 28067
rect 3513 28067 3571 28073
rect 3513 28064 3525 28067
rect 2639 28036 3525 28064
rect 2639 28033 2651 28036
rect 2593 28027 2651 28033
rect 3513 28033 3525 28036
rect 3559 28064 3571 28067
rect 4062 28064 4068 28076
rect 3559 28036 4068 28064
rect 3559 28033 3571 28036
rect 3513 28027 3571 28033
rect 4062 28024 4068 28036
rect 4120 28064 4126 28076
rect 4157 28067 4215 28073
rect 4157 28064 4169 28067
rect 4120 28036 4169 28064
rect 4120 28024 4126 28036
rect 4157 28033 4169 28036
rect 4203 28033 4215 28067
rect 4157 28027 4215 28033
rect 6638 28024 6644 28076
rect 6696 28064 6702 28076
rect 6733 28067 6791 28073
rect 6733 28064 6745 28067
rect 6696 28036 6745 28064
rect 6696 28024 6702 28036
rect 6733 28033 6745 28036
rect 6779 28033 6791 28067
rect 15838 28064 15844 28076
rect 15799 28036 15844 28064
rect 6733 28027 6791 28033
rect 15838 28024 15844 28036
rect 15896 28024 15902 28076
rect 16298 28024 16304 28076
rect 16356 28064 16362 28076
rect 16853 28067 16911 28073
rect 16853 28064 16865 28067
rect 16356 28036 16865 28064
rect 16356 28024 16362 28036
rect 16853 28033 16865 28036
rect 16899 28033 16911 28067
rect 33778 28064 33784 28076
rect 33739 28036 33784 28064
rect 16853 28027 16911 28033
rect 33778 28024 33784 28036
rect 33836 28024 33842 28076
rect 2038 27860 2044 27872
rect 1999 27832 2044 27860
rect 2038 27820 2044 27832
rect 2096 27820 2102 27872
rect 2682 27860 2688 27872
rect 2643 27832 2688 27860
rect 2682 27820 2688 27832
rect 2740 27820 2746 27872
rect 3605 27863 3663 27869
rect 3605 27829 3617 27863
rect 3651 27860 3663 27863
rect 3970 27860 3976 27872
rect 3651 27832 3976 27860
rect 3651 27829 3663 27832
rect 3605 27823 3663 27829
rect 3970 27820 3976 27832
rect 4028 27820 4034 27872
rect 4249 27863 4307 27869
rect 4249 27829 4261 27863
rect 4295 27860 4307 27863
rect 4982 27860 4988 27872
rect 4295 27832 4988 27860
rect 4295 27829 4307 27832
rect 4249 27823 4307 27829
rect 4982 27820 4988 27832
rect 5040 27820 5046 27872
rect 6825 27863 6883 27869
rect 6825 27829 6837 27863
rect 6871 27860 6883 27863
rect 7926 27860 7932 27872
rect 6871 27832 7932 27860
rect 6871 27829 6883 27832
rect 6825 27823 6883 27829
rect 7926 27820 7932 27832
rect 7984 27820 7990 27872
rect 15930 27820 15936 27872
rect 15988 27860 15994 27872
rect 16025 27863 16083 27869
rect 16025 27860 16037 27863
rect 15988 27832 16037 27860
rect 15988 27820 15994 27832
rect 16025 27829 16037 27832
rect 16071 27829 16083 27863
rect 16942 27860 16948 27872
rect 16903 27832 16948 27860
rect 16025 27823 16083 27829
rect 16942 27820 16948 27832
rect 17000 27820 17006 27872
rect 20714 27820 20720 27872
rect 20772 27860 20778 27872
rect 33689 27863 33747 27869
rect 33689 27860 33701 27863
rect 20772 27832 33701 27860
rect 20772 27820 20778 27832
rect 33689 27829 33701 27832
rect 33735 27829 33747 27863
rect 33689 27823 33747 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 16666 27588 16672 27600
rect 16627 27560 16672 27588
rect 16666 27548 16672 27560
rect 16724 27548 16730 27600
rect 17497 27591 17555 27597
rect 17497 27557 17509 27591
rect 17543 27557 17555 27591
rect 17497 27551 17555 27557
rect 2317 27523 2375 27529
rect 2317 27489 2329 27523
rect 2363 27520 2375 27523
rect 7098 27520 7104 27532
rect 2363 27492 7104 27520
rect 2363 27489 2375 27492
rect 2317 27483 2375 27489
rect 7098 27480 7104 27492
rect 7156 27480 7162 27532
rect 16853 27523 16911 27529
rect 16853 27489 16865 27523
rect 16899 27520 16911 27523
rect 17512 27520 17540 27551
rect 16899 27492 17540 27520
rect 16899 27489 16911 27492
rect 16853 27483 16911 27489
rect 1765 27455 1823 27461
rect 1765 27421 1777 27455
rect 1811 27452 1823 27455
rect 2222 27452 2228 27464
rect 1811 27424 2228 27452
rect 1811 27421 1823 27424
rect 1765 27415 1823 27421
rect 2222 27412 2228 27424
rect 2280 27412 2286 27464
rect 2409 27455 2467 27461
rect 2409 27452 2421 27455
rect 2332 27424 2421 27452
rect 2332 27396 2360 27424
rect 2409 27421 2421 27424
rect 2455 27421 2467 27455
rect 2409 27415 2467 27421
rect 3053 27455 3111 27461
rect 3053 27421 3065 27455
rect 3099 27421 3111 27455
rect 3053 27415 3111 27421
rect 2314 27344 2320 27396
rect 2372 27344 2378 27396
rect 3068 27384 3096 27415
rect 4062 27412 4068 27464
rect 4120 27452 4126 27464
rect 4157 27455 4215 27461
rect 4157 27452 4169 27455
rect 4120 27424 4169 27452
rect 4120 27412 4126 27424
rect 4157 27421 4169 27424
rect 4203 27452 4215 27455
rect 4617 27455 4675 27461
rect 4617 27452 4629 27455
rect 4203 27424 4629 27452
rect 4203 27421 4215 27424
rect 4157 27415 4215 27421
rect 4617 27421 4629 27424
rect 4663 27421 4675 27455
rect 4617 27415 4675 27421
rect 6733 27455 6791 27461
rect 6733 27421 6745 27455
rect 6779 27452 6791 27455
rect 6779 27424 7236 27452
rect 6779 27421 6791 27424
rect 6733 27415 6791 27421
rect 6822 27384 6828 27396
rect 3068 27356 6828 27384
rect 6822 27344 6828 27356
rect 6880 27344 6886 27396
rect 1673 27319 1731 27325
rect 1673 27285 1685 27319
rect 1719 27316 1731 27319
rect 1762 27316 1768 27328
rect 1719 27288 1768 27316
rect 1719 27285 1731 27288
rect 1673 27279 1731 27285
rect 1762 27276 1768 27288
rect 1820 27276 1826 27328
rect 2866 27316 2872 27328
rect 2827 27288 2872 27316
rect 2866 27276 2872 27288
rect 2924 27276 2930 27328
rect 3510 27276 3516 27328
rect 3568 27316 3574 27328
rect 4065 27319 4123 27325
rect 4065 27316 4077 27319
rect 3568 27288 4077 27316
rect 3568 27276 3574 27288
rect 4065 27285 4077 27288
rect 4111 27285 4123 27319
rect 4065 27279 4123 27285
rect 4709 27319 4767 27325
rect 4709 27285 4721 27319
rect 4755 27316 4767 27319
rect 5626 27316 5632 27328
rect 4755 27288 5632 27316
rect 4755 27285 4767 27288
rect 4709 27279 4767 27285
rect 5626 27276 5632 27288
rect 5684 27276 5690 27328
rect 5902 27316 5908 27328
rect 5863 27288 5908 27316
rect 5902 27276 5908 27288
rect 5960 27276 5966 27328
rect 6086 27276 6092 27328
rect 6144 27316 6150 27328
rect 7208 27325 7236 27424
rect 7282 27412 7288 27464
rect 7340 27452 7346 27464
rect 7377 27455 7435 27461
rect 7377 27452 7389 27455
rect 7340 27424 7389 27452
rect 7340 27412 7346 27424
rect 7377 27421 7389 27424
rect 7423 27421 7435 27455
rect 9122 27452 9128 27464
rect 9083 27424 9128 27452
rect 7377 27415 7435 27421
rect 9122 27412 9128 27424
rect 9180 27412 9186 27464
rect 12618 27412 12624 27464
rect 12676 27452 12682 27464
rect 13265 27455 13323 27461
rect 13265 27452 13277 27455
rect 12676 27424 13277 27452
rect 12676 27412 12682 27424
rect 13265 27421 13277 27424
rect 13311 27421 13323 27455
rect 15930 27452 15936 27464
rect 15891 27424 15936 27452
rect 13265 27415 13323 27421
rect 15930 27412 15936 27424
rect 15988 27412 15994 27464
rect 17037 27455 17095 27461
rect 17037 27421 17049 27455
rect 17083 27421 17095 27455
rect 17678 27452 17684 27464
rect 17639 27424 17684 27452
rect 17037 27415 17095 27421
rect 17052 27384 17080 27415
rect 17678 27412 17684 27424
rect 17736 27412 17742 27464
rect 18141 27387 18199 27393
rect 18141 27384 18153 27387
rect 17052 27356 18153 27384
rect 18141 27353 18153 27356
rect 18187 27353 18199 27387
rect 18141 27347 18199 27353
rect 6549 27319 6607 27325
rect 6549 27316 6561 27319
rect 6144 27288 6561 27316
rect 6144 27276 6150 27288
rect 6549 27285 6561 27288
rect 6595 27285 6607 27319
rect 6549 27279 6607 27285
rect 7193 27319 7251 27325
rect 7193 27285 7205 27319
rect 7239 27285 7251 27319
rect 9214 27316 9220 27328
rect 9175 27288 9220 27316
rect 7193 27279 7251 27285
rect 9214 27276 9220 27288
rect 9272 27276 9278 27328
rect 12250 27276 12256 27328
rect 12308 27316 12314 27328
rect 13081 27319 13139 27325
rect 13081 27316 13093 27319
rect 12308 27288 13093 27316
rect 12308 27276 12314 27288
rect 13081 27285 13093 27288
rect 13127 27285 13139 27319
rect 15746 27316 15752 27328
rect 15707 27288 15752 27316
rect 13081 27279 13139 27285
rect 15746 27276 15752 27288
rect 15804 27276 15810 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 3602 27112 3608 27124
rect 3563 27084 3608 27112
rect 3602 27072 3608 27084
rect 3660 27072 3666 27124
rect 6270 27072 6276 27124
rect 6328 27112 6334 27124
rect 6917 27115 6975 27121
rect 6917 27112 6929 27115
rect 6328 27084 6929 27112
rect 6328 27072 6334 27084
rect 6917 27081 6929 27084
rect 6963 27081 6975 27115
rect 6917 27075 6975 27081
rect 16666 27072 16672 27124
rect 16724 27112 16730 27124
rect 16853 27115 16911 27121
rect 16853 27112 16865 27115
rect 16724 27084 16865 27112
rect 16724 27072 16730 27084
rect 16853 27081 16865 27084
rect 16899 27081 16911 27115
rect 16853 27075 16911 27081
rect 29825 27115 29883 27121
rect 29825 27081 29837 27115
rect 29871 27112 29883 27115
rect 33226 27112 33232 27124
rect 29871 27084 33232 27112
rect 29871 27081 29883 27084
rect 29825 27075 29883 27081
rect 33226 27072 33232 27084
rect 33284 27072 33290 27124
rect 4062 27004 4068 27056
rect 4120 27044 4126 27056
rect 4120 27016 4936 27044
rect 4120 27004 4126 27016
rect 14 26936 20 26988
rect 72 26976 78 26988
rect 1581 26979 1639 26985
rect 1581 26976 1593 26979
rect 72 26948 1593 26976
rect 72 26936 78 26948
rect 1581 26945 1593 26948
rect 1627 26945 1639 26979
rect 2498 26976 2504 26988
rect 2459 26948 2504 26976
rect 1581 26939 1639 26945
rect 2498 26936 2504 26948
rect 2556 26976 2562 26988
rect 2961 26979 3019 26985
rect 2961 26976 2973 26979
rect 2556 26948 2973 26976
rect 2556 26936 2562 26948
rect 2961 26945 2973 26948
rect 3007 26945 3019 26979
rect 3786 26976 3792 26988
rect 3747 26948 3792 26976
rect 2961 26939 3019 26945
rect 2976 26908 3004 26939
rect 3786 26936 3792 26948
rect 3844 26936 3850 26988
rect 4433 26979 4491 26985
rect 4433 26945 4445 26979
rect 4479 26976 4491 26979
rect 4798 26976 4804 26988
rect 4479 26948 4804 26976
rect 4479 26945 4491 26948
rect 4433 26939 4491 26945
rect 4798 26936 4804 26948
rect 4856 26936 4862 26988
rect 4908 26985 4936 27016
rect 4893 26979 4951 26985
rect 4893 26945 4905 26979
rect 4939 26945 4951 26979
rect 4893 26939 4951 26945
rect 7282 26936 7288 26988
rect 7340 26976 7346 26988
rect 8021 26979 8079 26985
rect 8021 26976 8033 26979
rect 7340 26948 8033 26976
rect 7340 26936 7346 26948
rect 8021 26945 8033 26948
rect 8067 26945 8079 26979
rect 8021 26939 8079 26945
rect 8665 26979 8723 26985
rect 8665 26945 8677 26979
rect 8711 26976 8723 26979
rect 9030 26976 9036 26988
rect 8711 26948 9036 26976
rect 8711 26945 8723 26948
rect 8665 26939 8723 26945
rect 9030 26936 9036 26948
rect 9088 26936 9094 26988
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26945 11759 26979
rect 12618 26976 12624 26988
rect 12579 26948 12624 26976
rect 11701 26939 11759 26945
rect 5442 26908 5448 26920
rect 2976 26880 5448 26908
rect 5442 26868 5448 26880
rect 5500 26868 5506 26920
rect 7377 26911 7435 26917
rect 7377 26877 7389 26911
rect 7423 26877 7435 26911
rect 7377 26871 7435 26877
rect 7561 26911 7619 26917
rect 7561 26877 7573 26911
rect 7607 26908 7619 26911
rect 7650 26908 7656 26920
rect 7607 26880 7656 26908
rect 7607 26877 7619 26880
rect 7561 26871 7619 26877
rect 7392 26840 7420 26871
rect 7650 26868 7656 26880
rect 7708 26868 7714 26920
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 11716 26908 11744 26939
rect 12618 26936 12624 26948
rect 12676 26936 12682 26988
rect 13357 26979 13415 26985
rect 13357 26945 13369 26979
rect 13403 26945 13415 26979
rect 13357 26939 13415 26945
rect 14001 26979 14059 26985
rect 14001 26945 14013 26979
rect 14047 26945 14059 26979
rect 14001 26939 14059 26945
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26976 14887 26979
rect 16301 26979 16359 26985
rect 16301 26976 16313 26979
rect 14875 26948 16313 26976
rect 14875 26945 14887 26948
rect 14829 26939 14887 26945
rect 16301 26945 16313 26948
rect 16347 26945 16359 26979
rect 16301 26939 16359 26945
rect 13372 26908 13400 26939
rect 8628 26880 11744 26908
rect 11900 26880 13400 26908
rect 8628 26868 8634 26880
rect 11900 26849 11928 26880
rect 8113 26843 8171 26849
rect 8113 26840 8125 26843
rect 7392 26812 8125 26840
rect 8113 26809 8125 26812
rect 8159 26809 8171 26843
rect 8113 26803 8171 26809
rect 11885 26843 11943 26849
rect 11885 26809 11897 26843
rect 11931 26809 11943 26843
rect 11885 26803 11943 26809
rect 12434 26800 12440 26852
rect 12492 26840 12498 26852
rect 14016 26840 14044 26939
rect 15470 26908 15476 26920
rect 15431 26880 15476 26908
rect 15470 26868 15476 26880
rect 15528 26868 15534 26920
rect 16316 26908 16344 26939
rect 16942 26936 16948 26988
rect 17000 26976 17006 26988
rect 17313 26979 17371 26985
rect 17313 26976 17325 26979
rect 17000 26948 17325 26976
rect 17000 26936 17006 26948
rect 17313 26945 17325 26948
rect 17359 26945 17371 26979
rect 17313 26939 17371 26945
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26945 18475 26979
rect 18417 26939 18475 26945
rect 19061 26979 19119 26985
rect 19061 26945 19073 26979
rect 19107 26976 19119 26979
rect 20070 26976 20076 26988
rect 19107 26948 20076 26976
rect 19107 26945 19119 26948
rect 19061 26939 19119 26945
rect 17218 26908 17224 26920
rect 16316 26880 17224 26908
rect 17218 26868 17224 26880
rect 17276 26868 17282 26920
rect 17497 26911 17555 26917
rect 17497 26877 17509 26911
rect 17543 26908 17555 26911
rect 18138 26908 18144 26920
rect 17543 26880 18144 26908
rect 17543 26877 17555 26880
rect 17497 26871 17555 26877
rect 18138 26868 18144 26880
rect 18196 26868 18202 26920
rect 18432 26908 18460 26939
rect 20070 26936 20076 26948
rect 20128 26936 20134 26988
rect 29730 26976 29736 26988
rect 29691 26948 29736 26976
rect 29730 26936 29736 26948
rect 29788 26936 29794 26988
rect 35342 26936 35348 26988
rect 35400 26976 35406 26988
rect 38013 26979 38071 26985
rect 38013 26976 38025 26979
rect 35400 26948 38025 26976
rect 35400 26936 35406 26948
rect 38013 26945 38025 26948
rect 38059 26945 38071 26979
rect 38013 26939 38071 26945
rect 19426 26908 19432 26920
rect 18432 26880 19432 26908
rect 19426 26868 19432 26880
rect 19484 26868 19490 26920
rect 12492 26812 14044 26840
rect 12492 26800 12498 26812
rect 1765 26775 1823 26781
rect 1765 26741 1777 26775
rect 1811 26772 1823 26775
rect 1854 26772 1860 26784
rect 1811 26744 1860 26772
rect 1811 26741 1823 26744
rect 1765 26735 1823 26741
rect 1854 26732 1860 26744
rect 1912 26732 1918 26784
rect 2409 26775 2467 26781
rect 2409 26741 2421 26775
rect 2455 26772 2467 26775
rect 2498 26772 2504 26784
rect 2455 26744 2504 26772
rect 2455 26741 2467 26744
rect 2409 26735 2467 26741
rect 2498 26732 2504 26744
rect 2556 26732 2562 26784
rect 3053 26775 3111 26781
rect 3053 26741 3065 26775
rect 3099 26772 3111 26775
rect 3142 26772 3148 26784
rect 3099 26744 3148 26772
rect 3099 26741 3111 26744
rect 3053 26735 3111 26741
rect 3142 26732 3148 26744
rect 3200 26732 3206 26784
rect 4249 26775 4307 26781
rect 4249 26741 4261 26775
rect 4295 26772 4307 26775
rect 4706 26772 4712 26784
rect 4295 26744 4712 26772
rect 4295 26741 4307 26744
rect 4249 26735 4307 26741
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 4985 26775 5043 26781
rect 4985 26741 4997 26775
rect 5031 26772 5043 26775
rect 5074 26772 5080 26784
rect 5031 26744 5080 26772
rect 5031 26741 5043 26744
rect 4985 26735 5043 26741
rect 5074 26732 5080 26744
rect 5132 26732 5138 26784
rect 8849 26775 8907 26781
rect 8849 26741 8861 26775
rect 8895 26772 8907 26775
rect 9950 26772 9956 26784
rect 8895 26744 9956 26772
rect 8895 26741 8907 26744
rect 8849 26735 8907 26741
rect 9950 26732 9956 26744
rect 10008 26732 10014 26784
rect 12713 26775 12771 26781
rect 12713 26741 12725 26775
rect 12759 26772 12771 26775
rect 13354 26772 13360 26784
rect 12759 26744 13360 26772
rect 12759 26741 12771 26744
rect 12713 26735 12771 26741
rect 13354 26732 13360 26744
rect 13412 26732 13418 26784
rect 13541 26775 13599 26781
rect 13541 26741 13553 26775
rect 13587 26772 13599 26775
rect 13630 26772 13636 26784
rect 13587 26744 13636 26772
rect 13587 26741 13599 26744
rect 13541 26735 13599 26741
rect 13630 26732 13636 26744
rect 13688 26732 13694 26784
rect 14185 26775 14243 26781
rect 14185 26741 14197 26775
rect 14231 26772 14243 26775
rect 14826 26772 14832 26784
rect 14231 26744 14832 26772
rect 14231 26741 14243 26744
rect 14185 26735 14243 26741
rect 14826 26732 14832 26744
rect 14884 26732 14890 26784
rect 14921 26775 14979 26781
rect 14921 26741 14933 26775
rect 14967 26772 14979 26775
rect 15194 26772 15200 26784
rect 14967 26744 15200 26772
rect 14967 26741 14979 26744
rect 14921 26735 14979 26741
rect 15194 26732 15200 26744
rect 15252 26732 15258 26784
rect 15562 26732 15568 26784
rect 15620 26772 15626 26784
rect 16117 26775 16175 26781
rect 16117 26772 16129 26775
rect 15620 26744 16129 26772
rect 15620 26732 15626 26744
rect 16117 26741 16129 26744
rect 16163 26741 16175 26775
rect 16117 26735 16175 26741
rect 17678 26732 17684 26784
rect 17736 26772 17742 26784
rect 18233 26775 18291 26781
rect 18233 26772 18245 26775
rect 17736 26744 18245 26772
rect 17736 26732 17742 26744
rect 18233 26741 18245 26744
rect 18279 26741 18291 26775
rect 18874 26772 18880 26784
rect 18835 26744 18880 26772
rect 18233 26735 18291 26741
rect 18874 26732 18880 26744
rect 18932 26732 18938 26784
rect 38194 26772 38200 26784
rect 38155 26744 38200 26772
rect 38194 26732 38200 26744
rect 38252 26732 38258 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 4798 26528 4804 26580
rect 4856 26568 4862 26580
rect 4985 26571 5043 26577
rect 4985 26568 4997 26571
rect 4856 26540 4997 26568
rect 4856 26528 4862 26540
rect 4985 26537 4997 26540
rect 5031 26537 5043 26571
rect 6270 26568 6276 26580
rect 6231 26540 6276 26568
rect 4985 26531 5043 26537
rect 6270 26528 6276 26540
rect 6328 26528 6334 26580
rect 17037 26571 17095 26577
rect 17037 26537 17049 26571
rect 17083 26568 17095 26571
rect 18138 26568 18144 26580
rect 17083 26540 18000 26568
rect 18099 26540 18144 26568
rect 17083 26537 17095 26540
rect 17037 26531 17095 26537
rect 8202 26460 8208 26512
rect 8260 26500 8266 26512
rect 12437 26503 12495 26509
rect 8260 26472 9628 26500
rect 8260 26460 8266 26472
rect 5902 26432 5908 26444
rect 5863 26404 5908 26432
rect 5902 26392 5908 26404
rect 5960 26392 5966 26444
rect 6086 26432 6092 26444
rect 6047 26404 6092 26432
rect 6086 26392 6092 26404
rect 6144 26392 6150 26444
rect 8021 26435 8079 26441
rect 8021 26401 8033 26435
rect 8067 26432 8079 26435
rect 9217 26435 9275 26441
rect 9217 26432 9229 26435
rect 8067 26404 9229 26432
rect 8067 26401 8079 26404
rect 8021 26395 8079 26401
rect 9217 26401 9229 26404
rect 9263 26401 9275 26435
rect 9600 26432 9628 26472
rect 12437 26469 12449 26503
rect 12483 26500 12495 26503
rect 13538 26500 13544 26512
rect 12483 26472 13544 26500
rect 12483 26469 12495 26472
rect 12437 26463 12495 26469
rect 13538 26460 13544 26472
rect 13596 26460 13602 26512
rect 17497 26503 17555 26509
rect 17497 26469 17509 26503
rect 17543 26500 17555 26503
rect 17586 26500 17592 26512
rect 17543 26472 17592 26500
rect 17543 26469 17555 26472
rect 17497 26463 17555 26469
rect 17586 26460 17592 26472
rect 17644 26460 17650 26512
rect 17972 26500 18000 26540
rect 18138 26528 18144 26540
rect 18196 26528 18202 26580
rect 20438 26568 20444 26580
rect 18708 26540 20444 26568
rect 18708 26500 18736 26540
rect 20438 26528 20444 26540
rect 20496 26528 20502 26580
rect 36265 26571 36323 26577
rect 36265 26537 36277 26571
rect 36311 26568 36323 26571
rect 38010 26568 38016 26580
rect 36311 26540 38016 26568
rect 36311 26537 36323 26540
rect 36265 26531 36323 26537
rect 38010 26528 38016 26540
rect 38068 26528 38074 26580
rect 17972 26472 18736 26500
rect 14274 26432 14280 26444
rect 9600 26404 14280 26432
rect 9217 26395 9275 26401
rect 14274 26392 14280 26404
rect 14332 26392 14338 26444
rect 14458 26392 14464 26444
rect 14516 26432 14522 26444
rect 14516 26404 16896 26432
rect 14516 26392 14522 26404
rect 2314 26364 2320 26376
rect 2275 26336 2320 26364
rect 2314 26324 2320 26336
rect 2372 26324 2378 26376
rect 2777 26367 2835 26373
rect 2777 26333 2789 26367
rect 2823 26364 2835 26367
rect 2958 26364 2964 26376
rect 2823 26336 2964 26364
rect 2823 26333 2835 26336
rect 2777 26327 2835 26333
rect 2958 26324 2964 26336
rect 3016 26324 3022 26376
rect 4525 26367 4583 26373
rect 4525 26333 4537 26367
rect 4571 26333 4583 26367
rect 4525 26327 4583 26333
rect 1946 26256 1952 26308
rect 2004 26296 2010 26308
rect 2225 26299 2283 26305
rect 2225 26296 2237 26299
rect 2004 26268 2237 26296
rect 2004 26256 2010 26268
rect 2225 26265 2237 26268
rect 2271 26265 2283 26299
rect 2225 26259 2283 26265
rect 2869 26299 2927 26305
rect 2869 26265 2881 26299
rect 2915 26296 2927 26299
rect 4062 26296 4068 26308
rect 2915 26268 4068 26296
rect 2915 26265 2927 26268
rect 2869 26259 2927 26265
rect 4062 26256 4068 26268
rect 4120 26256 4126 26308
rect 4540 26296 4568 26327
rect 4798 26324 4804 26376
rect 4856 26364 4862 26376
rect 5169 26367 5227 26373
rect 5169 26364 5181 26367
rect 4856 26336 5181 26364
rect 4856 26324 4862 26336
rect 5169 26333 5181 26336
rect 5215 26333 5227 26367
rect 8202 26364 8208 26376
rect 8163 26336 8208 26364
rect 5169 26327 5227 26333
rect 8202 26324 8208 26336
rect 8260 26324 8266 26376
rect 9030 26324 9036 26376
rect 9088 26364 9094 26376
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 9088 26336 9137 26364
rect 9088 26324 9094 26336
rect 9125 26333 9137 26336
rect 9171 26333 9183 26367
rect 9950 26364 9956 26376
rect 9911 26336 9956 26364
rect 9125 26327 9183 26333
rect 9950 26324 9956 26336
rect 10008 26324 10014 26376
rect 10962 26364 10968 26376
rect 10923 26336 10968 26364
rect 10962 26324 10968 26336
rect 11020 26324 11026 26376
rect 11609 26367 11667 26373
rect 11609 26333 11621 26367
rect 11655 26364 11667 26367
rect 12066 26364 12072 26376
rect 11655 26336 12072 26364
rect 11655 26333 11667 26336
rect 11609 26327 11667 26333
rect 12066 26324 12072 26336
rect 12124 26324 12130 26376
rect 12250 26364 12256 26376
rect 12211 26336 12256 26364
rect 12250 26324 12256 26336
rect 12308 26324 12314 26376
rect 12526 26324 12532 26376
rect 12584 26364 12590 26376
rect 13081 26367 13139 26373
rect 13081 26364 13093 26367
rect 12584 26336 13093 26364
rect 12584 26324 12590 26336
rect 13081 26333 13093 26336
rect 13127 26333 13139 26367
rect 13081 26327 13139 26333
rect 13541 26367 13599 26373
rect 13541 26333 13553 26367
rect 13587 26364 13599 26367
rect 14369 26367 14427 26373
rect 14369 26364 14381 26367
rect 13587 26336 14381 26364
rect 13587 26333 13599 26336
rect 13541 26327 13599 26333
rect 14369 26333 14381 26336
rect 14415 26333 14427 26367
rect 15562 26364 15568 26376
rect 15523 26336 15568 26364
rect 14369 26327 14427 26333
rect 11054 26296 11060 26308
rect 4540 26268 5212 26296
rect 11015 26268 11060 26296
rect 5184 26240 5212 26268
rect 11054 26256 11060 26268
rect 11112 26256 11118 26308
rect 11701 26299 11759 26305
rect 11701 26265 11713 26299
rect 11747 26296 11759 26299
rect 11882 26296 11888 26308
rect 11747 26268 11888 26296
rect 11747 26265 11759 26268
rect 11701 26259 11759 26265
rect 11882 26256 11888 26268
rect 11940 26256 11946 26308
rect 12894 26256 12900 26308
rect 12952 26296 12958 26308
rect 13556 26296 13584 26327
rect 15562 26324 15568 26336
rect 15620 26324 15626 26376
rect 16868 26373 16896 26404
rect 17218 26392 17224 26444
rect 17276 26432 17282 26444
rect 17276 26404 18736 26432
rect 17276 26392 17282 26404
rect 16853 26367 16911 26373
rect 16853 26333 16865 26367
rect 16899 26333 16911 26367
rect 17678 26364 17684 26376
rect 17639 26336 17684 26364
rect 16853 26327 16911 26333
rect 17678 26324 17684 26336
rect 17736 26324 17742 26376
rect 18601 26367 18659 26373
rect 18601 26333 18613 26367
rect 18647 26333 18659 26367
rect 18708 26364 18736 26404
rect 18782 26392 18788 26444
rect 18840 26432 18846 26444
rect 18840 26404 18885 26432
rect 18840 26392 18846 26404
rect 19429 26367 19487 26373
rect 19429 26364 19441 26367
rect 18708 26336 19441 26364
rect 18601 26327 18659 26333
rect 19429 26333 19441 26336
rect 19475 26333 19487 26367
rect 36078 26364 36084 26376
rect 36039 26336 36084 26364
rect 19429 26327 19487 26333
rect 12952 26268 13584 26296
rect 14461 26299 14519 26305
rect 12952 26256 12958 26268
rect 14461 26265 14473 26299
rect 14507 26296 14519 26299
rect 15102 26296 15108 26308
rect 14507 26268 15108 26296
rect 14507 26265 14519 26268
rect 14461 26259 14519 26265
rect 15102 26256 15108 26268
rect 15160 26256 15166 26308
rect 18616 26296 18644 26327
rect 36078 26324 36084 26336
rect 36136 26324 36142 26376
rect 20622 26296 20628 26308
rect 18616 26268 20628 26296
rect 20622 26256 20628 26268
rect 20680 26256 20686 26308
rect 4338 26228 4344 26240
rect 4299 26200 4344 26228
rect 4338 26188 4344 26200
rect 4396 26188 4402 26240
rect 5166 26188 5172 26240
rect 5224 26188 5230 26240
rect 7561 26231 7619 26237
rect 7561 26197 7573 26231
rect 7607 26228 7619 26231
rect 7650 26228 7656 26240
rect 7607 26200 7656 26228
rect 7607 26197 7619 26200
rect 7561 26191 7619 26197
rect 7650 26188 7656 26200
rect 7708 26188 7714 26240
rect 9766 26228 9772 26240
rect 9727 26200 9772 26228
rect 9766 26188 9772 26200
rect 9824 26188 9830 26240
rect 12710 26188 12716 26240
rect 12768 26228 12774 26240
rect 12989 26231 13047 26237
rect 12989 26228 13001 26231
rect 12768 26200 13001 26228
rect 12768 26188 12774 26200
rect 12989 26197 13001 26200
rect 13035 26197 13047 26231
rect 13722 26228 13728 26240
rect 13683 26200 13728 26228
rect 12989 26191 13047 26197
rect 13722 26188 13728 26200
rect 13780 26188 13786 26240
rect 15749 26231 15807 26237
rect 15749 26197 15761 26231
rect 15795 26228 15807 26231
rect 16022 26228 16028 26240
rect 15795 26200 16028 26228
rect 15795 26197 15807 26200
rect 15749 26191 15807 26197
rect 16022 26188 16028 26200
rect 16080 26188 16086 26240
rect 16206 26228 16212 26240
rect 16167 26200 16212 26228
rect 16206 26188 16212 26200
rect 16264 26188 16270 26240
rect 19334 26188 19340 26240
rect 19392 26228 19398 26240
rect 19521 26231 19579 26237
rect 19521 26228 19533 26231
rect 19392 26200 19533 26228
rect 19392 26188 19398 26200
rect 19521 26197 19533 26200
rect 19567 26197 19579 26231
rect 19521 26191 19579 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 3786 26024 3792 26036
rect 3747 25996 3792 26024
rect 3786 25984 3792 25996
rect 3844 25984 3850 26036
rect 7650 26024 7656 26036
rect 7611 25996 7656 26024
rect 7650 25984 7656 25996
rect 7708 25984 7714 26036
rect 11885 26027 11943 26033
rect 11885 25993 11897 26027
rect 11931 26024 11943 26027
rect 12342 26024 12348 26036
rect 11931 25996 12348 26024
rect 11931 25993 11943 25996
rect 11885 25987 11943 25993
rect 12342 25984 12348 25996
rect 12400 25984 12406 26036
rect 15838 26024 15844 26036
rect 12728 25996 15844 26024
rect 4338 25956 4344 25968
rect 3252 25928 4344 25956
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 2222 25848 2228 25900
rect 2280 25888 2286 25900
rect 3252 25897 3280 25928
rect 4338 25916 4344 25928
rect 4396 25916 4402 25968
rect 4448 25928 6776 25956
rect 2409 25891 2467 25897
rect 2409 25888 2421 25891
rect 2280 25860 2421 25888
rect 2280 25848 2286 25860
rect 2409 25857 2421 25860
rect 2455 25857 2467 25891
rect 2409 25851 2467 25857
rect 3237 25891 3295 25897
rect 3237 25857 3249 25891
rect 3283 25857 3295 25891
rect 3237 25851 3295 25857
rect 3881 25891 3939 25897
rect 3881 25857 3893 25891
rect 3927 25888 3939 25891
rect 4448 25888 4476 25928
rect 3927 25860 4476 25888
rect 4525 25891 4583 25897
rect 3927 25857 3939 25860
rect 3881 25851 3939 25857
rect 4525 25857 4537 25891
rect 4571 25888 4583 25891
rect 4798 25888 4804 25900
rect 4571 25860 4804 25888
rect 4571 25857 4583 25860
rect 4525 25851 4583 25857
rect 4798 25848 4804 25860
rect 4856 25848 4862 25900
rect 5169 25891 5227 25897
rect 5169 25857 5181 25891
rect 5215 25888 5227 25891
rect 5997 25891 6055 25897
rect 5215 25860 5856 25888
rect 5215 25857 5227 25860
rect 5169 25851 5227 25857
rect 1302 25712 1308 25764
rect 1360 25752 1366 25764
rect 5828 25761 5856 25860
rect 5997 25857 6009 25891
rect 6043 25857 6055 25891
rect 6748 25888 6776 25928
rect 6822 25916 6828 25968
rect 6880 25956 6886 25968
rect 9033 25959 9091 25965
rect 9033 25956 9045 25959
rect 6880 25928 9045 25956
rect 6880 25916 6886 25928
rect 9033 25925 9045 25928
rect 9079 25925 9091 25959
rect 12434 25956 12440 25968
rect 9033 25919 9091 25925
rect 9140 25928 12440 25956
rect 7006 25888 7012 25900
rect 6748 25860 7012 25888
rect 5997 25851 6055 25857
rect 6012 25820 6040 25851
rect 7006 25848 7012 25860
rect 7064 25848 7070 25900
rect 7193 25891 7251 25897
rect 7193 25857 7205 25891
rect 7239 25888 7251 25891
rect 7374 25888 7380 25900
rect 7239 25860 7380 25888
rect 7239 25857 7251 25860
rect 7193 25851 7251 25857
rect 7374 25848 7380 25860
rect 7432 25848 7438 25900
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25888 8355 25891
rect 8386 25888 8392 25900
rect 8343 25860 8392 25888
rect 8343 25857 8355 25860
rect 8297 25851 8355 25857
rect 8386 25848 8392 25860
rect 8444 25848 8450 25900
rect 9140 25897 9168 25928
rect 12434 25916 12440 25928
rect 12492 25916 12498 25968
rect 9125 25891 9183 25897
rect 9125 25857 9137 25891
rect 9171 25857 9183 25891
rect 10226 25888 10232 25900
rect 10187 25860 10232 25888
rect 9125 25851 9183 25857
rect 10226 25848 10232 25860
rect 10284 25848 10290 25900
rect 10318 25848 10324 25900
rect 10376 25888 10382 25900
rect 10962 25888 10968 25900
rect 10376 25860 10968 25888
rect 10376 25848 10382 25860
rect 10962 25848 10968 25860
rect 11020 25888 11026 25900
rect 11149 25891 11207 25897
rect 11149 25888 11161 25891
rect 11020 25860 11161 25888
rect 11020 25848 11026 25860
rect 11149 25857 11161 25860
rect 11195 25857 11207 25891
rect 11149 25851 11207 25857
rect 6822 25820 6828 25832
rect 6012 25792 6828 25820
rect 6822 25780 6828 25792
rect 6880 25780 6886 25832
rect 8113 25823 8171 25829
rect 8113 25789 8125 25823
rect 8159 25820 8171 25823
rect 9766 25820 9772 25832
rect 8159 25792 9772 25820
rect 8159 25789 8171 25792
rect 8113 25783 8171 25789
rect 9766 25780 9772 25792
rect 9824 25780 9830 25832
rect 10042 25820 10048 25832
rect 10003 25792 10048 25820
rect 10042 25780 10048 25792
rect 10100 25780 10106 25832
rect 11164 25820 11192 25851
rect 11606 25848 11612 25900
rect 11664 25888 11670 25900
rect 11701 25891 11759 25897
rect 11701 25888 11713 25891
rect 11664 25860 11713 25888
rect 11664 25848 11670 25860
rect 11701 25857 11713 25860
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25888 12587 25891
rect 12618 25888 12624 25900
rect 12575 25860 12624 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 12618 25848 12624 25860
rect 12676 25848 12682 25900
rect 12728 25820 12756 25996
rect 13722 25916 13728 25968
rect 13780 25956 13786 25968
rect 13780 25928 14596 25956
rect 13780 25916 13786 25928
rect 13170 25888 13176 25900
rect 13131 25860 13176 25888
rect 13170 25848 13176 25860
rect 13228 25848 13234 25900
rect 14568 25897 14596 25928
rect 15488 25897 15516 25996
rect 15838 25984 15844 25996
rect 15896 25984 15902 26036
rect 19426 26024 19432 26036
rect 19306 25996 19432 26024
rect 19306 25956 19334 25996
rect 19426 25984 19432 25996
rect 19484 25984 19490 26036
rect 20070 26024 20076 26036
rect 20031 25996 20076 26024
rect 20070 25984 20076 25996
rect 20128 25984 20134 26036
rect 20622 25984 20628 26036
rect 20680 26024 20686 26036
rect 20809 26027 20867 26033
rect 20809 26024 20821 26027
rect 20680 25996 20821 26024
rect 20680 25984 20686 25996
rect 20809 25993 20821 25996
rect 20855 25993 20867 26027
rect 20809 25987 20867 25993
rect 29641 26027 29699 26033
rect 29641 25993 29653 26027
rect 29687 26024 29699 26027
rect 33870 26024 33876 26036
rect 29687 25996 33876 26024
rect 29687 25993 29699 25996
rect 29641 25987 29699 25993
rect 33870 25984 33876 25996
rect 33928 25984 33934 26036
rect 16132 25928 19334 25956
rect 14093 25891 14151 25897
rect 14093 25857 14105 25891
rect 14139 25857 14151 25891
rect 14093 25851 14151 25857
rect 14553 25891 14611 25897
rect 14553 25857 14565 25891
rect 14599 25857 14611 25891
rect 14553 25851 14611 25857
rect 15473 25891 15531 25897
rect 15473 25857 15485 25891
rect 15519 25857 15531 25891
rect 15473 25851 15531 25857
rect 11164 25792 12756 25820
rect 12802 25780 12808 25832
rect 12860 25820 12866 25832
rect 14108 25820 14136 25851
rect 15930 25848 15936 25900
rect 15988 25888 15994 25900
rect 16132 25897 16160 25928
rect 16117 25891 16175 25897
rect 16117 25888 16129 25891
rect 15988 25860 16129 25888
rect 15988 25848 15994 25860
rect 16117 25857 16129 25860
rect 16163 25857 16175 25891
rect 17494 25888 17500 25900
rect 17455 25860 17500 25888
rect 16117 25851 16175 25857
rect 17494 25848 17500 25860
rect 17552 25848 17558 25900
rect 18509 25891 18567 25897
rect 18509 25857 18521 25891
rect 18555 25888 18567 25891
rect 19334 25888 19340 25900
rect 18555 25860 19340 25888
rect 18555 25857 18567 25860
rect 18509 25851 18567 25857
rect 19334 25848 19340 25860
rect 19392 25848 19398 25900
rect 19429 25889 19487 25895
rect 19429 25855 19441 25889
rect 19475 25855 19487 25889
rect 20257 25891 20315 25897
rect 20257 25888 20269 25891
rect 19429 25849 19487 25855
rect 19812 25860 20269 25888
rect 12860 25792 14136 25820
rect 15565 25823 15623 25829
rect 12860 25780 12866 25792
rect 15565 25789 15577 25823
rect 15611 25820 15623 25823
rect 17313 25823 17371 25829
rect 17313 25820 17325 25823
rect 15611 25792 17325 25820
rect 15611 25789 15623 25792
rect 15565 25783 15623 25789
rect 17313 25789 17325 25792
rect 17359 25789 17371 25823
rect 18690 25820 18696 25832
rect 18651 25792 18696 25820
rect 17313 25783 17371 25789
rect 18690 25780 18696 25792
rect 18748 25780 18754 25832
rect 19444 25820 19472 25849
rect 19518 25820 19524 25832
rect 19444 25792 19524 25820
rect 19518 25780 19524 25792
rect 19576 25780 19582 25832
rect 2501 25755 2559 25761
rect 2501 25752 2513 25755
rect 1360 25724 2513 25752
rect 1360 25712 1366 25724
rect 2501 25721 2513 25724
rect 2547 25721 2559 25755
rect 2501 25715 2559 25721
rect 5813 25755 5871 25761
rect 5813 25721 5825 25755
rect 5859 25721 5871 25755
rect 5813 25715 5871 25721
rect 5902 25712 5908 25764
rect 5960 25752 5966 25764
rect 5960 25724 11100 25752
rect 5960 25712 5966 25724
rect 1765 25687 1823 25693
rect 1765 25653 1777 25687
rect 1811 25684 1823 25687
rect 1854 25684 1860 25696
rect 1811 25656 1860 25684
rect 1811 25653 1823 25656
rect 1765 25647 1823 25653
rect 1854 25644 1860 25656
rect 1912 25644 1918 25696
rect 3053 25687 3111 25693
rect 3053 25653 3065 25687
rect 3099 25684 3111 25687
rect 3234 25684 3240 25696
rect 3099 25656 3240 25684
rect 3099 25653 3111 25656
rect 3053 25647 3111 25653
rect 3234 25644 3240 25656
rect 3292 25644 3298 25696
rect 4433 25687 4491 25693
rect 4433 25653 4445 25687
rect 4479 25684 4491 25687
rect 4614 25684 4620 25696
rect 4479 25656 4620 25684
rect 4479 25653 4491 25656
rect 4433 25647 4491 25653
rect 4614 25644 4620 25656
rect 4672 25644 4678 25696
rect 5353 25687 5411 25693
rect 5353 25653 5365 25687
rect 5399 25684 5411 25687
rect 5534 25684 5540 25696
rect 5399 25656 5540 25684
rect 5399 25653 5411 25656
rect 5353 25647 5411 25653
rect 5534 25644 5540 25656
rect 5592 25644 5598 25696
rect 6454 25644 6460 25696
rect 6512 25684 6518 25696
rect 7009 25687 7067 25693
rect 7009 25684 7021 25687
rect 6512 25656 7021 25684
rect 6512 25644 6518 25656
rect 7009 25653 7021 25656
rect 7055 25653 7067 25687
rect 7009 25647 7067 25653
rect 8662 25644 8668 25696
rect 8720 25684 8726 25696
rect 9585 25687 9643 25693
rect 9585 25684 9597 25687
rect 8720 25656 9597 25684
rect 8720 25644 8726 25656
rect 9585 25653 9597 25656
rect 9631 25653 9643 25687
rect 9585 25647 9643 25653
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 10965 25687 11023 25693
rect 10965 25684 10977 25687
rect 9732 25656 10977 25684
rect 9732 25644 9738 25656
rect 10965 25653 10977 25656
rect 11011 25653 11023 25687
rect 11072 25684 11100 25724
rect 11698 25712 11704 25764
rect 11756 25752 11762 25764
rect 12989 25755 13047 25761
rect 12989 25752 13001 25755
rect 11756 25724 13001 25752
rect 11756 25712 11762 25724
rect 12989 25721 13001 25724
rect 13035 25721 13047 25755
rect 16390 25752 16396 25764
rect 12989 25715 13047 25721
rect 13096 25724 16396 25752
rect 11974 25684 11980 25696
rect 11072 25656 11980 25684
rect 10965 25647 11023 25653
rect 11974 25644 11980 25656
rect 12032 25644 12038 25696
rect 12342 25684 12348 25696
rect 12303 25656 12348 25684
rect 12342 25644 12348 25656
rect 12400 25644 12406 25696
rect 12434 25644 12440 25696
rect 12492 25684 12498 25696
rect 13096 25684 13124 25724
rect 16390 25712 16396 25724
rect 16448 25712 16454 25764
rect 16482 25712 16488 25764
rect 16540 25752 16546 25764
rect 19812 25752 19840 25860
rect 20257 25857 20269 25860
rect 20303 25888 20315 25891
rect 20717 25891 20775 25897
rect 20717 25888 20729 25891
rect 20303 25860 20729 25888
rect 20303 25857 20315 25860
rect 20257 25851 20315 25857
rect 20717 25857 20729 25860
rect 20763 25857 20775 25891
rect 20717 25851 20775 25857
rect 24026 25848 24032 25900
rect 24084 25888 24090 25900
rect 29549 25891 29607 25897
rect 29549 25888 29561 25891
rect 24084 25860 29561 25888
rect 24084 25848 24090 25860
rect 29549 25857 29561 25860
rect 29595 25857 29607 25891
rect 29549 25851 29607 25857
rect 16540 25724 19840 25752
rect 16540 25712 16546 25724
rect 12492 25656 13124 25684
rect 12492 25644 12498 25656
rect 13814 25644 13820 25696
rect 13872 25684 13878 25696
rect 13909 25687 13967 25693
rect 13909 25684 13921 25687
rect 13872 25656 13921 25684
rect 13872 25644 13878 25656
rect 13909 25653 13921 25656
rect 13955 25653 13967 25687
rect 14734 25684 14740 25696
rect 14695 25656 14740 25684
rect 13909 25647 13967 25653
rect 14734 25644 14740 25656
rect 14792 25644 14798 25696
rect 16209 25687 16267 25693
rect 16209 25653 16221 25687
rect 16255 25684 16267 25687
rect 16758 25684 16764 25696
rect 16255 25656 16764 25684
rect 16255 25653 16267 25656
rect 16209 25647 16267 25653
rect 16758 25644 16764 25656
rect 16816 25644 16822 25696
rect 16850 25644 16856 25696
rect 16908 25684 16914 25696
rect 18325 25687 18383 25693
rect 16908 25656 16953 25684
rect 16908 25644 16914 25656
rect 18325 25653 18337 25687
rect 18371 25684 18383 25687
rect 18506 25684 18512 25696
rect 18371 25656 18512 25684
rect 18371 25653 18383 25656
rect 18325 25647 18383 25653
rect 18506 25644 18512 25656
rect 18564 25644 18570 25696
rect 19521 25687 19579 25693
rect 19521 25653 19533 25687
rect 19567 25684 19579 25687
rect 20530 25684 20536 25696
rect 19567 25656 20536 25684
rect 19567 25653 19579 25656
rect 19521 25647 19579 25653
rect 20530 25644 20536 25656
rect 20588 25644 20594 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 8481 25483 8539 25489
rect 4120 25452 8432 25480
rect 4120 25440 4126 25452
rect 3237 25415 3295 25421
rect 3237 25381 3249 25415
rect 3283 25412 3295 25415
rect 8110 25412 8116 25424
rect 3283 25384 8116 25412
rect 3283 25381 3295 25384
rect 3237 25375 3295 25381
rect 8110 25372 8116 25384
rect 8168 25372 8174 25424
rect 8404 25412 8432 25452
rect 8481 25449 8493 25483
rect 8527 25480 8539 25483
rect 10042 25480 10048 25492
rect 8527 25452 10048 25480
rect 8527 25449 8539 25452
rect 8481 25443 8539 25449
rect 10042 25440 10048 25452
rect 10100 25440 10106 25492
rect 10410 25440 10416 25492
rect 10468 25480 10474 25492
rect 13170 25480 13176 25492
rect 10468 25452 13176 25480
rect 10468 25440 10474 25452
rect 13170 25440 13176 25452
rect 13228 25440 13234 25492
rect 14550 25480 14556 25492
rect 13556 25452 14556 25480
rect 9766 25412 9772 25424
rect 8404 25384 9772 25412
rect 9766 25372 9772 25384
rect 9824 25372 9830 25424
rect 13556 25412 13584 25452
rect 14550 25440 14556 25452
rect 14608 25440 14614 25492
rect 18138 25480 18144 25492
rect 18099 25452 18144 25480
rect 18138 25440 18144 25452
rect 18196 25440 18202 25492
rect 35713 25483 35771 25489
rect 35713 25449 35725 25483
rect 35759 25480 35771 25483
rect 36078 25480 36084 25492
rect 35759 25452 36084 25480
rect 35759 25449 35771 25452
rect 35713 25443 35771 25449
rect 36078 25440 36084 25452
rect 36136 25440 36142 25492
rect 15381 25415 15439 25421
rect 15381 25412 15393 25415
rect 10060 25384 13584 25412
rect 13648 25384 15393 25412
rect 2593 25347 2651 25353
rect 2593 25313 2605 25347
rect 2639 25344 2651 25347
rect 3694 25344 3700 25356
rect 2639 25316 3700 25344
rect 2639 25313 2651 25316
rect 2593 25307 2651 25313
rect 3694 25304 3700 25316
rect 3752 25304 3758 25356
rect 9953 25347 10011 25353
rect 9953 25344 9965 25347
rect 4724 25316 9965 25344
rect 1854 25276 1860 25288
rect 1815 25248 1860 25276
rect 1854 25236 1860 25248
rect 1912 25236 1918 25288
rect 2406 25236 2412 25288
rect 2464 25276 2470 25288
rect 4724 25285 4752 25316
rect 9953 25313 9965 25316
rect 9999 25313 10011 25347
rect 9953 25307 10011 25313
rect 2501 25279 2559 25285
rect 2501 25276 2513 25279
rect 2464 25248 2513 25276
rect 2464 25236 2470 25248
rect 2501 25245 2513 25248
rect 2547 25245 2559 25279
rect 2501 25239 2559 25245
rect 3145 25279 3203 25285
rect 3145 25245 3157 25279
rect 3191 25245 3203 25279
rect 3145 25239 3203 25245
rect 4709 25279 4767 25285
rect 4709 25245 4721 25279
rect 4755 25245 4767 25279
rect 5166 25276 5172 25288
rect 5079 25248 5172 25276
rect 4709 25239 4767 25245
rect 1949 25211 2007 25217
rect 1949 25177 1961 25211
rect 1995 25208 2007 25211
rect 3050 25208 3056 25220
rect 1995 25180 3056 25208
rect 1995 25177 2007 25180
rect 1949 25171 2007 25177
rect 3050 25168 3056 25180
rect 3108 25168 3114 25220
rect 2130 25100 2136 25152
rect 2188 25140 2194 25152
rect 3160 25140 3188 25239
rect 5166 25236 5172 25248
rect 5224 25236 5230 25288
rect 5810 25276 5816 25288
rect 5771 25248 5816 25276
rect 5810 25236 5816 25248
rect 5868 25236 5874 25288
rect 6454 25276 6460 25288
rect 6415 25248 6460 25276
rect 6454 25236 6460 25248
rect 6512 25236 6518 25288
rect 7285 25279 7343 25285
rect 7285 25245 7297 25279
rect 7331 25276 7343 25279
rect 7374 25276 7380 25288
rect 7331 25248 7380 25276
rect 7331 25245 7343 25248
rect 7285 25239 7343 25245
rect 7374 25236 7380 25248
rect 7432 25236 7438 25288
rect 7745 25279 7803 25285
rect 7745 25276 7757 25279
rect 7484 25248 7757 25276
rect 5184 25208 5212 25236
rect 6270 25208 6276 25220
rect 5184 25180 6276 25208
rect 6270 25168 6276 25180
rect 6328 25168 6334 25220
rect 6822 25168 6828 25220
rect 6880 25208 6886 25220
rect 7484 25208 7512 25248
rect 7745 25245 7757 25248
rect 7791 25245 7803 25279
rect 8570 25276 8576 25288
rect 8531 25248 8576 25276
rect 7745 25239 7803 25245
rect 8570 25236 8576 25248
rect 8628 25236 8634 25288
rect 8754 25236 8760 25288
rect 8812 25276 8818 25288
rect 10060 25285 10088 25384
rect 12986 25344 12992 25356
rect 12947 25316 12992 25344
rect 12986 25304 12992 25316
rect 13044 25304 13050 25356
rect 13648 25353 13676 25384
rect 15381 25381 15393 25384
rect 15427 25412 15439 25415
rect 16485 25415 16543 25421
rect 16485 25412 16497 25415
rect 15427 25384 16497 25412
rect 15427 25381 15439 25384
rect 15381 25375 15439 25381
rect 16485 25381 16497 25384
rect 16531 25381 16543 25415
rect 16485 25375 16543 25381
rect 13633 25347 13691 25353
rect 13633 25313 13645 25347
rect 13679 25313 13691 25347
rect 15194 25344 15200 25356
rect 15155 25316 15200 25344
rect 13633 25307 13691 25313
rect 15194 25304 15200 25316
rect 15252 25304 15258 25356
rect 16117 25347 16175 25353
rect 16117 25313 16129 25347
rect 16163 25344 16175 25347
rect 16206 25344 16212 25356
rect 16163 25316 16212 25344
rect 16163 25313 16175 25316
rect 16117 25307 16175 25313
rect 16206 25304 16212 25316
rect 16264 25304 16270 25356
rect 18509 25347 18567 25353
rect 18509 25313 18521 25347
rect 18555 25344 18567 25347
rect 18874 25344 18880 25356
rect 18555 25316 18880 25344
rect 18555 25313 18567 25316
rect 18509 25307 18567 25313
rect 18874 25304 18880 25316
rect 18932 25304 18938 25356
rect 9217 25279 9275 25285
rect 9217 25276 9229 25279
rect 8812 25248 9229 25276
rect 8812 25236 8818 25248
rect 9217 25245 9229 25248
rect 9263 25245 9275 25279
rect 9217 25239 9275 25245
rect 10045 25279 10103 25285
rect 10045 25245 10057 25279
rect 10091 25245 10103 25279
rect 10045 25239 10103 25245
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25245 10563 25279
rect 10505 25239 10563 25245
rect 11885 25279 11943 25285
rect 11885 25245 11897 25279
rect 11931 25276 11943 25279
rect 12710 25276 12716 25288
rect 11931 25248 12716 25276
rect 11931 25245 11943 25248
rect 11885 25239 11943 25245
rect 6880 25180 7512 25208
rect 6880 25168 6886 25180
rect 9490 25168 9496 25220
rect 9548 25208 9554 25220
rect 10520 25208 10548 25239
rect 12710 25236 12716 25248
rect 12768 25236 12774 25288
rect 15010 25276 15016 25288
rect 14971 25248 15016 25276
rect 15010 25236 15016 25248
rect 15068 25236 15074 25288
rect 16022 25236 16028 25288
rect 16080 25276 16086 25288
rect 16301 25279 16359 25285
rect 16301 25276 16313 25279
rect 16080 25248 16313 25276
rect 16080 25236 16086 25248
rect 16301 25245 16313 25248
rect 16347 25245 16359 25279
rect 16301 25239 16359 25245
rect 16666 25236 16672 25288
rect 16724 25276 16730 25288
rect 17405 25279 17463 25285
rect 17405 25276 17417 25279
rect 16724 25248 17417 25276
rect 16724 25236 16730 25248
rect 17405 25245 17417 25248
rect 17451 25245 17463 25279
rect 17405 25239 17463 25245
rect 18230 25236 18236 25288
rect 18288 25276 18294 25288
rect 18693 25279 18751 25285
rect 18693 25276 18705 25279
rect 18288 25248 18705 25276
rect 18288 25236 18294 25248
rect 18693 25245 18705 25248
rect 18739 25276 18751 25279
rect 18966 25276 18972 25288
rect 18739 25248 18972 25276
rect 18739 25245 18751 25248
rect 18693 25239 18751 25245
rect 18966 25236 18972 25248
rect 19024 25236 19030 25288
rect 19518 25236 19524 25288
rect 19576 25276 19582 25288
rect 19705 25279 19763 25285
rect 19705 25276 19717 25279
rect 19576 25248 19717 25276
rect 19576 25236 19582 25248
rect 19705 25245 19717 25248
rect 19751 25245 19763 25279
rect 20349 25279 20407 25285
rect 20349 25276 20361 25279
rect 19705 25239 19763 25245
rect 19904 25248 20361 25276
rect 13538 25208 13544 25220
rect 9548 25180 10548 25208
rect 13499 25180 13544 25208
rect 9548 25168 9554 25180
rect 13538 25168 13544 25180
rect 13596 25168 13602 25220
rect 2188 25112 3188 25140
rect 2188 25100 2194 25112
rect 3602 25100 3608 25152
rect 3660 25140 3666 25152
rect 4525 25143 4583 25149
rect 4525 25140 4537 25143
rect 3660 25112 4537 25140
rect 3660 25100 3666 25112
rect 4525 25109 4537 25112
rect 4571 25109 4583 25143
rect 5258 25140 5264 25152
rect 5219 25112 5264 25140
rect 4525 25103 4583 25109
rect 5258 25100 5264 25112
rect 5316 25100 5322 25152
rect 5997 25143 6055 25149
rect 5997 25109 6009 25143
rect 6043 25140 6055 25143
rect 6546 25140 6552 25152
rect 6043 25112 6552 25140
rect 6043 25109 6055 25112
rect 5997 25103 6055 25109
rect 6546 25100 6552 25112
rect 6604 25100 6610 25152
rect 6641 25143 6699 25149
rect 6641 25109 6653 25143
rect 6687 25140 6699 25143
rect 6730 25140 6736 25152
rect 6687 25112 6736 25140
rect 6687 25109 6699 25112
rect 6641 25103 6699 25109
rect 6730 25100 6736 25112
rect 6788 25100 6794 25152
rect 7193 25143 7251 25149
rect 7193 25109 7205 25143
rect 7239 25140 7251 25143
rect 7650 25140 7656 25152
rect 7239 25112 7656 25140
rect 7239 25109 7251 25112
rect 7193 25103 7251 25109
rect 7650 25100 7656 25112
rect 7708 25100 7714 25152
rect 7834 25140 7840 25152
rect 7795 25112 7840 25140
rect 7834 25100 7840 25112
rect 7892 25100 7898 25152
rect 9306 25140 9312 25152
rect 9267 25112 9312 25140
rect 9306 25100 9312 25112
rect 9364 25100 9370 25152
rect 9766 25100 9772 25152
rect 9824 25140 9830 25152
rect 10318 25140 10324 25152
rect 9824 25112 10324 25140
rect 9824 25100 9830 25112
rect 10318 25100 10324 25112
rect 10376 25100 10382 25152
rect 10594 25140 10600 25152
rect 10555 25112 10600 25140
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 11146 25100 11152 25152
rect 11204 25140 11210 25152
rect 11701 25143 11759 25149
rect 11701 25140 11713 25143
rect 11204 25112 11713 25140
rect 11204 25100 11210 25112
rect 11701 25109 11713 25112
rect 11747 25109 11759 25143
rect 11701 25103 11759 25109
rect 12529 25143 12587 25149
rect 12529 25109 12541 25143
rect 12575 25140 12587 25143
rect 13078 25140 13084 25152
rect 12575 25112 13084 25140
rect 12575 25109 12587 25112
rect 12529 25103 12587 25109
rect 13078 25100 13084 25112
rect 13136 25100 13142 25152
rect 14277 25143 14335 25149
rect 14277 25109 14289 25143
rect 14323 25140 14335 25143
rect 14366 25140 14372 25152
rect 14323 25112 14372 25140
rect 14323 25109 14335 25112
rect 14277 25103 14335 25109
rect 14366 25100 14372 25112
rect 14424 25100 14430 25152
rect 17589 25143 17647 25149
rect 17589 25109 17601 25143
rect 17635 25140 17647 25143
rect 17954 25140 17960 25152
rect 17635 25112 17960 25140
rect 17635 25109 17647 25112
rect 17589 25103 17647 25109
rect 17954 25100 17960 25112
rect 18012 25100 18018 25152
rect 19904 25149 19932 25248
rect 20349 25245 20361 25248
rect 20395 25245 20407 25279
rect 35618 25276 35624 25288
rect 35579 25248 35624 25276
rect 20349 25239 20407 25245
rect 35618 25236 35624 25248
rect 35676 25236 35682 25288
rect 38286 25276 38292 25288
rect 38247 25248 38292 25276
rect 38286 25236 38292 25248
rect 38344 25236 38350 25288
rect 19889 25143 19947 25149
rect 19889 25109 19901 25143
rect 19935 25109 19947 25143
rect 19889 25103 19947 25109
rect 20533 25143 20591 25149
rect 20533 25109 20545 25143
rect 20579 25140 20591 25143
rect 20898 25140 20904 25152
rect 20579 25112 20904 25140
rect 20579 25109 20591 25112
rect 20533 25103 20591 25109
rect 20898 25100 20904 25112
rect 20956 25100 20962 25152
rect 34790 25100 34796 25152
rect 34848 25140 34854 25152
rect 38105 25143 38163 25149
rect 38105 25140 38117 25143
rect 34848 25112 38117 25140
rect 34848 25100 34854 25112
rect 38105 25109 38117 25112
rect 38151 25109 38163 25143
rect 38105 25103 38163 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 5810 24896 5816 24948
rect 5868 24936 5874 24948
rect 5997 24939 6055 24945
rect 5997 24936 6009 24939
rect 5868 24908 6009 24936
rect 5868 24896 5874 24908
rect 5997 24905 6009 24908
rect 6043 24905 6055 24939
rect 5997 24899 6055 24905
rect 6086 24896 6092 24948
rect 6144 24936 6150 24948
rect 8754 24936 8760 24948
rect 6144 24908 8760 24936
rect 6144 24896 6150 24908
rect 8754 24896 8760 24908
rect 8812 24896 8818 24948
rect 9306 24896 9312 24948
rect 9364 24936 9370 24948
rect 11790 24936 11796 24948
rect 9364 24908 11796 24936
rect 9364 24896 9370 24908
rect 11790 24896 11796 24908
rect 11848 24896 11854 24948
rect 11974 24896 11980 24948
rect 12032 24936 12038 24948
rect 15930 24936 15936 24948
rect 12032 24908 15936 24936
rect 12032 24896 12038 24908
rect 15930 24896 15936 24908
rect 15988 24896 15994 24948
rect 5442 24828 5448 24880
rect 5500 24828 5506 24880
rect 12805 24871 12863 24877
rect 5828 24840 7328 24868
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24769 1915 24803
rect 2406 24800 2412 24812
rect 2367 24772 2412 24800
rect 1857 24763 1915 24769
rect 1872 24732 1900 24763
rect 2406 24760 2412 24772
rect 2464 24760 2470 24812
rect 3050 24800 3056 24812
rect 3011 24772 3056 24800
rect 3050 24760 3056 24772
rect 3108 24760 3114 24812
rect 3234 24800 3240 24812
rect 3195 24772 3240 24800
rect 3234 24760 3240 24772
rect 3292 24760 3298 24812
rect 4433 24803 4491 24809
rect 4433 24769 4445 24803
rect 4479 24800 4491 24803
rect 4614 24800 4620 24812
rect 4479 24772 4620 24800
rect 4479 24769 4491 24772
rect 4433 24763 4491 24769
rect 4614 24760 4620 24772
rect 4672 24760 4678 24812
rect 4890 24800 4896 24812
rect 4851 24772 4896 24800
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 5166 24760 5172 24812
rect 5224 24800 5230 24812
rect 5460 24800 5488 24828
rect 5828 24812 5856 24840
rect 5810 24800 5816 24812
rect 5224 24772 5488 24800
rect 5771 24772 5816 24800
rect 5224 24760 5230 24772
rect 5810 24760 5816 24772
rect 5868 24760 5874 24812
rect 7300 24809 7328 24840
rect 8312 24840 9812 24868
rect 6641 24803 6699 24809
rect 6641 24769 6653 24803
rect 6687 24769 6699 24803
rect 6641 24763 6699 24769
rect 7285 24803 7343 24809
rect 7285 24769 7297 24803
rect 7331 24769 7343 24803
rect 7285 24763 7343 24769
rect 3602 24732 3608 24744
rect 1872 24704 3608 24732
rect 3602 24692 3608 24704
rect 3660 24692 3666 24744
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24732 3755 24735
rect 4249 24735 4307 24741
rect 4249 24732 4261 24735
rect 3743 24704 4261 24732
rect 3743 24701 3755 24704
rect 3697 24695 3755 24701
rect 4249 24701 4261 24704
rect 4295 24732 4307 24735
rect 5442 24732 5448 24744
rect 4295 24704 5448 24732
rect 4295 24701 4307 24704
rect 4249 24695 4307 24701
rect 5442 24692 5448 24704
rect 5500 24692 5506 24744
rect 1854 24624 1860 24676
rect 1912 24664 1918 24676
rect 6656 24664 6684 24763
rect 7834 24760 7840 24812
rect 7892 24800 7898 24812
rect 8113 24803 8171 24809
rect 8113 24800 8125 24803
rect 7892 24772 8125 24800
rect 7892 24760 7898 24772
rect 8113 24769 8125 24772
rect 8159 24769 8171 24803
rect 8113 24763 8171 24769
rect 7926 24732 7932 24744
rect 7887 24704 7932 24732
rect 7926 24692 7932 24704
rect 7984 24732 7990 24744
rect 8312 24732 8340 24840
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 9033 24803 9091 24809
rect 9033 24800 9045 24803
rect 8444 24772 9045 24800
rect 8444 24760 8450 24772
rect 9033 24769 9045 24772
rect 9079 24769 9091 24803
rect 9674 24800 9680 24812
rect 9635 24772 9680 24800
rect 9033 24763 9091 24769
rect 9674 24760 9680 24772
rect 9732 24760 9738 24812
rect 9784 24800 9812 24840
rect 12805 24837 12817 24871
rect 12851 24868 12863 24871
rect 12986 24868 12992 24880
rect 12851 24840 12992 24868
rect 12851 24837 12863 24840
rect 12805 24831 12863 24837
rect 12986 24828 12992 24840
rect 13044 24828 13050 24880
rect 13354 24868 13360 24880
rect 13315 24840 13360 24868
rect 13354 24828 13360 24840
rect 13412 24828 13418 24880
rect 18690 24868 18696 24880
rect 18651 24840 18696 24868
rect 18690 24828 18696 24840
rect 18748 24828 18754 24880
rect 9950 24800 9956 24812
rect 9784 24772 9956 24800
rect 9950 24760 9956 24772
rect 10008 24760 10014 24812
rect 10318 24800 10324 24812
rect 10279 24772 10324 24800
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 11885 24803 11943 24809
rect 10980 24772 11836 24800
rect 7984 24704 8340 24732
rect 7984 24692 7990 24704
rect 8662 24692 8668 24744
rect 8720 24732 8726 24744
rect 10980 24732 11008 24772
rect 11146 24732 11152 24744
rect 8720 24704 11008 24732
rect 11107 24704 11152 24732
rect 8720 24692 8726 24704
rect 11146 24692 11152 24704
rect 11204 24692 11210 24744
rect 11701 24735 11759 24741
rect 11701 24701 11713 24735
rect 11747 24701 11759 24735
rect 11808 24732 11836 24772
rect 11885 24769 11897 24803
rect 11931 24800 11943 24803
rect 11974 24800 11980 24812
rect 11931 24772 11980 24800
rect 11931 24769 11943 24772
rect 11885 24763 11943 24769
rect 11974 24760 11980 24772
rect 12032 24760 12038 24812
rect 13630 24760 13636 24812
rect 13688 24800 13694 24812
rect 14645 24803 14703 24809
rect 14645 24800 14657 24803
rect 13688 24772 14657 24800
rect 13688 24760 13694 24772
rect 14645 24769 14657 24772
rect 14691 24769 14703 24803
rect 14645 24763 14703 24769
rect 15470 24760 15476 24812
rect 15528 24800 15534 24812
rect 15565 24803 15623 24809
rect 15565 24800 15577 24803
rect 15528 24772 15577 24800
rect 15528 24760 15534 24772
rect 15565 24769 15577 24772
rect 15611 24769 15623 24803
rect 15746 24800 15752 24812
rect 15707 24772 15752 24800
rect 15565 24763 15623 24769
rect 15746 24760 15752 24772
rect 15804 24760 15810 24812
rect 16758 24760 16764 24812
rect 16816 24800 16822 24812
rect 17589 24803 17647 24809
rect 17589 24800 17601 24803
rect 16816 24772 17601 24800
rect 16816 24760 16822 24772
rect 17589 24769 17601 24772
rect 17635 24769 17647 24803
rect 17589 24763 17647 24769
rect 17678 24760 17684 24812
rect 17736 24800 17742 24812
rect 18414 24800 18420 24812
rect 17736 24772 18420 24800
rect 17736 24760 17742 24772
rect 18414 24760 18420 24772
rect 18472 24760 18478 24812
rect 20530 24800 20536 24812
rect 20491 24772 20536 24800
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 20714 24800 20720 24812
rect 20675 24772 20720 24800
rect 20714 24760 20720 24772
rect 20772 24760 20778 24812
rect 37550 24800 37556 24812
rect 20824 24772 37556 24800
rect 13449 24735 13507 24741
rect 11808 24704 13308 24732
rect 11701 24695 11759 24701
rect 1912 24636 6684 24664
rect 6733 24667 6791 24673
rect 1912 24624 1918 24636
rect 6733 24633 6745 24667
rect 6779 24664 6791 24667
rect 11716 24664 11744 24695
rect 6779 24636 11744 24664
rect 13280 24664 13308 24704
rect 13449 24701 13461 24735
rect 13495 24732 13507 24735
rect 14829 24735 14887 24741
rect 13495 24704 14780 24732
rect 13495 24701 13507 24704
rect 13449 24695 13507 24701
rect 14185 24667 14243 24673
rect 14185 24664 14197 24667
rect 13280 24636 14197 24664
rect 6779 24633 6791 24636
rect 6733 24627 6791 24633
rect 14185 24633 14197 24636
rect 14231 24633 14243 24667
rect 14185 24627 14243 24633
rect 1670 24596 1676 24608
rect 1631 24568 1676 24596
rect 1670 24556 1676 24568
rect 1728 24556 1734 24608
rect 2501 24599 2559 24605
rect 2501 24565 2513 24599
rect 2547 24596 2559 24599
rect 5994 24596 6000 24608
rect 2547 24568 6000 24596
rect 2547 24565 2559 24568
rect 2501 24559 2559 24565
rect 5994 24556 6000 24568
rect 6052 24556 6058 24608
rect 7377 24599 7435 24605
rect 7377 24565 7389 24599
rect 7423 24596 7435 24599
rect 7834 24596 7840 24608
rect 7423 24568 7840 24596
rect 7423 24565 7435 24568
rect 7377 24559 7435 24565
rect 7834 24556 7840 24568
rect 7892 24556 7898 24608
rect 8573 24599 8631 24605
rect 8573 24565 8585 24599
rect 8619 24596 8631 24599
rect 8938 24596 8944 24608
rect 8619 24568 8944 24596
rect 8619 24565 8631 24568
rect 8573 24559 8631 24565
rect 8938 24556 8944 24568
rect 8996 24556 9002 24608
rect 9122 24596 9128 24608
rect 9083 24568 9128 24596
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 9858 24596 9864 24608
rect 9819 24568 9864 24596
rect 9858 24556 9864 24568
rect 9916 24556 9922 24608
rect 10410 24596 10416 24608
rect 10371 24568 10416 24596
rect 10410 24556 10416 24568
rect 10468 24556 10474 24608
rect 11238 24556 11244 24608
rect 11296 24596 11302 24608
rect 12069 24599 12127 24605
rect 12069 24596 12081 24599
rect 11296 24568 12081 24596
rect 11296 24556 11302 24568
rect 12069 24565 12081 24568
rect 12115 24565 12127 24599
rect 14752 24596 14780 24704
rect 14829 24701 14841 24735
rect 14875 24701 14887 24735
rect 14829 24695 14887 24701
rect 16209 24735 16267 24741
rect 16209 24701 16221 24735
rect 16255 24732 16267 24735
rect 16574 24732 16580 24744
rect 16255 24704 16580 24732
rect 16255 24701 16267 24704
rect 16209 24695 16267 24701
rect 14844 24664 14872 24695
rect 16574 24692 16580 24704
rect 16632 24732 16638 24744
rect 16850 24732 16856 24744
rect 16632 24704 16856 24732
rect 16632 24692 16638 24704
rect 16850 24692 16856 24704
rect 16908 24692 16914 24744
rect 17405 24735 17463 24741
rect 17405 24701 17417 24735
rect 17451 24732 17463 24735
rect 17862 24732 17868 24744
rect 17451 24704 17868 24732
rect 17451 24701 17463 24704
rect 17405 24695 17463 24701
rect 17862 24692 17868 24704
rect 17920 24692 17926 24744
rect 18601 24735 18659 24741
rect 18601 24701 18613 24735
rect 18647 24732 18659 24735
rect 18782 24732 18788 24744
rect 18647 24704 18788 24732
rect 18647 24701 18659 24704
rect 18601 24695 18659 24701
rect 18782 24692 18788 24704
rect 18840 24692 18846 24744
rect 19613 24735 19671 24741
rect 19613 24701 19625 24735
rect 19659 24732 19671 24735
rect 19978 24732 19984 24744
rect 19659 24704 19984 24732
rect 19659 24701 19671 24704
rect 19613 24695 19671 24701
rect 19978 24692 19984 24704
rect 20036 24732 20042 24744
rect 20824 24732 20852 24772
rect 37550 24760 37556 24772
rect 37608 24760 37614 24812
rect 20036 24704 20852 24732
rect 20036 24692 20042 24704
rect 21082 24692 21088 24744
rect 21140 24732 21146 24744
rect 21177 24735 21235 24741
rect 21177 24732 21189 24735
rect 21140 24704 21189 24732
rect 21140 24692 21146 24704
rect 21177 24701 21189 24704
rect 21223 24701 21235 24735
rect 21177 24695 21235 24701
rect 15010 24664 15016 24676
rect 14844 24636 15016 24664
rect 15010 24624 15016 24636
rect 15068 24664 15074 24676
rect 20806 24664 20812 24676
rect 15068 24636 20812 24664
rect 15068 24624 15074 24636
rect 20806 24624 20812 24636
rect 20864 24624 20870 24676
rect 17678 24596 17684 24608
rect 14752 24568 17684 24596
rect 12069 24559 12127 24565
rect 17678 24556 17684 24568
rect 17736 24556 17742 24608
rect 17770 24556 17776 24608
rect 17828 24596 17834 24608
rect 17957 24599 18015 24605
rect 17957 24596 17969 24599
rect 17828 24568 17969 24596
rect 17828 24556 17834 24568
rect 17957 24565 17969 24568
rect 18003 24565 18015 24599
rect 20070 24596 20076 24608
rect 20031 24568 20076 24596
rect 17957 24559 18015 24565
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 2406 24352 2412 24404
rect 2464 24392 2470 24404
rect 4246 24392 4252 24404
rect 2464 24364 4252 24392
rect 2464 24352 2470 24364
rect 4246 24352 4252 24364
rect 4304 24352 4310 24404
rect 4617 24395 4675 24401
rect 4617 24361 4629 24395
rect 4663 24392 4675 24395
rect 4890 24392 4896 24404
rect 4663 24364 4896 24392
rect 4663 24361 4675 24364
rect 4617 24355 4675 24361
rect 4890 24352 4896 24364
rect 4948 24352 4954 24404
rect 7558 24392 7564 24404
rect 5000 24364 7564 24392
rect 2958 24284 2964 24336
rect 3016 24324 3022 24336
rect 5000 24324 5028 24364
rect 7558 24352 7564 24364
rect 7616 24352 7622 24404
rect 7742 24352 7748 24404
rect 7800 24392 7806 24404
rect 9766 24392 9772 24404
rect 7800 24364 9772 24392
rect 7800 24352 7806 24364
rect 9766 24352 9772 24364
rect 9824 24352 9830 24404
rect 9858 24352 9864 24404
rect 9916 24392 9922 24404
rect 11882 24392 11888 24404
rect 9916 24364 11888 24392
rect 9916 24352 9922 24364
rect 11882 24352 11888 24364
rect 11940 24352 11946 24404
rect 12710 24352 12716 24404
rect 12768 24392 12774 24404
rect 16482 24392 16488 24404
rect 12768 24364 16488 24392
rect 12768 24352 12774 24364
rect 16482 24352 16488 24364
rect 16540 24352 16546 24404
rect 16945 24395 17003 24401
rect 16945 24361 16957 24395
rect 16991 24392 17003 24395
rect 18690 24392 18696 24404
rect 16991 24364 18696 24392
rect 16991 24361 17003 24364
rect 16945 24355 17003 24361
rect 18690 24352 18696 24364
rect 18748 24352 18754 24404
rect 35342 24392 35348 24404
rect 35303 24364 35348 24392
rect 35342 24352 35348 24364
rect 35400 24352 35406 24404
rect 3016 24296 5028 24324
rect 5997 24327 6055 24333
rect 3016 24284 3022 24296
rect 5997 24293 6009 24327
rect 6043 24324 6055 24327
rect 8938 24324 8944 24336
rect 6043 24296 8944 24324
rect 6043 24293 6055 24296
rect 5997 24287 6055 24293
rect 8938 24284 8944 24296
rect 8996 24284 9002 24336
rect 12342 24324 12348 24336
rect 10980 24296 12348 24324
rect 2777 24259 2835 24265
rect 2777 24225 2789 24259
rect 2823 24256 2835 24259
rect 3973 24259 4031 24265
rect 3973 24256 3985 24259
rect 2823 24228 3985 24256
rect 2823 24225 2835 24228
rect 2777 24219 2835 24225
rect 3973 24225 3985 24228
rect 4019 24225 4031 24259
rect 3973 24219 4031 24225
rect 4157 24259 4215 24265
rect 4157 24225 4169 24259
rect 4203 24256 4215 24259
rect 4706 24256 4712 24268
rect 4203 24228 4712 24256
rect 4203 24225 4215 24228
rect 4157 24219 4215 24225
rect 4706 24216 4712 24228
rect 4764 24216 4770 24268
rect 5166 24256 5172 24268
rect 5000 24228 5172 24256
rect 5000 24200 5028 24228
rect 5166 24216 5172 24228
rect 5224 24216 5230 24268
rect 5350 24256 5356 24268
rect 5311 24228 5356 24256
rect 5350 24216 5356 24228
rect 5408 24216 5414 24268
rect 5534 24256 5540 24268
rect 5495 24228 5540 24256
rect 5534 24216 5540 24228
rect 5592 24216 5598 24268
rect 6178 24216 6184 24268
rect 6236 24256 6242 24268
rect 6549 24259 6607 24265
rect 6549 24256 6561 24259
rect 6236 24228 6561 24256
rect 6236 24216 6242 24228
rect 6549 24225 6561 24228
rect 6595 24225 6607 24259
rect 6549 24219 6607 24225
rect 7193 24259 7251 24265
rect 7193 24225 7205 24259
rect 7239 24256 7251 24259
rect 7668 24256 7880 24268
rect 8021 24259 8079 24265
rect 8021 24256 8033 24259
rect 7239 24240 8033 24256
rect 7239 24228 7696 24240
rect 7852 24228 8033 24240
rect 7239 24225 7251 24228
rect 7193 24219 7251 24225
rect 8021 24225 8033 24228
rect 8067 24256 8079 24259
rect 10042 24256 10048 24268
rect 8067 24228 10048 24256
rect 8067 24225 8079 24228
rect 8021 24219 8079 24225
rect 10042 24216 10048 24228
rect 10100 24216 10106 24268
rect 1486 24148 1492 24200
rect 1544 24188 1550 24200
rect 1949 24191 2007 24197
rect 1949 24188 1961 24191
rect 1544 24160 1961 24188
rect 1544 24148 1550 24160
rect 1949 24157 1961 24160
rect 1995 24188 2007 24191
rect 2130 24188 2136 24200
rect 1995 24160 2136 24188
rect 1995 24157 2007 24160
rect 1949 24151 2007 24157
rect 2130 24148 2136 24160
rect 2188 24148 2194 24200
rect 2222 24148 2228 24200
rect 2280 24188 2286 24200
rect 3421 24191 3479 24197
rect 3421 24188 3433 24191
rect 2280 24160 3433 24188
rect 2280 24148 2286 24160
rect 3421 24157 3433 24160
rect 3467 24157 3479 24191
rect 3421 24151 3479 24157
rect 4982 24148 4988 24200
rect 5040 24148 5046 24200
rect 5810 24148 5816 24200
rect 5868 24188 5874 24200
rect 6270 24188 6276 24200
rect 5868 24160 6276 24188
rect 5868 24148 5874 24160
rect 6270 24148 6276 24160
rect 6328 24148 6334 24200
rect 9306 24188 9312 24200
rect 8496 24160 9312 24188
rect 2041 24123 2099 24129
rect 2041 24089 2053 24123
rect 2087 24120 2099 24123
rect 5166 24120 5172 24132
rect 2087 24092 5172 24120
rect 2087 24089 2099 24092
rect 2041 24083 2099 24089
rect 5166 24080 5172 24092
rect 5224 24080 5230 24132
rect 6638 24080 6644 24132
rect 6696 24120 6702 24132
rect 7742 24120 7748 24132
rect 6696 24092 6741 24120
rect 7703 24092 7748 24120
rect 6696 24080 6702 24092
rect 7742 24080 7748 24092
rect 7800 24080 7806 24132
rect 7834 24080 7840 24132
rect 7892 24120 7898 24132
rect 7892 24092 7937 24120
rect 7892 24080 7898 24092
rect 8202 24080 8208 24132
rect 8260 24120 8266 24132
rect 8496 24120 8524 24160
rect 9306 24148 9312 24160
rect 9364 24148 9370 24200
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24157 10011 24191
rect 9953 24151 10011 24157
rect 10597 24191 10655 24197
rect 10597 24157 10609 24191
rect 10643 24188 10655 24191
rect 10980 24188 11008 24296
rect 12342 24284 12348 24296
rect 12400 24284 12406 24336
rect 14642 24324 14648 24336
rect 14603 24296 14648 24324
rect 14642 24284 14648 24296
rect 14700 24284 14706 24336
rect 25406 24324 25412 24336
rect 17512 24296 25412 24324
rect 11054 24216 11060 24268
rect 11112 24256 11118 24268
rect 11425 24259 11483 24265
rect 11425 24256 11437 24259
rect 11112 24228 11437 24256
rect 11112 24216 11118 24228
rect 11425 24225 11437 24228
rect 11471 24225 11483 24259
rect 11425 24219 11483 24225
rect 11514 24216 11520 24268
rect 11572 24256 11578 24268
rect 17512 24265 17540 24296
rect 25406 24284 25412 24296
rect 25464 24284 25470 24336
rect 17497 24259 17555 24265
rect 17497 24256 17509 24259
rect 11572 24228 17509 24256
rect 11572 24216 11578 24228
rect 17497 24225 17509 24228
rect 17543 24225 17555 24259
rect 17497 24219 17555 24225
rect 17586 24216 17592 24268
rect 17644 24256 17650 24268
rect 17681 24259 17739 24265
rect 17681 24256 17693 24259
rect 17644 24228 17693 24256
rect 17644 24216 17650 24228
rect 17681 24225 17693 24228
rect 17727 24225 17739 24259
rect 17681 24219 17739 24225
rect 17862 24216 17868 24268
rect 17920 24256 17926 24268
rect 20898 24256 20904 24268
rect 17920 24228 18828 24256
rect 20859 24228 20904 24256
rect 17920 24216 17926 24228
rect 10643 24160 11008 24188
rect 11241 24191 11299 24197
rect 10643 24157 10655 24160
rect 10597 24151 10655 24157
rect 11241 24157 11253 24191
rect 11287 24188 11299 24191
rect 11330 24188 11336 24200
rect 11287 24160 11336 24188
rect 11287 24157 11299 24160
rect 11241 24151 11299 24157
rect 8260 24092 8524 24120
rect 8260 24080 8266 24092
rect 8570 24080 8576 24132
rect 8628 24120 8634 24132
rect 9968 24120 9996 24151
rect 11330 24148 11336 24160
rect 11388 24148 11394 24200
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 14458 24188 14464 24200
rect 13587 24160 14464 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 14458 24148 14464 24160
rect 14516 24148 14522 24200
rect 16298 24148 16304 24200
rect 16356 24188 16362 24200
rect 16393 24191 16451 24197
rect 16393 24188 16405 24191
rect 16356 24160 16405 24188
rect 16356 24148 16362 24160
rect 16393 24157 16405 24160
rect 16439 24157 16451 24191
rect 16393 24151 16451 24157
rect 16666 24148 16672 24200
rect 16724 24188 16730 24200
rect 16853 24191 16911 24197
rect 16853 24188 16865 24191
rect 16724 24160 16865 24188
rect 16724 24148 16730 24160
rect 16853 24157 16865 24160
rect 16899 24157 16911 24191
rect 16853 24151 16911 24157
rect 17954 24148 17960 24200
rect 18012 24188 18018 24200
rect 18693 24191 18751 24197
rect 18693 24188 18705 24191
rect 18012 24160 18705 24188
rect 18012 24148 18018 24160
rect 18693 24157 18705 24160
rect 18739 24157 18751 24191
rect 18800 24188 18828 24228
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 21082 24256 21088 24268
rect 21043 24228 21088 24256
rect 21082 24216 21088 24228
rect 21140 24216 21146 24268
rect 27246 24188 27252 24200
rect 18800 24160 27252 24188
rect 18693 24151 18751 24157
rect 27246 24148 27252 24160
rect 27304 24148 27310 24200
rect 33134 24148 33140 24200
rect 33192 24188 33198 24200
rect 35161 24191 35219 24197
rect 35161 24188 35173 24191
rect 33192 24160 35173 24188
rect 33192 24148 33198 24160
rect 35161 24157 35173 24160
rect 35207 24157 35219 24191
rect 35161 24151 35219 24157
rect 14182 24120 14188 24132
rect 8628 24092 9996 24120
rect 10796 24092 14188 24120
rect 8628 24080 8634 24092
rect 3326 24052 3332 24064
rect 3287 24024 3332 24052
rect 3326 24012 3332 24024
rect 3384 24012 3390 24064
rect 7374 24012 7380 24064
rect 7432 24052 7438 24064
rect 8846 24052 8852 24064
rect 7432 24024 8852 24052
rect 7432 24012 7438 24024
rect 8846 24012 8852 24024
rect 8904 24012 8910 24064
rect 9398 24052 9404 24064
rect 9359 24024 9404 24052
rect 9398 24012 9404 24024
rect 9456 24012 9462 24064
rect 10134 24052 10140 24064
rect 10095 24024 10140 24052
rect 10134 24012 10140 24024
rect 10192 24012 10198 24064
rect 10796 24061 10824 24092
rect 14182 24080 14188 24092
rect 14240 24080 14246 24132
rect 14826 24080 14832 24132
rect 14884 24120 14890 24132
rect 15105 24123 15163 24129
rect 15105 24120 15117 24123
rect 14884 24092 15117 24120
rect 14884 24080 14890 24092
rect 15105 24089 15117 24092
rect 15151 24089 15163 24123
rect 15105 24083 15163 24089
rect 15197 24123 15255 24129
rect 15197 24089 15209 24123
rect 15243 24120 15255 24123
rect 16574 24120 16580 24132
rect 15243 24092 16580 24120
rect 15243 24089 15255 24092
rect 15197 24083 15255 24089
rect 16574 24080 16580 24092
rect 16632 24080 16638 24132
rect 17402 24080 17408 24132
rect 17460 24120 17466 24132
rect 20070 24120 20076 24132
rect 17460 24092 20076 24120
rect 17460 24080 17466 24092
rect 20070 24080 20076 24092
rect 20128 24120 20134 24132
rect 20441 24123 20499 24129
rect 20441 24120 20453 24123
rect 20128 24092 20453 24120
rect 20128 24080 20134 24092
rect 20441 24089 20453 24092
rect 20487 24089 20499 24123
rect 20441 24083 20499 24089
rect 10781 24055 10839 24061
rect 10781 24021 10793 24055
rect 10827 24021 10839 24055
rect 10781 24015 10839 24021
rect 11885 24055 11943 24061
rect 11885 24021 11897 24055
rect 11931 24052 11943 24055
rect 11974 24052 11980 24064
rect 11931 24024 11980 24052
rect 11931 24021 11943 24024
rect 11885 24015 11943 24021
rect 11974 24012 11980 24024
rect 12032 24012 12038 24064
rect 13081 24055 13139 24061
rect 13081 24021 13093 24055
rect 13127 24052 13139 24055
rect 13446 24052 13452 24064
rect 13127 24024 13452 24052
rect 13127 24021 13139 24024
rect 13081 24015 13139 24021
rect 13446 24012 13452 24024
rect 13504 24012 13510 24064
rect 13630 24052 13636 24064
rect 13591 24024 13636 24052
rect 13630 24012 13636 24024
rect 13688 24012 13694 24064
rect 13906 24012 13912 24064
rect 13964 24052 13970 24064
rect 16209 24055 16267 24061
rect 16209 24052 16221 24055
rect 13964 24024 16221 24052
rect 13964 24012 13970 24024
rect 16209 24021 16221 24024
rect 16255 24021 16267 24055
rect 16209 24015 16267 24021
rect 17770 24012 17776 24064
rect 17828 24052 17834 24064
rect 18141 24055 18199 24061
rect 18141 24052 18153 24055
rect 17828 24024 18153 24052
rect 17828 24012 17834 24024
rect 18141 24021 18153 24024
rect 18187 24021 18199 24055
rect 18141 24015 18199 24021
rect 18877 24055 18935 24061
rect 18877 24021 18889 24055
rect 18923 24052 18935 24055
rect 18966 24052 18972 24064
rect 18923 24024 18972 24052
rect 18923 24021 18935 24024
rect 18877 24015 18935 24021
rect 18966 24012 18972 24024
rect 19024 24012 19030 24064
rect 19426 24052 19432 24064
rect 19387 24024 19432 24052
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1765 23851 1823 23857
rect 1765 23817 1777 23851
rect 1811 23848 1823 23851
rect 1854 23848 1860 23860
rect 1811 23820 1860 23848
rect 1811 23817 1823 23820
rect 1765 23811 1823 23817
rect 1854 23808 1860 23820
rect 1912 23808 1918 23860
rect 3878 23808 3884 23860
rect 3936 23848 3942 23860
rect 3936 23820 4476 23848
rect 3936 23808 3942 23820
rect 4338 23780 4344 23792
rect 4299 23752 4344 23780
rect 4338 23740 4344 23752
rect 4396 23740 4402 23792
rect 4448 23780 4476 23820
rect 5258 23808 5264 23860
rect 5316 23848 5322 23860
rect 5316 23820 8800 23848
rect 5316 23808 5322 23820
rect 4448 23752 5856 23780
rect 1581 23715 1639 23721
rect 1581 23681 1593 23715
rect 1627 23681 1639 23715
rect 1581 23675 1639 23681
rect 2501 23715 2559 23721
rect 2501 23681 2513 23715
rect 2547 23712 2559 23715
rect 2590 23712 2596 23724
rect 2547 23684 2596 23712
rect 2547 23681 2559 23684
rect 2501 23675 2559 23681
rect 1596 23644 1624 23675
rect 2590 23672 2596 23684
rect 2648 23712 2654 23724
rect 2648 23684 2912 23712
rect 2648 23672 2654 23684
rect 2774 23644 2780 23656
rect 1596 23616 2780 23644
rect 2774 23604 2780 23616
rect 2832 23604 2838 23656
rect 2884 23644 2912 23684
rect 2958 23672 2964 23724
rect 3016 23712 3022 23724
rect 3605 23715 3663 23721
rect 3016 23684 3061 23712
rect 3016 23672 3022 23684
rect 3605 23681 3617 23715
rect 3651 23712 3663 23715
rect 3878 23712 3884 23724
rect 3651 23684 3884 23712
rect 3651 23681 3663 23684
rect 3605 23675 3663 23681
rect 3878 23672 3884 23684
rect 3936 23672 3942 23724
rect 4246 23712 4252 23724
rect 4159 23684 4252 23712
rect 4246 23672 4252 23684
rect 4304 23712 4310 23724
rect 4706 23712 4712 23724
rect 4304 23684 4712 23712
rect 4304 23672 4310 23684
rect 4706 23672 4712 23684
rect 4764 23672 4770 23724
rect 4982 23672 4988 23724
rect 5040 23712 5046 23724
rect 5828 23721 5856 23752
rect 7006 23740 7012 23792
rect 7064 23780 7070 23792
rect 7101 23783 7159 23789
rect 7101 23780 7113 23783
rect 7064 23752 7113 23780
rect 7064 23740 7070 23752
rect 7101 23749 7113 23752
rect 7147 23749 7159 23783
rect 7650 23780 7656 23792
rect 7611 23752 7656 23780
rect 7101 23743 7159 23749
rect 7650 23740 7656 23752
rect 7708 23740 7714 23792
rect 7745 23783 7803 23789
rect 7745 23749 7757 23783
rect 7791 23780 7803 23783
rect 8662 23780 8668 23792
rect 7791 23752 8668 23780
rect 7791 23749 7803 23752
rect 7745 23743 7803 23749
rect 8662 23740 8668 23752
rect 8720 23740 8726 23792
rect 5077 23715 5135 23721
rect 5077 23712 5089 23715
rect 5040 23684 5089 23712
rect 5040 23672 5046 23684
rect 5077 23681 5089 23684
rect 5123 23681 5135 23715
rect 5077 23675 5135 23681
rect 5813 23715 5871 23721
rect 5813 23681 5825 23715
rect 5859 23681 5871 23715
rect 5813 23675 5871 23681
rect 4614 23644 4620 23656
rect 2884 23616 4620 23644
rect 4614 23604 4620 23616
rect 4672 23604 4678 23656
rect 5092 23644 5120 23675
rect 8570 23672 8576 23724
rect 8628 23672 8634 23724
rect 8772 23721 8800 23820
rect 9306 23808 9312 23860
rect 9364 23848 9370 23860
rect 11606 23848 11612 23860
rect 9364 23820 11612 23848
rect 9364 23808 9370 23820
rect 11606 23808 11612 23820
rect 11664 23808 11670 23860
rect 13446 23808 13452 23860
rect 13504 23848 13510 23860
rect 20530 23848 20536 23860
rect 13504 23820 17540 23848
rect 13504 23808 13510 23820
rect 9398 23740 9404 23792
rect 9456 23780 9462 23792
rect 12069 23783 12127 23789
rect 12069 23780 12081 23783
rect 9456 23752 12081 23780
rect 9456 23740 9462 23752
rect 12069 23749 12081 23752
rect 12115 23749 12127 23783
rect 12069 23743 12127 23749
rect 13630 23740 13636 23792
rect 13688 23780 13694 23792
rect 13688 23752 16160 23780
rect 13688 23740 13694 23752
rect 8757 23715 8815 23721
rect 8757 23681 8769 23715
rect 8803 23681 8815 23715
rect 8757 23675 8815 23681
rect 9122 23672 9128 23724
rect 9180 23712 9186 23724
rect 9861 23715 9919 23721
rect 9861 23712 9873 23715
rect 9180 23684 9873 23712
rect 9180 23672 9186 23684
rect 9861 23681 9873 23684
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23712 11023 23715
rect 11698 23712 11704 23724
rect 11011 23684 11704 23712
rect 11011 23681 11023 23684
rect 10965 23675 11023 23681
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23681 13323 23715
rect 13906 23712 13912 23724
rect 13867 23684 13912 23712
rect 13265 23675 13323 23681
rect 5258 23644 5264 23656
rect 5092 23616 5264 23644
rect 5258 23604 5264 23616
rect 5316 23604 5322 23656
rect 6362 23604 6368 23656
rect 6420 23644 6426 23656
rect 8202 23644 8208 23656
rect 6420 23616 8208 23644
rect 6420 23604 6426 23616
rect 8202 23604 8208 23616
rect 8260 23604 8266 23656
rect 3050 23576 3056 23588
rect 3011 23548 3056 23576
rect 3050 23536 3056 23548
rect 3108 23536 3114 23588
rect 3697 23579 3755 23585
rect 3697 23545 3709 23579
rect 3743 23576 3755 23579
rect 5350 23576 5356 23588
rect 3743 23548 5356 23576
rect 3743 23545 3755 23548
rect 3697 23539 3755 23545
rect 5350 23536 5356 23548
rect 5408 23536 5414 23588
rect 5442 23536 5448 23588
rect 5500 23576 5506 23588
rect 8389 23579 8447 23585
rect 8389 23576 8401 23579
rect 5500 23548 8401 23576
rect 5500 23536 5506 23548
rect 8389 23545 8401 23548
rect 8435 23545 8447 23579
rect 8389 23539 8447 23545
rect 8588 23520 8616 23672
rect 8941 23647 8999 23653
rect 8941 23613 8953 23647
rect 8987 23644 8999 23647
rect 9677 23647 9735 23653
rect 9677 23644 9689 23647
rect 8987 23616 9689 23644
rect 8987 23613 8999 23616
rect 8941 23607 8999 23613
rect 9677 23613 9689 23616
rect 9723 23644 9735 23647
rect 11514 23644 11520 23656
rect 9723 23616 11520 23644
rect 9723 23613 9735 23616
rect 9677 23607 9735 23613
rect 11514 23604 11520 23616
rect 11572 23604 11578 23656
rect 11974 23644 11980 23656
rect 11935 23616 11980 23644
rect 11974 23604 11980 23616
rect 12032 23604 12038 23656
rect 13280 23644 13308 23675
rect 13906 23672 13912 23684
rect 13964 23672 13970 23724
rect 14550 23712 14556 23724
rect 14511 23684 14556 23712
rect 14550 23672 14556 23684
rect 14608 23672 14614 23724
rect 14734 23672 14740 23724
rect 14792 23712 14798 23724
rect 16132 23721 16160 23752
rect 15013 23715 15071 23721
rect 15013 23712 15025 23715
rect 14792 23684 15025 23712
rect 14792 23672 14798 23684
rect 15013 23681 15025 23684
rect 15059 23681 15071 23715
rect 15013 23675 15071 23681
rect 16117 23715 16175 23721
rect 16117 23681 16129 23715
rect 16163 23681 16175 23715
rect 17402 23712 17408 23724
rect 16117 23675 16175 23681
rect 16224 23684 17408 23712
rect 13814 23644 13820 23656
rect 13280 23616 13820 23644
rect 13814 23604 13820 23616
rect 13872 23604 13878 23656
rect 13998 23604 14004 23656
rect 14056 23644 14062 23656
rect 14918 23644 14924 23656
rect 14056 23616 14924 23644
rect 14056 23604 14062 23616
rect 14918 23604 14924 23616
rect 14976 23604 14982 23656
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23644 15255 23647
rect 16224 23644 16252 23684
rect 17402 23672 17408 23684
rect 17460 23672 17466 23724
rect 17512 23721 17540 23820
rect 18156 23820 20536 23848
rect 18156 23721 18184 23820
rect 20530 23808 20536 23820
rect 20588 23808 20594 23860
rect 18966 23780 18972 23792
rect 18927 23752 18972 23780
rect 18966 23740 18972 23752
rect 19024 23740 19030 23792
rect 19889 23783 19947 23789
rect 19889 23749 19901 23783
rect 19935 23780 19947 23783
rect 19978 23780 19984 23792
rect 19935 23752 19984 23780
rect 19935 23749 19947 23752
rect 19889 23743 19947 23749
rect 19978 23740 19984 23752
rect 20036 23740 20042 23792
rect 17497 23715 17555 23721
rect 17497 23681 17509 23715
rect 17543 23681 17555 23715
rect 17497 23675 17555 23681
rect 18141 23715 18199 23721
rect 18141 23681 18153 23715
rect 18187 23681 18199 23715
rect 18141 23675 18199 23681
rect 20438 23672 20444 23724
rect 20496 23712 20502 23724
rect 20533 23715 20591 23721
rect 20533 23712 20545 23715
rect 20496 23684 20545 23712
rect 20496 23672 20502 23684
rect 20533 23681 20545 23684
rect 20579 23681 20591 23715
rect 20533 23675 20591 23681
rect 33965 23715 34023 23721
rect 33965 23681 33977 23715
rect 34011 23712 34023 23715
rect 34790 23712 34796 23724
rect 34011 23684 34796 23712
rect 34011 23681 34023 23684
rect 33965 23675 34023 23681
rect 34790 23672 34796 23684
rect 34848 23672 34854 23724
rect 38286 23712 38292 23724
rect 38247 23684 38292 23712
rect 38286 23672 38292 23684
rect 38344 23672 38350 23724
rect 15243 23616 16252 23644
rect 16301 23647 16359 23653
rect 15243 23613 15255 23616
rect 15197 23607 15255 23613
rect 16301 23613 16313 23647
rect 16347 23644 16359 23647
rect 17313 23647 17371 23653
rect 16347 23616 17264 23644
rect 16347 23613 16359 23616
rect 16301 23607 16359 23613
rect 9950 23536 9956 23588
rect 10008 23576 10014 23588
rect 10962 23576 10968 23588
rect 10008 23548 10968 23576
rect 10008 23536 10014 23548
rect 10962 23536 10968 23548
rect 11020 23536 11026 23588
rect 12529 23579 12587 23585
rect 12529 23545 12541 23579
rect 12575 23576 12587 23579
rect 14642 23576 14648 23588
rect 12575 23548 14648 23576
rect 12575 23545 12587 23548
rect 12529 23539 12587 23545
rect 14642 23536 14648 23548
rect 14700 23536 14706 23588
rect 2409 23511 2467 23517
rect 2409 23477 2421 23511
rect 2455 23508 2467 23511
rect 2590 23508 2596 23520
rect 2455 23480 2596 23508
rect 2455 23477 2467 23480
rect 2409 23471 2467 23477
rect 2590 23468 2596 23480
rect 2648 23468 2654 23520
rect 4982 23508 4988 23520
rect 4943 23480 4988 23508
rect 4982 23468 4988 23480
rect 5040 23468 5046 23520
rect 5905 23511 5963 23517
rect 5905 23477 5917 23511
rect 5951 23508 5963 23511
rect 8478 23508 8484 23520
rect 5951 23480 8484 23508
rect 5951 23477 5963 23480
rect 5905 23471 5963 23477
rect 8478 23468 8484 23480
rect 8536 23468 8542 23520
rect 8570 23468 8576 23520
rect 8628 23468 8634 23520
rect 8938 23468 8944 23520
rect 8996 23508 9002 23520
rect 9398 23508 9404 23520
rect 8996 23480 9404 23508
rect 8996 23468 9002 23480
rect 9398 23468 9404 23480
rect 9456 23468 9462 23520
rect 10321 23511 10379 23517
rect 10321 23477 10333 23511
rect 10367 23508 10379 23511
rect 11054 23508 11060 23520
rect 10367 23480 11060 23508
rect 10367 23477 10379 23480
rect 10321 23471 10379 23477
rect 11054 23468 11060 23480
rect 11112 23468 11118 23520
rect 11149 23511 11207 23517
rect 11149 23477 11161 23511
rect 11195 23508 11207 23511
rect 13170 23508 13176 23520
rect 11195 23480 13176 23508
rect 11195 23477 11207 23480
rect 11149 23471 11207 23477
rect 13170 23468 13176 23480
rect 13228 23468 13234 23520
rect 13449 23511 13507 23517
rect 13449 23477 13461 23511
rect 13495 23508 13507 23511
rect 13906 23508 13912 23520
rect 13495 23480 13912 23508
rect 13495 23477 13507 23480
rect 13449 23471 13507 23477
rect 13906 23468 13912 23480
rect 13964 23468 13970 23520
rect 14090 23508 14096 23520
rect 14051 23480 14096 23508
rect 14090 23468 14096 23480
rect 14148 23468 14154 23520
rect 15470 23468 15476 23520
rect 15528 23508 15534 23520
rect 15933 23511 15991 23517
rect 15933 23508 15945 23511
rect 15528 23480 15945 23508
rect 15528 23468 15534 23480
rect 15933 23477 15945 23480
rect 15979 23508 15991 23511
rect 16853 23511 16911 23517
rect 16853 23508 16865 23511
rect 15979 23480 16865 23508
rect 15979 23477 15991 23480
rect 15933 23471 15991 23477
rect 16853 23477 16865 23480
rect 16899 23477 16911 23511
rect 17236 23508 17264 23616
rect 17313 23613 17325 23647
rect 17359 23613 17371 23647
rect 17313 23607 17371 23613
rect 18877 23647 18935 23653
rect 18877 23613 18889 23647
rect 18923 23644 18935 23647
rect 19426 23644 19432 23656
rect 18923 23616 19432 23644
rect 18923 23613 18935 23616
rect 18877 23607 18935 23613
rect 17328 23576 17356 23607
rect 19426 23604 19432 23616
rect 19484 23604 19490 23656
rect 20349 23579 20407 23585
rect 20349 23576 20361 23579
rect 17328 23548 20361 23576
rect 20349 23545 20361 23548
rect 20395 23545 20407 23579
rect 20349 23539 20407 23545
rect 18138 23508 18144 23520
rect 17236 23480 18144 23508
rect 16853 23471 16911 23477
rect 18138 23468 18144 23480
rect 18196 23468 18202 23520
rect 18322 23508 18328 23520
rect 18283 23480 18328 23508
rect 18322 23468 18328 23480
rect 18380 23468 18386 23520
rect 21910 23468 21916 23520
rect 21968 23508 21974 23520
rect 33873 23511 33931 23517
rect 33873 23508 33885 23511
rect 21968 23480 33885 23508
rect 21968 23468 21974 23480
rect 33873 23477 33885 23480
rect 33919 23477 33931 23511
rect 33873 23471 33931 23477
rect 34514 23468 34520 23520
rect 34572 23508 34578 23520
rect 38105 23511 38163 23517
rect 38105 23508 38117 23511
rect 34572 23480 38117 23508
rect 34572 23468 34578 23480
rect 38105 23477 38117 23480
rect 38151 23477 38163 23511
rect 38105 23471 38163 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1854 23264 1860 23316
rect 1912 23304 1918 23316
rect 6086 23304 6092 23316
rect 1912 23276 6092 23304
rect 1912 23264 1918 23276
rect 6086 23264 6092 23276
rect 6144 23264 6150 23316
rect 7763 23307 7821 23313
rect 7763 23273 7775 23307
rect 7809 23304 7821 23307
rect 10318 23304 10324 23316
rect 7809 23276 10324 23304
rect 7809 23273 7821 23276
rect 7763 23267 7821 23273
rect 10318 23264 10324 23276
rect 10376 23264 10382 23316
rect 12526 23304 12532 23316
rect 12487 23276 12532 23304
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 14550 23264 14556 23316
rect 14608 23304 14614 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14608 23276 14657 23304
rect 14608 23264 14614 23276
rect 14645 23273 14657 23276
rect 14691 23273 14703 23307
rect 20530 23304 20536 23316
rect 20491 23276 20536 23304
rect 14645 23267 14703 23273
rect 20530 23264 20536 23276
rect 20588 23264 20594 23316
rect 4065 23239 4123 23245
rect 4065 23205 4077 23239
rect 4111 23236 4123 23239
rect 5534 23236 5540 23248
rect 4111 23208 5540 23236
rect 4111 23205 4123 23208
rect 4065 23199 4123 23205
rect 5534 23196 5540 23208
rect 5592 23196 5598 23248
rect 8294 23196 8300 23248
rect 8352 23236 8358 23248
rect 17770 23236 17776 23248
rect 8352 23208 12112 23236
rect 8352 23196 8358 23208
rect 1581 23171 1639 23177
rect 1581 23137 1593 23171
rect 1627 23168 1639 23171
rect 2222 23168 2228 23180
rect 1627 23140 2228 23168
rect 1627 23137 1639 23140
rect 1581 23131 1639 23137
rect 2222 23128 2228 23140
rect 2280 23128 2286 23180
rect 5258 23128 5264 23180
rect 5316 23168 5322 23180
rect 5316 23140 8340 23168
rect 5316 23128 5322 23140
rect 3878 23060 3884 23112
rect 3936 23100 3942 23112
rect 3973 23103 4031 23109
rect 3973 23100 3985 23103
rect 3936 23072 3985 23100
rect 3936 23060 3942 23072
rect 3973 23069 3985 23072
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 4617 23103 4675 23109
rect 4617 23069 4629 23103
rect 4663 23100 4675 23103
rect 4706 23100 4712 23112
rect 4663 23072 4712 23100
rect 4663 23069 4675 23072
rect 4617 23063 4675 23069
rect 4706 23060 4712 23072
rect 4764 23100 4770 23112
rect 5442 23100 5448 23112
rect 4764 23072 5448 23100
rect 4764 23060 4770 23072
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 8021 23103 8079 23109
rect 8021 23069 8033 23103
rect 8067 23100 8079 23103
rect 8202 23100 8208 23112
rect 8067 23072 8208 23100
rect 8067 23069 8079 23072
rect 8021 23063 8079 23069
rect 8202 23060 8208 23072
rect 8260 23060 8266 23112
rect 8312 23100 8340 23140
rect 8478 23128 8484 23180
rect 8536 23168 8542 23180
rect 8536 23140 9904 23168
rect 8536 23128 8542 23140
rect 9876 23100 9904 23140
rect 10594 23128 10600 23180
rect 10652 23168 10658 23180
rect 10873 23171 10931 23177
rect 10873 23168 10885 23171
rect 10652 23140 10885 23168
rect 10652 23128 10658 23140
rect 10873 23137 10885 23140
rect 10919 23137 10931 23171
rect 10873 23131 10931 23137
rect 11146 23128 11152 23180
rect 11204 23168 11210 23180
rect 12084 23177 12112 23208
rect 15304 23208 17776 23236
rect 11885 23171 11943 23177
rect 11885 23168 11897 23171
rect 11204 23140 11897 23168
rect 11204 23128 11210 23140
rect 11885 23137 11897 23140
rect 11931 23137 11943 23171
rect 11885 23131 11943 23137
rect 12069 23171 12127 23177
rect 12069 23137 12081 23171
rect 12115 23137 12127 23171
rect 13078 23168 13084 23180
rect 13039 23140 13084 23168
rect 12069 23131 12127 23137
rect 13078 23128 13084 23140
rect 13136 23128 13142 23180
rect 13538 23168 13544 23180
rect 13499 23140 13544 23168
rect 13538 23128 13544 23140
rect 13596 23168 13602 23180
rect 13998 23168 14004 23180
rect 13596 23140 14004 23168
rect 13596 23128 13602 23140
rect 13998 23128 14004 23140
rect 14056 23128 14062 23180
rect 14090 23128 14096 23180
rect 14148 23168 14154 23180
rect 14148 23140 15240 23168
rect 14148 23128 14154 23140
rect 10689 23103 10747 23109
rect 10689 23100 10701 23103
rect 8312 23072 9076 23100
rect 9876 23072 10701 23100
rect 1857 23035 1915 23041
rect 1857 23001 1869 23035
rect 1903 23032 1915 23035
rect 2130 23032 2136 23044
rect 1903 23004 2136 23032
rect 1903 23001 1915 23004
rect 1857 22995 1915 23001
rect 2130 22992 2136 23004
rect 2188 22992 2194 23044
rect 4982 23032 4988 23044
rect 3082 23004 4988 23032
rect 4982 22992 4988 23004
rect 5040 22992 5046 23044
rect 5166 22992 5172 23044
rect 5224 23032 5230 23044
rect 5224 23004 6578 23032
rect 5224 22992 5230 23004
rect 3326 22964 3332 22976
rect 3287 22936 3332 22964
rect 3326 22924 3332 22936
rect 3384 22924 3390 22976
rect 4706 22964 4712 22976
rect 4667 22936 4712 22964
rect 4706 22924 4712 22936
rect 4764 22924 4770 22976
rect 5813 22967 5871 22973
rect 5813 22933 5825 22967
rect 5859 22964 5871 22967
rect 6178 22964 6184 22976
rect 5859 22936 6184 22964
rect 5859 22933 5871 22936
rect 5813 22927 5871 22933
rect 6178 22924 6184 22936
rect 6236 22924 6242 22976
rect 6273 22967 6331 22973
rect 6273 22933 6285 22967
rect 6319 22964 6331 22967
rect 8938 22964 8944 22976
rect 6319 22936 8944 22964
rect 6319 22933 6331 22936
rect 6273 22927 6331 22933
rect 8938 22924 8944 22936
rect 8996 22924 9002 22976
rect 9048 22964 9076 23072
rect 10689 23069 10701 23072
rect 10735 23069 10747 23103
rect 10689 23063 10747 23069
rect 13722 23060 13728 23112
rect 13780 23100 13786 23112
rect 15102 23100 15108 23112
rect 13780 23072 14964 23100
rect 15063 23072 15108 23100
rect 13780 23060 13786 23072
rect 9214 23032 9220 23044
rect 9176 23004 9220 23032
rect 9214 22992 9220 23004
rect 9272 22992 9278 23044
rect 9318 23035 9376 23041
rect 9318 23001 9330 23035
rect 9364 23032 9376 23035
rect 9858 23032 9864 23044
rect 9364 23004 9444 23032
rect 9819 23004 9864 23032
rect 9364 23001 9376 23004
rect 9318 22995 9376 23001
rect 9416 22964 9444 23004
rect 9858 22992 9864 23004
rect 9916 22992 9922 23044
rect 13170 22992 13176 23044
rect 13228 23032 13234 23044
rect 14826 23032 14832 23044
rect 13228 23004 13273 23032
rect 13740 23004 14832 23032
rect 13228 22992 13234 23004
rect 9048 22936 9444 22964
rect 11333 22967 11391 22973
rect 11333 22933 11345 22967
rect 11379 22964 11391 22967
rect 13740 22964 13768 23004
rect 14826 22992 14832 23004
rect 14884 22992 14890 23044
rect 11379 22936 13768 22964
rect 11379 22933 11391 22936
rect 11333 22927 11391 22933
rect 14090 22924 14096 22976
rect 14148 22964 14154 22976
rect 14274 22964 14280 22976
rect 14148 22936 14280 22964
rect 14148 22924 14154 22936
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 14936 22964 14964 23072
rect 15102 23060 15108 23072
rect 15160 23060 15166 23112
rect 15212 23032 15240 23140
rect 15304 23109 15332 23208
rect 17770 23196 17776 23208
rect 17828 23196 17834 23248
rect 15930 23128 15936 23180
rect 15988 23168 15994 23180
rect 16117 23171 16175 23177
rect 16117 23168 16129 23171
rect 15988 23140 16129 23168
rect 15988 23128 15994 23140
rect 16117 23137 16129 23140
rect 16163 23137 16175 23171
rect 18230 23168 18236 23180
rect 18191 23140 18236 23168
rect 16117 23131 16175 23137
rect 18230 23128 18236 23140
rect 18288 23128 18294 23180
rect 18322 23128 18328 23180
rect 18380 23168 18386 23180
rect 18417 23171 18475 23177
rect 18417 23168 18429 23171
rect 18380 23140 18429 23168
rect 18380 23128 18386 23140
rect 18417 23137 18429 23140
rect 18463 23137 18475 23171
rect 18417 23131 18475 23137
rect 20073 23171 20131 23177
rect 20073 23137 20085 23171
rect 20119 23168 20131 23171
rect 33226 23168 33232 23180
rect 20119 23140 33232 23168
rect 20119 23137 20131 23140
rect 20073 23131 20131 23137
rect 33226 23128 33232 23140
rect 33284 23128 33290 23180
rect 15289 23103 15347 23109
rect 15289 23069 15301 23103
rect 15335 23069 15347 23103
rect 17310 23100 17316 23112
rect 17271 23072 17316 23100
rect 15289 23063 15347 23069
rect 17310 23060 17316 23072
rect 17368 23060 17374 23112
rect 19242 23060 19248 23112
rect 19300 23100 19306 23112
rect 19889 23103 19947 23109
rect 19889 23100 19901 23103
rect 19300 23072 19901 23100
rect 19300 23060 19306 23072
rect 19889 23069 19901 23072
rect 19935 23069 19947 23103
rect 20714 23100 20720 23112
rect 20675 23072 20720 23100
rect 19889 23063 19947 23069
rect 20714 23060 20720 23072
rect 20772 23060 20778 23112
rect 16209 23035 16267 23041
rect 15212 23004 15976 23032
rect 15654 22964 15660 22976
rect 14936 22936 15660 22964
rect 15654 22924 15660 22936
rect 15712 22924 15718 22976
rect 15948 22964 15976 23004
rect 16209 23001 16221 23035
rect 16255 23001 16267 23035
rect 16758 23032 16764 23044
rect 16719 23004 16764 23032
rect 16209 22995 16267 23001
rect 16224 22964 16252 22995
rect 16758 22992 16764 23004
rect 16816 22992 16822 23044
rect 17402 22964 17408 22976
rect 15948 22936 16252 22964
rect 17363 22936 17408 22964
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 18874 22964 18880 22976
rect 18835 22936 18880 22964
rect 18874 22924 18880 22936
rect 18932 22964 18938 22976
rect 19429 22967 19487 22973
rect 19429 22964 19441 22967
rect 18932 22936 19441 22964
rect 18932 22924 18938 22936
rect 19429 22933 19441 22936
rect 19475 22933 19487 22967
rect 19429 22927 19487 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1765 22763 1823 22769
rect 1765 22729 1777 22763
rect 1811 22760 1823 22763
rect 1854 22760 1860 22772
rect 1811 22732 1860 22760
rect 1811 22729 1823 22732
rect 1765 22723 1823 22729
rect 1854 22720 1860 22732
rect 1912 22720 1918 22772
rect 2130 22720 2136 22772
rect 2188 22760 2194 22772
rect 3418 22760 3424 22772
rect 2188 22732 3424 22760
rect 2188 22720 2194 22732
rect 3418 22720 3424 22732
rect 3476 22760 3482 22772
rect 7745 22763 7803 22769
rect 3476 22732 5856 22760
rect 3476 22720 3482 22732
rect 3786 22692 3792 22704
rect 3726 22664 3792 22692
rect 3786 22652 3792 22664
rect 3844 22652 3850 22704
rect 5258 22692 5264 22704
rect 5219 22664 5264 22692
rect 5258 22652 5264 22664
rect 5316 22652 5322 22704
rect 1578 22624 1584 22636
rect 1539 22596 1584 22624
rect 1578 22584 1584 22596
rect 1636 22584 1642 22636
rect 2222 22624 2228 22636
rect 2183 22596 2228 22624
rect 2222 22584 2228 22596
rect 2280 22584 2286 22636
rect 4614 22624 4620 22636
rect 4575 22596 4620 22624
rect 4614 22584 4620 22596
rect 4672 22624 4678 22636
rect 4982 22624 4988 22636
rect 4672 22596 4988 22624
rect 4672 22584 4678 22596
rect 4982 22584 4988 22596
rect 5040 22584 5046 22636
rect 5828 22633 5856 22732
rect 7745 22729 7757 22763
rect 7791 22760 7803 22763
rect 7926 22760 7932 22772
rect 7791 22732 7932 22760
rect 7791 22729 7803 22732
rect 7745 22723 7803 22729
rect 7926 22720 7932 22732
rect 7984 22720 7990 22772
rect 8202 22720 8208 22772
rect 8260 22760 8266 22772
rect 9122 22760 9128 22772
rect 8260 22732 9128 22760
rect 8260 22720 8266 22732
rect 9122 22720 9128 22732
rect 9180 22760 9186 22772
rect 9180 22732 9444 22760
rect 9180 22720 9186 22732
rect 6178 22652 6184 22704
rect 6236 22692 6242 22704
rect 6641 22695 6699 22701
rect 6641 22692 6653 22695
rect 6236 22664 6653 22692
rect 6236 22652 6242 22664
rect 6641 22661 6653 22664
rect 6687 22661 6699 22695
rect 6641 22655 6699 22661
rect 6730 22652 6736 22704
rect 6788 22692 6794 22704
rect 6788 22664 6833 22692
rect 6788 22652 6794 22664
rect 6914 22652 6920 22704
rect 6972 22692 6978 22704
rect 7285 22695 7343 22701
rect 7285 22692 7297 22695
rect 6972 22664 7297 22692
rect 6972 22652 6978 22664
rect 7285 22661 7297 22664
rect 7331 22661 7343 22695
rect 7285 22655 7343 22661
rect 8938 22652 8944 22704
rect 8996 22692 9002 22704
rect 9217 22695 9275 22701
rect 9217 22692 9229 22695
rect 8996 22664 9229 22692
rect 8996 22652 9002 22664
rect 9217 22661 9229 22664
rect 9263 22661 9275 22695
rect 9416 22692 9444 22732
rect 9582 22720 9588 22772
rect 9640 22760 9646 22772
rect 9640 22720 9674 22760
rect 12986 22720 12992 22772
rect 13044 22760 13050 22772
rect 13044 22732 14872 22760
rect 13044 22720 13050 22732
rect 9646 22692 9674 22720
rect 9416 22664 9536 22692
rect 9646 22664 10824 22692
rect 9217 22655 9275 22661
rect 5353 22627 5411 22633
rect 5353 22593 5365 22627
rect 5399 22593 5411 22627
rect 5353 22587 5411 22593
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22593 5871 22627
rect 5813 22587 5871 22593
rect 2501 22559 2559 22565
rect 2501 22556 2513 22559
rect 2332 22528 2513 22556
rect 2332 22432 2360 22528
rect 2501 22525 2513 22528
rect 2547 22525 2559 22559
rect 5166 22556 5172 22568
rect 2501 22519 2559 22525
rect 3528 22528 5172 22556
rect 2314 22380 2320 22432
rect 2372 22380 2378 22432
rect 2590 22380 2596 22432
rect 2648 22420 2654 22432
rect 3528 22420 3556 22528
rect 5166 22516 5172 22528
rect 5224 22516 5230 22568
rect 3602 22448 3608 22500
rect 3660 22488 3666 22500
rect 4525 22491 4583 22497
rect 4525 22488 4537 22491
rect 3660 22460 4537 22488
rect 3660 22448 3666 22460
rect 4525 22457 4537 22460
rect 4571 22457 4583 22491
rect 5368 22488 5396 22587
rect 5828 22556 5856 22587
rect 8110 22584 8116 22636
rect 8168 22584 8174 22636
rect 9508 22633 9536 22664
rect 9493 22627 9551 22633
rect 9493 22593 9505 22627
rect 9539 22593 9551 22627
rect 9493 22587 9551 22593
rect 9582 22584 9588 22636
rect 9640 22624 9646 22636
rect 9950 22624 9956 22636
rect 9640 22596 9956 22624
rect 9640 22584 9646 22596
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 10134 22584 10140 22636
rect 10192 22624 10198 22636
rect 10689 22627 10747 22633
rect 10689 22624 10701 22627
rect 10192 22596 10701 22624
rect 10192 22584 10198 22596
rect 10689 22593 10701 22596
rect 10735 22593 10747 22627
rect 10796 22624 10824 22664
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 11149 22695 11207 22701
rect 11149 22692 11161 22695
rect 11112 22664 11161 22692
rect 11112 22652 11118 22664
rect 11149 22661 11161 22664
rect 11195 22692 11207 22695
rect 11422 22692 11428 22704
rect 11195 22664 11428 22692
rect 11195 22661 11207 22664
rect 11149 22655 11207 22661
rect 11422 22652 11428 22664
rect 11480 22652 11486 22704
rect 13814 22692 13820 22704
rect 13775 22664 13820 22692
rect 13814 22652 13820 22664
rect 13872 22652 13878 22704
rect 14844 22692 14872 22732
rect 14918 22720 14924 22772
rect 14976 22760 14982 22772
rect 19242 22760 19248 22772
rect 14976 22732 15608 22760
rect 19203 22732 19248 22760
rect 14976 22720 14982 22732
rect 15286 22692 15292 22704
rect 14844 22664 15292 22692
rect 15286 22652 15292 22664
rect 15344 22652 15350 22704
rect 15470 22692 15476 22704
rect 15431 22664 15476 22692
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 15580 22701 15608 22732
rect 19242 22720 19248 22732
rect 19300 22720 19306 22772
rect 15565 22695 15623 22701
rect 15565 22661 15577 22695
rect 15611 22661 15623 22695
rect 17402 22692 17408 22704
rect 17363 22664 17408 22692
rect 15565 22655 15623 22661
rect 17402 22652 17408 22664
rect 17460 22652 17466 22704
rect 17862 22652 17868 22704
rect 17920 22692 17926 22704
rect 20714 22692 20720 22704
rect 17920 22664 20720 22692
rect 17920 22652 17926 22664
rect 12710 22624 12716 22636
rect 10796 22596 12716 22624
rect 10689 22587 10747 22593
rect 12710 22584 12716 22596
rect 12768 22584 12774 22636
rect 12989 22627 13047 22633
rect 12989 22593 13001 22627
rect 13035 22624 13047 22627
rect 13078 22624 13084 22636
rect 13035 22596 13084 22624
rect 13035 22593 13047 22596
rect 12989 22587 13047 22593
rect 13078 22584 13084 22596
rect 13136 22584 13142 22636
rect 17954 22584 17960 22636
rect 18012 22624 18018 22636
rect 18233 22627 18291 22633
rect 18233 22624 18245 22627
rect 18012 22596 18245 22624
rect 18012 22584 18018 22596
rect 18233 22593 18245 22596
rect 18279 22593 18291 22627
rect 18233 22587 18291 22593
rect 18414 22584 18420 22636
rect 18472 22624 18478 22636
rect 19168 22633 19196 22664
rect 20714 22652 20720 22664
rect 20772 22652 20778 22704
rect 18693 22627 18751 22633
rect 18693 22624 18705 22627
rect 18472 22596 18705 22624
rect 18472 22584 18478 22596
rect 18693 22593 18705 22596
rect 18739 22593 18751 22627
rect 18693 22587 18751 22593
rect 19153 22627 19211 22633
rect 19153 22593 19165 22627
rect 19199 22593 19211 22627
rect 19153 22587 19211 22593
rect 19242 22584 19248 22636
rect 19300 22624 19306 22636
rect 21174 22624 21180 22636
rect 19300 22596 21180 22624
rect 19300 22584 19306 22596
rect 21174 22584 21180 22596
rect 21232 22584 21238 22636
rect 21450 22624 21456 22636
rect 21411 22596 21456 22624
rect 21450 22584 21456 22596
rect 21508 22584 21514 22636
rect 5828 22528 7788 22556
rect 7098 22488 7104 22500
rect 5368 22460 7104 22488
rect 4525 22451 4583 22457
rect 7098 22448 7104 22460
rect 7156 22448 7162 22500
rect 2648 22392 3556 22420
rect 3973 22423 4031 22429
rect 2648 22380 2654 22392
rect 3973 22389 3985 22423
rect 4019 22420 4031 22423
rect 5810 22420 5816 22432
rect 4019 22392 5816 22420
rect 4019 22389 4031 22392
rect 3973 22383 4031 22389
rect 5810 22380 5816 22392
rect 5868 22380 5874 22432
rect 5905 22423 5963 22429
rect 5905 22389 5917 22423
rect 5951 22420 5963 22423
rect 7650 22420 7656 22432
rect 5951 22392 7656 22420
rect 5951 22389 5963 22392
rect 5905 22383 5963 22389
rect 7650 22380 7656 22392
rect 7708 22380 7714 22432
rect 7760 22420 7788 22528
rect 9766 22516 9772 22568
rect 9824 22556 9830 22568
rect 10505 22559 10563 22565
rect 10505 22556 10517 22559
rect 9824 22528 10517 22556
rect 9824 22516 9830 22528
rect 10505 22525 10517 22528
rect 10551 22556 10563 22559
rect 10551 22528 10824 22556
rect 10551 22525 10563 22528
rect 10505 22519 10563 22525
rect 10796 22500 10824 22528
rect 10962 22516 10968 22568
rect 11020 22556 11026 22568
rect 11701 22559 11759 22565
rect 11701 22556 11713 22559
rect 11020 22528 11713 22556
rect 11020 22516 11026 22528
rect 11701 22525 11713 22528
rect 11747 22525 11759 22559
rect 11882 22556 11888 22568
rect 11843 22528 11888 22556
rect 11701 22519 11759 22525
rect 11882 22516 11888 22528
rect 11940 22516 11946 22568
rect 13722 22556 13728 22568
rect 13683 22528 13728 22556
rect 13722 22516 13728 22528
rect 13780 22516 13786 22568
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 17221 22559 17279 22565
rect 17221 22556 17233 22559
rect 16816 22528 17233 22556
rect 16816 22516 16822 22528
rect 17221 22525 17233 22528
rect 17267 22525 17279 22559
rect 17221 22519 17279 22525
rect 10778 22448 10784 22500
rect 10836 22448 10842 22500
rect 11974 22448 11980 22500
rect 12032 22488 12038 22500
rect 12069 22491 12127 22497
rect 12069 22488 12081 22491
rect 12032 22460 12081 22488
rect 12032 22448 12038 22460
rect 12069 22457 12081 22460
rect 12115 22457 12127 22491
rect 12069 22451 12127 22457
rect 14277 22491 14335 22497
rect 14277 22457 14289 22491
rect 14323 22488 14335 22491
rect 16025 22491 16083 22497
rect 16025 22488 16037 22491
rect 14323 22460 16037 22488
rect 14323 22457 14335 22460
rect 14277 22451 14335 22457
rect 16025 22457 16037 22460
rect 16071 22488 16083 22491
rect 17034 22488 17040 22500
rect 16071 22460 17040 22488
rect 16071 22457 16083 22460
rect 16025 22451 16083 22457
rect 17034 22448 17040 22460
rect 17092 22448 17098 22500
rect 17236 22488 17264 22519
rect 17402 22516 17408 22568
rect 17460 22556 17466 22568
rect 17497 22559 17555 22565
rect 17497 22556 17509 22559
rect 17460 22528 17509 22556
rect 17460 22516 17466 22528
rect 17497 22525 17509 22528
rect 17543 22525 17555 22559
rect 18046 22556 18052 22568
rect 17959 22528 18052 22556
rect 17497 22519 17555 22525
rect 18046 22516 18052 22528
rect 18104 22556 18110 22568
rect 18598 22556 18604 22568
rect 18104 22528 18604 22556
rect 18104 22516 18110 22528
rect 18598 22516 18604 22528
rect 18656 22516 18662 22568
rect 20625 22559 20683 22565
rect 20625 22525 20637 22559
rect 20671 22525 20683 22559
rect 20625 22519 20683 22525
rect 20640 22488 20668 22519
rect 20806 22516 20812 22568
rect 20864 22556 20870 22568
rect 30466 22556 30472 22568
rect 20864 22528 30472 22556
rect 20864 22516 20870 22528
rect 30466 22516 30472 22528
rect 30524 22516 30530 22568
rect 21269 22491 21327 22497
rect 21269 22488 21281 22491
rect 17236 22460 20576 22488
rect 20640 22460 21281 22488
rect 9766 22420 9772 22432
rect 7760 22392 9772 22420
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 9858 22380 9864 22432
rect 9916 22420 9922 22432
rect 12986 22420 12992 22432
rect 9916 22392 12992 22420
rect 9916 22380 9922 22392
rect 12986 22380 12992 22392
rect 13044 22380 13050 22432
rect 13173 22423 13231 22429
rect 13173 22389 13185 22423
rect 13219 22420 13231 22423
rect 15194 22420 15200 22432
rect 13219 22392 15200 22420
rect 13219 22389 13231 22392
rect 13173 22383 13231 22389
rect 15194 22380 15200 22392
rect 15252 22380 15258 22432
rect 15286 22380 15292 22432
rect 15344 22420 15350 22432
rect 18782 22420 18788 22432
rect 15344 22392 18788 22420
rect 15344 22380 15350 22392
rect 18782 22380 18788 22392
rect 18840 22380 18846 22432
rect 20438 22420 20444 22432
rect 20399 22392 20444 22420
rect 20438 22380 20444 22392
rect 20496 22380 20502 22432
rect 20548 22420 20576 22460
rect 21269 22457 21281 22460
rect 21315 22457 21327 22491
rect 21269 22451 21327 22457
rect 33318 22420 33324 22432
rect 20548 22392 33324 22420
rect 33318 22380 33324 22392
rect 33376 22380 33382 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 2958 22176 2964 22228
rect 3016 22216 3022 22228
rect 3157 22219 3215 22225
rect 3157 22216 3169 22219
rect 3016 22188 3169 22216
rect 3016 22176 3022 22188
rect 3157 22185 3169 22188
rect 3203 22216 3215 22219
rect 4062 22216 4068 22228
rect 3203 22188 4068 22216
rect 3203 22185 3215 22188
rect 3157 22179 3215 22185
rect 4062 22176 4068 22188
rect 4120 22176 4126 22228
rect 5258 22176 5264 22228
rect 5316 22216 5322 22228
rect 5442 22216 5448 22228
rect 5316 22188 5448 22216
rect 5316 22176 5322 22188
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 8315 22219 8373 22225
rect 8315 22185 8327 22219
rect 8361 22216 8373 22219
rect 9030 22216 9036 22228
rect 8361 22188 9036 22216
rect 8361 22185 8373 22188
rect 8315 22179 8373 22185
rect 9030 22176 9036 22188
rect 9088 22216 9094 22228
rect 9214 22216 9220 22228
rect 9088 22188 9220 22216
rect 9088 22176 9094 22188
rect 9214 22176 9220 22188
rect 9272 22176 9278 22228
rect 12526 22176 12532 22228
rect 12584 22216 12590 22228
rect 12897 22219 12955 22225
rect 12897 22216 12909 22219
rect 12584 22188 12909 22216
rect 12584 22176 12590 22188
rect 12897 22185 12909 22188
rect 12943 22185 12955 22219
rect 12897 22179 12955 22185
rect 13446 22176 13452 22228
rect 13504 22216 13510 22228
rect 18874 22216 18880 22228
rect 13504 22188 18880 22216
rect 13504 22176 13510 22188
rect 18874 22176 18880 22188
rect 18932 22176 18938 22228
rect 6825 22151 6883 22157
rect 6825 22117 6837 22151
rect 6871 22148 6883 22151
rect 7282 22148 7288 22160
rect 6871 22120 7288 22148
rect 6871 22117 6883 22120
rect 6825 22111 6883 22117
rect 7282 22108 7288 22120
rect 7340 22108 7346 22160
rect 9306 22108 9312 22160
rect 9364 22148 9370 22160
rect 13538 22148 13544 22160
rect 9364 22120 13544 22148
rect 9364 22108 9370 22120
rect 13538 22108 13544 22120
rect 13596 22108 13602 22160
rect 14200 22120 14780 22148
rect 2130 22040 2136 22092
rect 2188 22080 2194 22092
rect 3421 22083 3479 22089
rect 3421 22080 3433 22083
rect 2188 22052 3433 22080
rect 2188 22040 2194 22052
rect 3421 22049 3433 22052
rect 3467 22080 3479 22083
rect 4522 22080 4528 22092
rect 3467 22052 4528 22080
rect 3467 22049 3479 22052
rect 3421 22043 3479 22049
rect 4522 22040 4528 22052
rect 4580 22080 4586 22092
rect 4617 22083 4675 22089
rect 4617 22080 4629 22083
rect 4580 22052 4629 22080
rect 4580 22040 4586 22052
rect 4617 22049 4629 22052
rect 4663 22049 4675 22083
rect 4617 22043 4675 22049
rect 5534 22040 5540 22092
rect 5592 22080 5598 22092
rect 5592 22052 7236 22080
rect 5592 22040 5598 22052
rect 3878 21972 3884 22024
rect 3936 22012 3942 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3936 21984 3985 22012
rect 3936 21972 3942 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 7208 21998 7236 22052
rect 8938 22040 8944 22092
rect 8996 22080 9002 22092
rect 9582 22080 9588 22092
rect 8996 22052 9588 22080
rect 8996 22040 9002 22052
rect 9582 22040 9588 22052
rect 9640 22040 9646 22092
rect 11238 22040 11244 22092
rect 11296 22080 11302 22092
rect 11425 22083 11483 22089
rect 11425 22080 11437 22083
rect 11296 22052 11437 22080
rect 11296 22040 11302 22052
rect 11425 22049 11437 22052
rect 11471 22080 11483 22083
rect 11698 22080 11704 22092
rect 11471 22052 11704 22080
rect 11471 22049 11483 22052
rect 11425 22043 11483 22049
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 11882 22040 11888 22092
rect 11940 22080 11946 22092
rect 12713 22083 12771 22089
rect 12713 22080 12725 22083
rect 11940 22052 12725 22080
rect 11940 22040 11946 22052
rect 12713 22049 12725 22052
rect 12759 22049 12771 22083
rect 12713 22043 12771 22049
rect 13630 22040 13636 22092
rect 13688 22080 13694 22092
rect 14200 22080 14228 22120
rect 14366 22080 14372 22092
rect 13688 22052 14228 22080
rect 14327 22052 14372 22080
rect 13688 22040 13694 22052
rect 14366 22040 14372 22052
rect 14424 22040 14430 22092
rect 14642 22080 14648 22092
rect 14603 22052 14648 22080
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 14752 22080 14780 22120
rect 15948 22120 18552 22148
rect 15948 22080 15976 22120
rect 16114 22080 16120 22092
rect 14752 22052 15976 22080
rect 16075 22052 16120 22080
rect 16114 22040 16120 22052
rect 16172 22040 16178 22092
rect 16761 22083 16819 22089
rect 16761 22049 16773 22083
rect 16807 22080 16819 22083
rect 18414 22080 18420 22092
rect 16807 22052 18420 22080
rect 16807 22049 16819 22052
rect 16761 22043 16819 22049
rect 18414 22040 18420 22052
rect 18472 22040 18478 22092
rect 18524 22080 18552 22120
rect 18690 22080 18696 22092
rect 18524 22052 18696 22080
rect 18690 22040 18696 22052
rect 18748 22040 18754 22092
rect 18874 22080 18880 22092
rect 18835 22052 18880 22080
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 21910 22080 21916 22092
rect 21871 22052 21916 22080
rect 21910 22040 21916 22052
rect 21968 22040 21974 22092
rect 8573 22015 8631 22021
rect 3973 21975 4031 21981
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 8619 21984 9168 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 2590 21904 2596 21956
rect 2648 21904 2654 21956
rect 1394 21836 1400 21888
rect 1452 21876 1458 21888
rect 1673 21879 1731 21885
rect 1673 21876 1685 21879
rect 1452 21848 1685 21876
rect 1452 21836 1458 21848
rect 1673 21845 1685 21848
rect 1719 21845 1731 21879
rect 1673 21839 1731 21845
rect 1854 21836 1860 21888
rect 1912 21876 1918 21888
rect 3988 21876 4016 21975
rect 9140 21956 9168 21984
rect 10410 21972 10416 22024
rect 10468 22012 10474 22024
rect 10468 21984 11008 22012
rect 10468 21972 10474 21984
rect 4246 21904 4252 21956
rect 4304 21944 4310 21956
rect 4798 21944 4804 21956
rect 4304 21916 4804 21944
rect 4304 21904 4310 21916
rect 4798 21904 4804 21916
rect 4856 21944 4862 21956
rect 4893 21947 4951 21953
rect 4893 21944 4905 21947
rect 4856 21916 4905 21944
rect 4856 21904 4862 21916
rect 4893 21913 4905 21916
rect 4939 21913 4951 21947
rect 4893 21907 4951 21913
rect 5350 21904 5356 21956
rect 5408 21904 5414 21956
rect 9122 21944 9128 21956
rect 9083 21916 9128 21944
rect 9122 21904 9128 21916
rect 9180 21904 9186 21956
rect 10873 21947 10931 21953
rect 10873 21913 10885 21947
rect 10919 21913 10931 21947
rect 10873 21907 10931 21913
rect 1912 21848 4016 21876
rect 4065 21879 4123 21885
rect 1912 21836 1918 21848
rect 4065 21845 4077 21879
rect 4111 21876 4123 21879
rect 5810 21876 5816 21888
rect 4111 21848 5816 21876
rect 4111 21845 4123 21848
rect 4065 21839 4123 21845
rect 5810 21836 5816 21848
rect 5868 21836 5874 21888
rect 6270 21836 6276 21888
rect 6328 21876 6334 21888
rect 6365 21879 6423 21885
rect 6365 21876 6377 21879
rect 6328 21848 6377 21876
rect 6328 21836 6334 21848
rect 6365 21845 6377 21848
rect 6411 21876 6423 21879
rect 6638 21876 6644 21888
rect 6411 21848 6644 21876
rect 6411 21845 6423 21848
rect 6365 21839 6423 21845
rect 6638 21836 6644 21848
rect 6696 21836 6702 21888
rect 6822 21836 6828 21888
rect 6880 21876 6886 21888
rect 10888 21876 10916 21907
rect 6880 21848 10916 21876
rect 10980 21876 11008 21984
rect 12342 21972 12348 22024
rect 12400 22012 12406 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12400 21984 12541 22012
rect 12400 21972 12406 21984
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 15102 21972 15108 22024
rect 15160 22012 15166 22024
rect 15657 22015 15715 22021
rect 15657 22012 15669 22015
rect 15160 21984 15669 22012
rect 15160 21972 15166 21984
rect 15657 21981 15669 21984
rect 15703 21981 15715 22015
rect 15657 21975 15715 21981
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 21981 16359 22015
rect 17494 22012 17500 22024
rect 17455 21984 17500 22012
rect 16301 21975 16359 21981
rect 11517 21947 11575 21953
rect 11517 21944 11529 21947
rect 11348 21916 11529 21944
rect 11348 21876 11376 21916
rect 11517 21913 11529 21916
rect 11563 21913 11575 21947
rect 12066 21944 12072 21956
rect 12027 21916 12072 21944
rect 11517 21907 11575 21913
rect 12066 21904 12072 21916
rect 12124 21904 12130 21956
rect 12250 21904 12256 21956
rect 12308 21944 12314 21956
rect 13814 21944 13820 21956
rect 12308 21916 13820 21944
rect 12308 21904 12314 21916
rect 13814 21904 13820 21916
rect 13872 21904 13878 21956
rect 14182 21904 14188 21956
rect 14240 21944 14246 21956
rect 14461 21947 14519 21953
rect 14461 21944 14473 21947
rect 14240 21916 14473 21944
rect 14240 21904 14246 21916
rect 14461 21913 14473 21916
rect 14507 21913 14519 21947
rect 14461 21907 14519 21913
rect 14550 21904 14556 21956
rect 14608 21944 14614 21956
rect 16316 21944 16344 21975
rect 17494 21972 17500 21984
rect 17552 21972 17558 22024
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 19613 22015 19671 22021
rect 19613 22012 19625 22015
rect 19392 21984 19625 22012
rect 19392 21972 19398 21984
rect 19613 21981 19625 21984
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 20162 21972 20168 22024
rect 20220 22012 20226 22024
rect 20257 22015 20315 22021
rect 20257 22012 20269 22015
rect 20220 21984 20269 22012
rect 20220 21972 20226 21984
rect 20257 21981 20269 21984
rect 20303 21981 20315 22015
rect 38286 22012 38292 22024
rect 38247 21984 38292 22012
rect 20257 21975 20315 21981
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 14608 21916 16344 21944
rect 14608 21904 14614 21916
rect 18046 21904 18052 21956
rect 18104 21944 18110 21956
rect 18322 21953 18328 21956
rect 18222 21947 18280 21953
rect 18222 21944 18234 21947
rect 18104 21916 18234 21944
rect 18104 21904 18110 21916
rect 18222 21913 18234 21916
rect 18268 21913 18280 21947
rect 18222 21907 18280 21913
rect 18318 21907 18328 21953
rect 18380 21944 18386 21956
rect 18380 21916 18418 21944
rect 18322 21904 18328 21907
rect 18380 21904 18386 21916
rect 18690 21904 18696 21956
rect 18748 21944 18754 21956
rect 21266 21944 21272 21956
rect 18748 21916 21272 21944
rect 18748 21904 18754 21916
rect 21266 21904 21272 21916
rect 21324 21904 21330 21956
rect 21818 21944 21824 21956
rect 21779 21916 21824 21944
rect 21818 21904 21824 21916
rect 21876 21904 21882 21956
rect 10980 21848 11376 21876
rect 6880 21836 6886 21848
rect 13538 21836 13544 21888
rect 13596 21876 13602 21888
rect 15473 21879 15531 21885
rect 15473 21876 15485 21879
rect 13596 21848 15485 21876
rect 13596 21836 13602 21848
rect 15473 21845 15485 21848
rect 15519 21845 15531 21879
rect 15473 21839 15531 21845
rect 17681 21879 17739 21885
rect 17681 21845 17693 21879
rect 17727 21876 17739 21879
rect 17954 21876 17960 21888
rect 17727 21848 17960 21876
rect 17727 21845 17739 21848
rect 17681 21839 17739 21845
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 18966 21836 18972 21888
rect 19024 21876 19030 21888
rect 19521 21879 19579 21885
rect 19521 21876 19533 21879
rect 19024 21848 19533 21876
rect 19024 21836 19030 21848
rect 19521 21845 19533 21848
rect 19567 21845 19579 21879
rect 19521 21839 19579 21845
rect 19978 21836 19984 21888
rect 20036 21876 20042 21888
rect 20073 21879 20131 21885
rect 20073 21876 20085 21879
rect 20036 21848 20085 21876
rect 20036 21836 20042 21848
rect 20073 21845 20085 21848
rect 20119 21845 20131 21879
rect 20073 21839 20131 21845
rect 32214 21836 32220 21888
rect 32272 21876 32278 21888
rect 38105 21879 38163 21885
rect 38105 21876 38117 21879
rect 32272 21848 38117 21876
rect 32272 21836 32278 21848
rect 38105 21845 38117 21848
rect 38151 21845 38163 21879
rect 38105 21839 38163 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 4246 21672 4252 21684
rect 4207 21644 4252 21672
rect 4246 21632 4252 21644
rect 4304 21632 4310 21684
rect 7285 21675 7343 21681
rect 4448 21644 7236 21672
rect 2038 21564 2044 21616
rect 2096 21604 2102 21616
rect 2096 21576 2162 21604
rect 2096 21564 2102 21576
rect 3234 21564 3240 21616
rect 3292 21604 3298 21616
rect 3329 21607 3387 21613
rect 3329 21604 3341 21607
rect 3292 21576 3341 21604
rect 3292 21564 3298 21576
rect 3329 21573 3341 21576
rect 3375 21604 3387 21607
rect 4448 21604 4476 21644
rect 3375 21576 4476 21604
rect 5721 21607 5779 21613
rect 3375 21573 3387 21576
rect 3329 21567 3387 21573
rect 5721 21573 5733 21607
rect 5767 21604 5779 21607
rect 6454 21604 6460 21616
rect 5767 21576 6460 21604
rect 5767 21573 5779 21576
rect 5721 21567 5779 21573
rect 6454 21564 6460 21576
rect 6512 21564 6518 21616
rect 3694 21496 3700 21548
rect 3752 21536 3758 21548
rect 3752 21508 4646 21536
rect 3752 21496 3758 21508
rect 6178 21496 6184 21548
rect 6236 21536 6242 21548
rect 7101 21539 7159 21545
rect 7101 21536 7113 21539
rect 6236 21508 7113 21536
rect 6236 21496 6242 21508
rect 7101 21505 7113 21508
rect 7147 21505 7159 21539
rect 7101 21499 7159 21505
rect 1581 21471 1639 21477
rect 1581 21437 1593 21471
rect 1627 21468 1639 21471
rect 2130 21468 2136 21480
rect 1627 21440 2136 21468
rect 1627 21437 1639 21440
rect 1581 21431 1639 21437
rect 2130 21428 2136 21440
rect 2188 21428 2194 21480
rect 3605 21471 3663 21477
rect 3605 21468 3617 21471
rect 2240 21440 3617 21468
rect 2240 21412 2268 21440
rect 3605 21437 3617 21440
rect 3651 21437 3663 21471
rect 5997 21471 6055 21477
rect 5997 21468 6009 21471
rect 3605 21431 3663 21437
rect 4632 21440 6009 21468
rect 4632 21412 4660 21440
rect 5997 21437 6009 21440
rect 6043 21437 6055 21471
rect 7208 21468 7236 21644
rect 7285 21641 7297 21675
rect 7331 21672 7343 21675
rect 8294 21672 8300 21684
rect 7331 21644 8300 21672
rect 7331 21641 7343 21644
rect 7285 21635 7343 21641
rect 8294 21632 8300 21644
rect 8352 21632 8358 21684
rect 8478 21632 8484 21684
rect 8536 21672 8542 21684
rect 10781 21675 10839 21681
rect 8536 21644 9536 21672
rect 8536 21632 8542 21644
rect 7466 21564 7472 21616
rect 7524 21604 7530 21616
rect 7524 21576 8050 21604
rect 7524 21564 7530 21576
rect 9508 21536 9536 21644
rect 10781 21641 10793 21675
rect 10827 21672 10839 21675
rect 12250 21672 12256 21684
rect 10827 21644 12256 21672
rect 10827 21641 10839 21644
rect 10781 21635 10839 21641
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 12897 21675 12955 21681
rect 12897 21641 12909 21675
rect 12943 21672 12955 21675
rect 16850 21672 16856 21684
rect 12943 21644 16856 21672
rect 12943 21641 12955 21644
rect 12897 21635 12955 21641
rect 16850 21632 16856 21644
rect 16908 21632 16914 21684
rect 17494 21632 17500 21684
rect 17552 21672 17558 21684
rect 18141 21675 18199 21681
rect 18141 21672 18153 21675
rect 17552 21644 18153 21672
rect 17552 21632 17558 21644
rect 18141 21641 18153 21644
rect 18187 21641 18199 21675
rect 20162 21672 20168 21684
rect 20123 21644 20168 21672
rect 18141 21635 18199 21641
rect 20162 21632 20168 21644
rect 20220 21632 20226 21684
rect 21269 21675 21327 21681
rect 21269 21641 21281 21675
rect 21315 21672 21327 21675
rect 21818 21672 21824 21684
rect 21315 21644 21824 21672
rect 21315 21641 21327 21644
rect 21269 21635 21327 21641
rect 21818 21632 21824 21644
rect 21876 21632 21882 21684
rect 29457 21675 29515 21681
rect 29457 21641 29469 21675
rect 29503 21672 29515 21675
rect 33134 21672 33140 21684
rect 29503 21644 33140 21672
rect 29503 21641 29515 21644
rect 29457 21635 29515 21641
rect 33134 21632 33140 21644
rect 33192 21632 33198 21684
rect 10134 21604 10140 21616
rect 10095 21576 10140 21604
rect 10134 21564 10140 21576
rect 10192 21564 10198 21616
rect 14458 21564 14464 21616
rect 14516 21604 14522 21616
rect 14553 21607 14611 21613
rect 14553 21604 14565 21607
rect 14516 21576 14565 21604
rect 14516 21564 14522 21576
rect 14553 21573 14565 21576
rect 14599 21573 14611 21607
rect 14553 21567 14611 21573
rect 14645 21607 14703 21613
rect 14645 21573 14657 21607
rect 14691 21604 14703 21607
rect 16942 21604 16948 21616
rect 14691 21576 16948 21604
rect 14691 21573 14703 21576
rect 14645 21567 14703 21573
rect 16942 21564 16948 21576
rect 17000 21564 17006 21616
rect 17126 21604 17132 21616
rect 17052 21576 17132 21604
rect 10045 21539 10103 21545
rect 9508 21508 9674 21536
rect 8478 21468 8484 21480
rect 7208 21440 8484 21468
rect 5997 21431 6055 21437
rect 8478 21428 8484 21440
rect 8536 21428 8542 21480
rect 8846 21428 8852 21480
rect 8904 21468 8910 21480
rect 9214 21468 9220 21480
rect 8904 21440 9220 21468
rect 8904 21428 8910 21440
rect 9214 21428 9220 21440
rect 9272 21428 9278 21480
rect 9493 21471 9551 21477
rect 9493 21468 9505 21471
rect 9416 21440 9505 21468
rect 2222 21360 2228 21412
rect 2280 21360 2286 21412
rect 4614 21360 4620 21412
rect 4672 21360 4678 21412
rect 7098 21292 7104 21344
rect 7156 21332 7162 21344
rect 7745 21335 7803 21341
rect 7745 21332 7757 21335
rect 7156 21304 7757 21332
rect 7156 21292 7162 21304
rect 7745 21301 7757 21304
rect 7791 21332 7803 21335
rect 8478 21332 8484 21344
rect 7791 21304 8484 21332
rect 7791 21301 7803 21304
rect 7745 21295 7803 21301
rect 8478 21292 8484 21304
rect 8536 21292 8542 21344
rect 9122 21292 9128 21344
rect 9180 21332 9186 21344
rect 9416 21332 9444 21440
rect 9493 21437 9505 21440
rect 9539 21437 9551 21471
rect 9646 21468 9674 21508
rect 10045 21505 10057 21539
rect 10091 21536 10103 21539
rect 10318 21536 10324 21548
rect 10091 21508 10324 21536
rect 10091 21505 10103 21508
rect 10045 21499 10103 21505
rect 10318 21496 10324 21508
rect 10376 21496 10382 21548
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21536 10747 21539
rect 12802 21536 12808 21548
rect 10735 21508 12808 21536
rect 10735 21505 10747 21508
rect 10689 21499 10747 21505
rect 10704 21468 10732 21499
rect 12802 21496 12808 21508
rect 12860 21496 12866 21548
rect 13354 21536 13360 21548
rect 13315 21508 13360 21536
rect 13354 21496 13360 21508
rect 13412 21496 13418 21548
rect 13998 21536 14004 21548
rect 13959 21508 14004 21536
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 15838 21536 15844 21548
rect 15799 21508 15844 21536
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 16850 21536 16856 21548
rect 16811 21508 16856 21536
rect 16850 21496 16856 21508
rect 16908 21496 16914 21548
rect 17052 21545 17080 21576
rect 17126 21564 17132 21576
rect 17184 21564 17190 21616
rect 18966 21604 18972 21616
rect 18927 21576 18972 21604
rect 18966 21564 18972 21576
rect 19024 21564 19030 21616
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 18138 21496 18144 21548
rect 18196 21536 18202 21548
rect 18325 21539 18383 21545
rect 18325 21536 18337 21539
rect 18196 21508 18337 21536
rect 18196 21496 18202 21508
rect 18325 21505 18337 21508
rect 18371 21505 18383 21539
rect 18325 21499 18383 21505
rect 19981 21539 20039 21545
rect 19981 21505 19993 21539
rect 20027 21505 20039 21539
rect 21174 21536 21180 21548
rect 21087 21508 21180 21536
rect 19981 21499 20039 21505
rect 9646 21440 10732 21468
rect 12253 21471 12311 21477
rect 9493 21431 9551 21437
rect 12253 21437 12265 21471
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 9582 21360 9588 21412
rect 9640 21400 9646 21412
rect 11882 21400 11888 21412
rect 9640 21372 11888 21400
rect 9640 21360 9646 21372
rect 11882 21360 11888 21372
rect 11940 21360 11946 21412
rect 9180 21304 9444 21332
rect 12268 21332 12296 21431
rect 13262 21428 13268 21480
rect 13320 21468 13326 21480
rect 15654 21468 15660 21480
rect 13320 21440 15056 21468
rect 15615 21440 15660 21468
rect 13320 21428 13326 21440
rect 13449 21403 13507 21409
rect 13449 21369 13461 21403
rect 13495 21400 13507 21403
rect 14550 21400 14556 21412
rect 13495 21372 14556 21400
rect 13495 21369 13507 21372
rect 13449 21363 13507 21369
rect 14550 21360 14556 21372
rect 14608 21360 14614 21412
rect 14918 21332 14924 21344
rect 12268 21304 14924 21332
rect 9180 21292 9186 21304
rect 14918 21292 14924 21304
rect 14976 21292 14982 21344
rect 15028 21332 15056 21440
rect 15654 21428 15660 21440
rect 15712 21428 15718 21480
rect 18414 21428 18420 21480
rect 18472 21468 18478 21480
rect 18877 21471 18935 21477
rect 18877 21468 18889 21471
rect 18472 21440 18889 21468
rect 18472 21428 18478 21440
rect 18877 21437 18889 21440
rect 18923 21437 18935 21471
rect 19334 21468 19340 21480
rect 19247 21440 19340 21468
rect 18877 21431 18935 21437
rect 19334 21428 19340 21440
rect 19392 21468 19398 21480
rect 19996 21468 20024 21499
rect 21174 21496 21180 21508
rect 21232 21536 21238 21548
rect 21358 21536 21364 21548
rect 21232 21508 21364 21536
rect 21232 21496 21238 21508
rect 21358 21496 21364 21508
rect 21416 21496 21422 21548
rect 21542 21496 21548 21548
rect 21600 21536 21606 21548
rect 22833 21539 22891 21545
rect 22833 21536 22845 21539
rect 21600 21508 22845 21536
rect 21600 21496 21606 21508
rect 22833 21505 22845 21508
rect 22879 21505 22891 21539
rect 22833 21499 22891 21505
rect 25314 21496 25320 21548
rect 25372 21536 25378 21548
rect 29365 21539 29423 21545
rect 29365 21536 29377 21539
rect 25372 21508 29377 21536
rect 25372 21496 25378 21508
rect 29365 21505 29377 21508
rect 29411 21505 29423 21539
rect 29365 21499 29423 21505
rect 30745 21539 30803 21545
rect 30745 21505 30757 21539
rect 30791 21536 30803 21539
rect 34514 21536 34520 21548
rect 30791 21508 34520 21536
rect 30791 21505 30803 21508
rect 30745 21499 30803 21505
rect 34514 21496 34520 21508
rect 34572 21496 34578 21548
rect 19392 21440 20024 21468
rect 19392 21428 19398 21440
rect 21910 21428 21916 21480
rect 21968 21468 21974 21480
rect 22005 21471 22063 21477
rect 22005 21468 22017 21471
rect 21968 21440 22017 21468
rect 21968 21428 21974 21440
rect 22005 21437 22017 21440
rect 22051 21437 22063 21471
rect 22005 21431 22063 21437
rect 19352 21400 19380 21428
rect 15764 21372 19380 21400
rect 19429 21403 19487 21409
rect 15764 21332 15792 21372
rect 19429 21369 19441 21403
rect 19475 21400 19487 21403
rect 20070 21400 20076 21412
rect 19475 21372 20076 21400
rect 19475 21369 19487 21372
rect 19429 21363 19487 21369
rect 20070 21360 20076 21372
rect 20128 21400 20134 21412
rect 35618 21400 35624 21412
rect 20128 21372 35624 21400
rect 20128 21360 20134 21372
rect 35618 21360 35624 21372
rect 35676 21360 35682 21412
rect 15028 21304 15792 21332
rect 16301 21335 16359 21341
rect 16301 21301 16313 21335
rect 16347 21332 16359 21335
rect 16850 21332 16856 21344
rect 16347 21304 16856 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 16850 21292 16856 21304
rect 16908 21332 16914 21344
rect 17221 21335 17279 21341
rect 17221 21332 17233 21335
rect 16908 21304 17233 21332
rect 16908 21292 16914 21304
rect 17221 21301 17233 21304
rect 17267 21301 17279 21335
rect 17221 21295 17279 21301
rect 23017 21335 23075 21341
rect 23017 21301 23029 21335
rect 23063 21332 23075 21335
rect 23658 21332 23664 21344
rect 23063 21304 23664 21332
rect 23063 21301 23075 21304
rect 23017 21295 23075 21301
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 28994 21292 29000 21344
rect 29052 21332 29058 21344
rect 30653 21335 30711 21341
rect 30653 21332 30665 21335
rect 29052 21304 30665 21332
rect 29052 21292 29058 21304
rect 30653 21301 30665 21304
rect 30699 21301 30711 21335
rect 30653 21295 30711 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 2038 21088 2044 21140
rect 2096 21128 2102 21140
rect 2133 21131 2191 21137
rect 2133 21128 2145 21131
rect 2096 21100 2145 21128
rect 2096 21088 2102 21100
rect 2133 21097 2145 21100
rect 2179 21128 2191 21131
rect 2222 21128 2228 21140
rect 2179 21100 2228 21128
rect 2179 21097 2191 21100
rect 2133 21091 2191 21097
rect 2222 21088 2228 21100
rect 2280 21088 2286 21140
rect 5169 21131 5227 21137
rect 5169 21097 5181 21131
rect 5215 21128 5227 21131
rect 5350 21128 5356 21140
rect 5215 21100 5356 21128
rect 5215 21097 5227 21100
rect 5169 21091 5227 21097
rect 5350 21088 5356 21100
rect 5408 21088 5414 21140
rect 7929 21131 7987 21137
rect 7929 21097 7941 21131
rect 7975 21128 7987 21131
rect 13725 21131 13783 21137
rect 7975 21100 12480 21128
rect 7975 21097 7987 21100
rect 7929 21091 7987 21097
rect 1394 21020 1400 21072
rect 1452 21060 1458 21072
rect 4154 21060 4160 21072
rect 1452 21032 4160 21060
rect 1452 21020 1458 21032
rect 4154 21020 4160 21032
rect 4212 21020 4218 21072
rect 4706 21020 4712 21072
rect 4764 21060 4770 21072
rect 4890 21060 4896 21072
rect 4764 21032 4896 21060
rect 4764 21020 4770 21032
rect 4890 21020 4896 21032
rect 4948 21020 4954 21072
rect 4525 20995 4583 21001
rect 4525 20961 4537 20995
rect 4571 20992 4583 20995
rect 11606 20992 11612 21004
rect 4571 20964 11612 20992
rect 4571 20961 4583 20964
rect 4525 20955 4583 20961
rect 11606 20952 11612 20964
rect 11664 20952 11670 21004
rect 11885 20995 11943 21001
rect 11885 20961 11897 20995
rect 11931 20992 11943 20995
rect 12158 20992 12164 21004
rect 11931 20964 12164 20992
rect 11931 20961 11943 20964
rect 11885 20955 11943 20961
rect 12158 20952 12164 20964
rect 12216 20952 12222 21004
rect 12452 20992 12480 21100
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 17126 21128 17132 21140
rect 13771 21100 17132 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 17126 21088 17132 21100
rect 17184 21088 17190 21140
rect 13906 21020 13912 21072
rect 13964 21060 13970 21072
rect 16574 21060 16580 21072
rect 13964 21032 16580 21060
rect 13964 21020 13970 21032
rect 16574 21020 16580 21032
rect 16632 21020 16638 21072
rect 18509 21063 18567 21069
rect 18509 21029 18521 21063
rect 18555 21060 18567 21063
rect 19058 21060 19064 21072
rect 18555 21032 19064 21060
rect 18555 21029 18567 21032
rect 18509 21023 18567 21029
rect 19058 21020 19064 21032
rect 19116 21060 19122 21072
rect 20070 21060 20076 21072
rect 19116 21032 19564 21060
rect 20031 21032 20076 21060
rect 19116 21020 19122 21032
rect 14461 20995 14519 21001
rect 14461 20992 14473 20995
rect 12452 20964 14473 20992
rect 14461 20961 14473 20964
rect 14507 20961 14519 20995
rect 14461 20955 14519 20961
rect 15654 20952 15660 21004
rect 15712 20992 15718 21004
rect 16025 20995 16083 21001
rect 16025 20992 16037 20995
rect 15712 20964 16037 20992
rect 15712 20952 15718 20964
rect 16025 20961 16037 20964
rect 16071 20992 16083 20995
rect 16482 20992 16488 21004
rect 16071 20964 16488 20992
rect 16071 20961 16083 20964
rect 16025 20955 16083 20961
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 16850 20992 16856 21004
rect 16811 20964 16856 20992
rect 16850 20952 16856 20964
rect 16908 20952 16914 21004
rect 18693 20995 18751 21001
rect 18693 20961 18705 20995
rect 18739 20992 18751 20995
rect 19334 20992 19340 21004
rect 18739 20964 19340 20992
rect 18739 20961 18751 20964
rect 18693 20955 18751 20961
rect 19334 20952 19340 20964
rect 19392 20952 19398 21004
rect 19536 21001 19564 21032
rect 20070 21020 20076 21032
rect 20128 21020 20134 21072
rect 21266 21020 21272 21072
rect 21324 21060 21330 21072
rect 21361 21063 21419 21069
rect 21361 21060 21373 21063
rect 21324 21032 21373 21060
rect 21324 21020 21330 21032
rect 21361 21029 21373 21032
rect 21407 21029 21419 21063
rect 21361 21023 21419 21029
rect 23382 21020 23388 21072
rect 23440 21020 23446 21072
rect 19521 20995 19579 21001
rect 19521 20961 19533 20995
rect 19567 20961 19579 20995
rect 21910 20992 21916 21004
rect 21871 20964 21916 20992
rect 19521 20955 19579 20961
rect 21910 20952 21916 20964
rect 21968 20952 21974 21004
rect 22462 20952 22468 21004
rect 22520 20992 22526 21004
rect 23109 20995 23167 21001
rect 23109 20992 23121 20995
rect 22520 20964 23121 20992
rect 22520 20952 22526 20964
rect 23109 20961 23121 20964
rect 23155 20992 23167 20995
rect 23400 20992 23428 21020
rect 23155 20964 23428 20992
rect 23155 20961 23167 20964
rect 23109 20955 23167 20961
rect 4433 20927 4491 20933
rect 4433 20893 4445 20927
rect 4479 20924 4491 20927
rect 4890 20924 4896 20936
rect 4479 20896 4896 20924
rect 4479 20893 4491 20896
rect 4433 20887 4491 20893
rect 4890 20884 4896 20896
rect 4948 20884 4954 20936
rect 5166 20884 5172 20936
rect 5224 20924 5230 20936
rect 5350 20924 5356 20936
rect 5224 20896 5356 20924
rect 5224 20884 5230 20896
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 6917 20927 6975 20933
rect 6917 20893 6929 20927
rect 6963 20924 6975 20927
rect 7466 20924 7472 20936
rect 6963 20896 7472 20924
rect 6963 20893 6975 20896
rect 6917 20887 6975 20893
rect 7466 20884 7472 20896
rect 7524 20884 7530 20936
rect 7745 20927 7803 20933
rect 7745 20893 7757 20927
rect 7791 20924 7803 20927
rect 8573 20927 8631 20933
rect 7791 20896 8432 20924
rect 7791 20893 7803 20896
rect 7745 20887 7803 20893
rect 3421 20859 3479 20865
rect 3421 20825 3433 20859
rect 3467 20825 3479 20859
rect 3421 20819 3479 20825
rect 3436 20788 3464 20819
rect 5902 20816 5908 20868
rect 5960 20816 5966 20868
rect 6641 20859 6699 20865
rect 6641 20825 6653 20859
rect 6687 20856 6699 20859
rect 8202 20856 8208 20868
rect 6687 20828 8208 20856
rect 6687 20825 6699 20828
rect 6641 20819 6699 20825
rect 8202 20816 8208 20828
rect 8260 20816 8266 20868
rect 6822 20788 6828 20800
rect 3436 20760 6828 20788
rect 6822 20748 6828 20760
rect 6880 20748 6886 20800
rect 7282 20748 7288 20800
rect 7340 20788 7346 20800
rect 7742 20788 7748 20800
rect 7340 20760 7748 20788
rect 7340 20748 7346 20760
rect 7742 20748 7748 20760
rect 7800 20748 7806 20800
rect 8404 20797 8432 20896
rect 8573 20893 8585 20927
rect 8619 20924 8631 20927
rect 8846 20924 8852 20936
rect 8619 20896 8852 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 8846 20884 8852 20896
rect 8904 20884 8910 20936
rect 9122 20924 9128 20936
rect 9083 20896 9128 20924
rect 9122 20884 9128 20896
rect 9180 20884 9186 20936
rect 11054 20884 11060 20936
rect 11112 20924 11118 20936
rect 12069 20927 12127 20933
rect 12069 20924 12081 20927
rect 11112 20896 12081 20924
rect 11112 20884 11118 20896
rect 12069 20893 12081 20896
rect 12115 20893 12127 20927
rect 13538 20924 13544 20936
rect 13499 20896 13544 20924
rect 12069 20887 12127 20893
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 14274 20924 14280 20936
rect 14235 20896 14280 20924
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 14366 20884 14372 20936
rect 14424 20924 14430 20936
rect 15841 20927 15899 20933
rect 15841 20924 15853 20927
rect 14424 20896 15853 20924
rect 14424 20884 14430 20896
rect 15841 20893 15853 20896
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 20625 20927 20683 20933
rect 20625 20893 20637 20927
rect 20671 20924 20683 20927
rect 21174 20924 21180 20936
rect 20671 20896 21180 20924
rect 20671 20893 20683 20896
rect 20625 20887 20683 20893
rect 8478 20816 8484 20868
rect 8536 20856 8542 20868
rect 9401 20859 9459 20865
rect 9401 20856 9413 20859
rect 8536 20828 9413 20856
rect 8536 20816 8542 20828
rect 9401 20825 9413 20828
rect 9447 20825 9459 20859
rect 9401 20819 9459 20825
rect 9858 20816 9864 20868
rect 9916 20816 9922 20868
rect 13906 20856 13912 20868
rect 10888 20828 13912 20856
rect 8389 20791 8447 20797
rect 8389 20757 8401 20791
rect 8435 20757 8447 20791
rect 8389 20751 8447 20757
rect 8846 20748 8852 20800
rect 8904 20788 8910 20800
rect 9490 20788 9496 20800
rect 8904 20760 9496 20788
rect 8904 20748 8910 20760
rect 9490 20748 9496 20760
rect 9548 20748 9554 20800
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 10888 20797 10916 20828
rect 13906 20816 13912 20828
rect 13964 20816 13970 20868
rect 13998 20816 14004 20868
rect 14056 20856 14062 20868
rect 15102 20856 15108 20868
rect 14056 20828 15108 20856
rect 14056 20816 14062 20828
rect 15102 20816 15108 20828
rect 15160 20816 15166 20868
rect 15654 20816 15660 20868
rect 15712 20856 15718 20868
rect 16945 20859 17003 20865
rect 16945 20856 16957 20859
rect 15712 20828 16957 20856
rect 15712 20816 15718 20828
rect 16945 20825 16957 20828
rect 16991 20825 17003 20859
rect 16945 20819 17003 20825
rect 17497 20859 17555 20865
rect 17497 20825 17509 20859
rect 17543 20856 17555 20859
rect 18782 20856 18788 20868
rect 17543 20828 18788 20856
rect 17543 20825 17555 20828
rect 17497 20819 17555 20825
rect 10873 20791 10931 20797
rect 10873 20788 10885 20791
rect 9732 20760 10885 20788
rect 9732 20748 9738 20760
rect 10873 20757 10885 20760
rect 10919 20757 10931 20791
rect 10873 20751 10931 20757
rect 12342 20748 12348 20800
rect 12400 20788 12406 20800
rect 12529 20791 12587 20797
rect 12529 20788 12541 20791
rect 12400 20760 12541 20788
rect 12400 20748 12406 20760
rect 12529 20757 12541 20760
rect 12575 20757 12587 20791
rect 12529 20751 12587 20757
rect 14921 20791 14979 20797
rect 14921 20757 14933 20791
rect 14967 20788 14979 20791
rect 15010 20788 15016 20800
rect 14967 20760 15016 20788
rect 14967 20757 14979 20760
rect 14921 20751 14979 20757
rect 15010 20748 15016 20760
rect 15068 20748 15074 20800
rect 15381 20791 15439 20797
rect 15381 20757 15393 20791
rect 15427 20788 15439 20791
rect 15470 20788 15476 20800
rect 15427 20760 15476 20788
rect 15427 20757 15439 20760
rect 15381 20751 15439 20757
rect 15470 20748 15476 20760
rect 15528 20748 15534 20800
rect 15930 20748 15936 20800
rect 15988 20788 15994 20800
rect 17512 20788 17540 20819
rect 18782 20816 18788 20828
rect 18840 20816 18846 20868
rect 15988 20760 17540 20788
rect 18892 20788 18920 20887
rect 21174 20884 21180 20896
rect 21232 20884 21238 20936
rect 32214 20924 32220 20936
rect 32175 20896 32220 20924
rect 32214 20884 32220 20896
rect 32272 20884 32278 20936
rect 19613 20859 19671 20865
rect 19613 20825 19625 20859
rect 19659 20856 19671 20859
rect 19978 20856 19984 20868
rect 19659 20828 19984 20856
rect 19659 20825 19671 20828
rect 19613 20819 19671 20825
rect 19978 20816 19984 20828
rect 20036 20816 20042 20868
rect 21821 20859 21879 20865
rect 21821 20825 21833 20859
rect 21867 20825 21879 20859
rect 22830 20856 22836 20868
rect 22791 20828 22836 20856
rect 21821 20819 21879 20825
rect 20070 20788 20076 20800
rect 18892 20760 20076 20788
rect 15988 20748 15994 20760
rect 20070 20748 20076 20760
rect 20128 20748 20134 20800
rect 20809 20791 20867 20797
rect 20809 20757 20821 20791
rect 20855 20788 20867 20791
rect 21836 20788 21864 20819
rect 22830 20816 22836 20828
rect 22888 20816 22894 20868
rect 22925 20859 22983 20865
rect 22925 20825 22937 20859
rect 22971 20825 22983 20859
rect 22925 20819 22983 20825
rect 20855 20760 21864 20788
rect 22940 20788 22968 20819
rect 23566 20788 23572 20800
rect 22940 20760 23572 20788
rect 20855 20757 20867 20760
rect 20809 20751 20867 20757
rect 23566 20748 23572 20760
rect 23624 20748 23630 20800
rect 32122 20788 32128 20800
rect 32083 20760 32128 20788
rect 32122 20748 32128 20760
rect 32180 20748 32186 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1670 20584 1676 20596
rect 1631 20556 1676 20584
rect 1670 20544 1676 20556
rect 1728 20544 1734 20596
rect 3970 20544 3976 20596
rect 4028 20584 4034 20596
rect 6914 20584 6920 20596
rect 4028 20556 6920 20584
rect 4028 20544 4034 20556
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 7009 20587 7067 20593
rect 7009 20553 7021 20587
rect 7055 20584 7067 20587
rect 10226 20584 10232 20596
rect 7055 20556 9996 20584
rect 10187 20556 10232 20584
rect 7055 20553 7067 20556
rect 7009 20547 7067 20553
rect 3142 20476 3148 20528
rect 3200 20476 3206 20528
rect 4154 20516 4160 20528
rect 4067 20488 4160 20516
rect 4154 20476 4160 20488
rect 4212 20516 4218 20528
rect 4212 20488 4752 20516
rect 4212 20476 4218 20488
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20448 1915 20451
rect 2866 20448 2872 20460
rect 1903 20420 2872 20448
rect 1903 20417 1915 20420
rect 1857 20411 1915 20417
rect 2866 20408 2872 20420
rect 2924 20408 2930 20460
rect 2409 20383 2467 20389
rect 2409 20349 2421 20383
rect 2455 20380 2467 20383
rect 3418 20380 3424 20392
rect 2455 20352 3424 20380
rect 2455 20349 2467 20352
rect 2409 20343 2467 20349
rect 3418 20340 3424 20352
rect 3476 20340 3482 20392
rect 4433 20383 4491 20389
rect 4433 20349 4445 20383
rect 4479 20380 4491 20383
rect 4614 20380 4620 20392
rect 4479 20352 4620 20380
rect 4479 20349 4491 20352
rect 4433 20343 4491 20349
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 4724 20380 4752 20488
rect 5534 20476 5540 20528
rect 5592 20516 5598 20528
rect 7834 20516 7840 20528
rect 5592 20488 7840 20516
rect 5592 20476 5598 20488
rect 7834 20476 7840 20488
rect 7892 20476 7898 20528
rect 8754 20476 8760 20528
rect 8812 20476 8818 20528
rect 5166 20448 5172 20460
rect 5127 20420 5172 20448
rect 5166 20408 5172 20420
rect 5224 20408 5230 20460
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20448 5871 20451
rect 6270 20448 6276 20460
rect 5859 20420 6276 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 6270 20408 6276 20420
rect 6328 20408 6334 20460
rect 6825 20451 6883 20457
rect 6825 20417 6837 20451
rect 6871 20448 6883 20451
rect 7098 20448 7104 20460
rect 6871 20420 7104 20448
rect 6871 20417 6883 20420
rect 6825 20411 6883 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 9030 20408 9036 20460
rect 9088 20448 9094 20460
rect 9858 20448 9864 20460
rect 9088 20420 9864 20448
rect 9088 20408 9094 20420
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 9968 20448 9996 20556
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 12342 20584 12348 20596
rect 12303 20556 12348 20584
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 14093 20587 14151 20593
rect 14093 20553 14105 20587
rect 14139 20584 14151 20587
rect 14182 20584 14188 20596
rect 14139 20556 14188 20584
rect 14139 20553 14151 20556
rect 14093 20547 14151 20553
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 14826 20584 14832 20596
rect 14787 20556 14832 20584
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 15933 20587 15991 20593
rect 15933 20553 15945 20587
rect 15979 20584 15991 20587
rect 16022 20584 16028 20596
rect 15979 20556 16028 20584
rect 15979 20553 15991 20556
rect 15933 20547 15991 20553
rect 16022 20544 16028 20556
rect 16080 20544 16086 20596
rect 18417 20587 18475 20593
rect 18417 20553 18429 20587
rect 18463 20584 18475 20587
rect 18506 20584 18512 20596
rect 18463 20556 18512 20584
rect 18463 20553 18475 20556
rect 18417 20547 18475 20553
rect 18506 20544 18512 20556
rect 18564 20544 18570 20596
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19521 20587 19579 20593
rect 19521 20584 19533 20587
rect 19392 20556 19533 20584
rect 19392 20544 19398 20556
rect 19521 20553 19533 20556
rect 19567 20553 19579 20587
rect 19521 20547 19579 20553
rect 20070 20544 20076 20596
rect 20128 20584 20134 20596
rect 20165 20587 20223 20593
rect 20165 20584 20177 20587
rect 20128 20556 20177 20584
rect 20128 20544 20134 20556
rect 20165 20553 20177 20556
rect 20211 20553 20223 20587
rect 20165 20547 20223 20553
rect 21174 20544 21180 20596
rect 21232 20584 21238 20596
rect 21269 20587 21327 20593
rect 21269 20584 21281 20587
rect 21232 20556 21281 20584
rect 21232 20544 21238 20556
rect 21269 20553 21281 20556
rect 21315 20553 21327 20587
rect 22830 20584 22836 20596
rect 22791 20556 22836 20584
rect 21269 20547 21327 20553
rect 22830 20544 22836 20556
rect 22888 20544 22894 20596
rect 23477 20587 23535 20593
rect 23477 20553 23489 20587
rect 23523 20584 23535 20587
rect 23566 20584 23572 20596
rect 23523 20556 23572 20584
rect 23523 20553 23535 20556
rect 23477 20547 23535 20553
rect 23566 20544 23572 20556
rect 23624 20544 23630 20596
rect 10873 20519 10931 20525
rect 10873 20485 10885 20519
rect 10919 20516 10931 20519
rect 14274 20516 14280 20528
rect 10919 20488 14280 20516
rect 10919 20485 10931 20488
rect 10873 20479 10931 20485
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 10045 20451 10103 20457
rect 10045 20448 10057 20451
rect 9968 20420 10057 20448
rect 10045 20417 10057 20420
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 11606 20408 11612 20460
rect 11664 20448 11670 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11664 20420 11897 20448
rect 11664 20408 11670 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 13357 20451 13415 20457
rect 13357 20448 13369 20451
rect 12768 20420 13369 20448
rect 12768 20408 12774 20420
rect 13357 20417 13369 20420
rect 13403 20417 13415 20451
rect 13998 20448 14004 20460
rect 13959 20420 14004 20448
rect 13357 20411 13415 20417
rect 13998 20408 14004 20420
rect 14056 20408 14062 20460
rect 14645 20451 14703 20457
rect 14645 20417 14657 20451
rect 14691 20417 14703 20451
rect 14645 20411 14703 20417
rect 6362 20380 6368 20392
rect 4724 20352 6368 20380
rect 6362 20340 6368 20352
rect 6420 20340 6426 20392
rect 7466 20380 7472 20392
rect 7427 20352 7472 20380
rect 7466 20340 7472 20352
rect 7524 20340 7530 20392
rect 7745 20383 7803 20389
rect 7745 20380 7757 20383
rect 7576 20352 7757 20380
rect 7282 20312 7288 20324
rect 4356 20284 7288 20312
rect 3418 20204 3424 20256
rect 3476 20244 3482 20256
rect 4356 20244 4384 20284
rect 7282 20272 7288 20284
rect 7340 20312 7346 20324
rect 7576 20312 7604 20352
rect 7745 20349 7757 20352
rect 7791 20349 7803 20383
rect 7745 20343 7803 20349
rect 7834 20340 7840 20392
rect 7892 20380 7898 20392
rect 9490 20380 9496 20392
rect 7892 20352 8800 20380
rect 9451 20352 9496 20380
rect 7892 20340 7898 20352
rect 7340 20284 7604 20312
rect 8772 20312 8800 20352
rect 9490 20340 9496 20352
rect 9548 20340 9554 20392
rect 11054 20380 11060 20392
rect 9600 20352 11060 20380
rect 9600 20312 9628 20352
rect 11054 20340 11060 20352
rect 11112 20340 11118 20392
rect 11330 20340 11336 20392
rect 11388 20380 11394 20392
rect 11701 20383 11759 20389
rect 11701 20380 11713 20383
rect 11388 20352 11713 20380
rect 11388 20340 11394 20352
rect 11701 20349 11713 20352
rect 11747 20349 11759 20383
rect 11701 20343 11759 20349
rect 8772 20284 9628 20312
rect 14660 20312 14688 20411
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 15289 20451 15347 20457
rect 15289 20448 15301 20451
rect 14976 20420 15301 20448
rect 14976 20408 14982 20420
rect 15289 20417 15301 20420
rect 15335 20417 15347 20451
rect 15289 20411 15347 20417
rect 15378 20408 15384 20460
rect 15436 20448 15442 20460
rect 15473 20451 15531 20457
rect 15473 20448 15485 20451
rect 15436 20420 15485 20448
rect 15436 20408 15442 20420
rect 15473 20417 15485 20420
rect 15519 20417 15531 20451
rect 17310 20448 17316 20460
rect 17271 20420 17316 20448
rect 15473 20411 15531 20417
rect 17310 20408 17316 20420
rect 17368 20408 17374 20460
rect 17678 20408 17684 20460
rect 17736 20448 17742 20460
rect 17957 20451 18015 20457
rect 17957 20448 17969 20451
rect 17736 20420 17969 20448
rect 17736 20408 17742 20420
rect 17957 20417 17969 20420
rect 18003 20417 18015 20451
rect 17957 20411 18015 20417
rect 18138 20408 18144 20460
rect 18196 20448 18202 20460
rect 18690 20448 18696 20460
rect 18196 20420 18696 20448
rect 18196 20408 18202 20420
rect 18690 20408 18696 20420
rect 18748 20448 18754 20460
rect 18877 20451 18935 20457
rect 18877 20448 18889 20451
rect 18748 20420 18889 20448
rect 18748 20408 18754 20420
rect 18877 20417 18889 20420
rect 18923 20417 18935 20451
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 18877 20411 18935 20417
rect 19076 20420 19717 20448
rect 17773 20383 17831 20389
rect 17773 20349 17785 20383
rect 17819 20380 17831 20383
rect 18046 20380 18052 20392
rect 17819 20352 18052 20380
rect 17819 20349 17831 20352
rect 17773 20343 17831 20349
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 19076 20321 19104 20420
rect 19705 20417 19717 20420
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 21358 20408 21364 20460
rect 21416 20448 21422 20460
rect 21453 20451 21511 20457
rect 21453 20448 21465 20451
rect 21416 20420 21465 20448
rect 21416 20408 21422 20420
rect 21453 20417 21465 20420
rect 21499 20417 21511 20451
rect 22002 20448 22008 20460
rect 21963 20420 22008 20448
rect 21453 20411 21511 20417
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 23658 20448 23664 20460
rect 23619 20420 23664 20448
rect 23658 20408 23664 20420
rect 23716 20408 23722 20460
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20417 24179 20451
rect 24121 20411 24179 20417
rect 21082 20340 21088 20392
rect 21140 20380 21146 20392
rect 24136 20380 24164 20411
rect 24578 20380 24584 20392
rect 21140 20352 24584 20380
rect 21140 20340 21146 20352
rect 24578 20340 24584 20352
rect 24636 20340 24642 20392
rect 17129 20315 17187 20321
rect 17129 20312 17141 20315
rect 14660 20284 17141 20312
rect 7340 20272 7346 20284
rect 17129 20281 17141 20284
rect 17175 20281 17187 20315
rect 17129 20275 17187 20281
rect 19061 20315 19119 20321
rect 19061 20281 19073 20315
rect 19107 20281 19119 20315
rect 19061 20275 19119 20281
rect 3476 20216 4384 20244
rect 5353 20247 5411 20253
rect 3476 20204 3482 20216
rect 5353 20213 5365 20247
rect 5399 20244 5411 20247
rect 5534 20244 5540 20256
rect 5399 20216 5540 20244
rect 5399 20213 5411 20216
rect 5353 20207 5411 20213
rect 5534 20204 5540 20216
rect 5592 20204 5598 20256
rect 5905 20247 5963 20253
rect 5905 20213 5917 20247
rect 5951 20244 5963 20247
rect 7374 20244 7380 20256
rect 5951 20216 7380 20244
rect 5951 20213 5963 20216
rect 5905 20207 5963 20213
rect 7374 20204 7380 20216
rect 7432 20204 7438 20256
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 9122 20244 9128 20256
rect 7524 20216 9128 20244
rect 7524 20204 7530 20216
rect 9122 20204 9128 20216
rect 9180 20204 9186 20256
rect 9582 20204 9588 20256
rect 9640 20244 9646 20256
rect 13262 20244 13268 20256
rect 9640 20216 13268 20244
rect 9640 20204 9646 20216
rect 13262 20204 13268 20216
rect 13320 20204 13326 20256
rect 13538 20244 13544 20256
rect 13499 20216 13544 20244
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 15470 20244 15476 20256
rect 13780 20216 15476 20244
rect 13780 20204 13786 20216
rect 15470 20204 15476 20216
rect 15528 20204 15534 20256
rect 22097 20247 22155 20253
rect 22097 20213 22109 20247
rect 22143 20244 22155 20247
rect 22278 20244 22284 20256
rect 22143 20216 22284 20244
rect 22143 20213 22155 20216
rect 22097 20207 22155 20213
rect 22278 20204 22284 20216
rect 22336 20204 22342 20256
rect 24305 20247 24363 20253
rect 24305 20213 24317 20247
rect 24351 20244 24363 20247
rect 25498 20244 25504 20256
rect 24351 20216 25504 20244
rect 24351 20213 24363 20216
rect 24305 20207 24363 20213
rect 25498 20204 25504 20216
rect 25556 20204 25562 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 3418 20040 3424 20052
rect 3379 20012 3424 20040
rect 3418 20000 3424 20012
rect 3476 20000 3482 20052
rect 4433 20043 4491 20049
rect 4433 20009 4445 20043
rect 4479 20040 4491 20043
rect 5166 20040 5172 20052
rect 4479 20012 5172 20040
rect 4479 20009 4491 20012
rect 4433 20003 4491 20009
rect 5166 20000 5172 20012
rect 5224 20000 5230 20052
rect 6178 20040 6184 20052
rect 5644 20012 6184 20040
rect 4890 19972 4896 19984
rect 4264 19944 4896 19972
rect 1673 19907 1731 19913
rect 1673 19873 1685 19907
rect 1719 19904 1731 19907
rect 2038 19904 2044 19916
rect 1719 19876 2044 19904
rect 1719 19873 1731 19876
rect 1673 19867 1731 19873
rect 2038 19864 2044 19876
rect 2096 19864 2102 19916
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 4264 19845 4292 19944
rect 4890 19932 4896 19944
rect 4948 19932 4954 19984
rect 5077 19975 5135 19981
rect 5077 19941 5089 19975
rect 5123 19972 5135 19975
rect 5644 19972 5672 20012
rect 6178 20000 6184 20012
rect 6236 20000 6242 20052
rect 6270 20000 6276 20052
rect 6328 20040 6334 20052
rect 6914 20040 6920 20052
rect 6328 20012 6920 20040
rect 6328 20000 6334 20012
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 9030 20040 9036 20052
rect 7024 20012 9036 20040
rect 7024 19972 7052 20012
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 9214 20040 9220 20052
rect 9171 20012 9220 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 9214 20000 9220 20012
rect 9272 20000 9278 20052
rect 12066 20040 12072 20052
rect 9600 20012 12072 20040
rect 5123 19944 5672 19972
rect 6840 19944 7052 19972
rect 5123 19941 5135 19944
rect 5077 19935 5135 19941
rect 6270 19904 6276 19916
rect 4908 19876 6276 19904
rect 4908 19845 4936 19876
rect 6270 19864 6276 19876
rect 6328 19864 6334 19916
rect 6362 19864 6368 19916
rect 6420 19904 6426 19916
rect 6840 19904 6868 19944
rect 7374 19932 7380 19984
rect 7432 19972 7438 19984
rect 9600 19972 9628 20012
rect 12066 20000 12072 20012
rect 12124 20000 12130 20052
rect 15197 20043 15255 20049
rect 15197 20009 15209 20043
rect 15243 20040 15255 20043
rect 16022 20040 16028 20052
rect 15243 20012 16028 20040
rect 15243 20009 15255 20012
rect 15197 20003 15255 20009
rect 16022 20000 16028 20012
rect 16080 20000 16086 20052
rect 16942 20000 16948 20052
rect 17000 20040 17006 20052
rect 18049 20043 18107 20049
rect 18049 20040 18061 20043
rect 17000 20012 18061 20040
rect 17000 20000 17006 20012
rect 18049 20009 18061 20012
rect 18095 20040 18107 20043
rect 18230 20040 18236 20052
rect 18095 20012 18236 20040
rect 18095 20009 18107 20012
rect 18049 20003 18107 20009
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 29178 20040 29184 20052
rect 19306 20012 29184 20040
rect 7432 19944 9628 19972
rect 13725 19975 13783 19981
rect 7432 19932 7438 19944
rect 13725 19941 13737 19975
rect 13771 19972 13783 19975
rect 14366 19972 14372 19984
rect 13771 19944 14372 19972
rect 13771 19941 13783 19944
rect 13725 19935 13783 19941
rect 14366 19932 14372 19944
rect 14424 19932 14430 19984
rect 16482 19932 16488 19984
rect 16540 19972 16546 19984
rect 16540 19944 17448 19972
rect 16540 19932 16546 19944
rect 7006 19904 7012 19916
rect 6420 19876 6868 19904
rect 6932 19876 7012 19904
rect 6420 19864 6426 19876
rect 4249 19839 4307 19845
rect 4249 19836 4261 19839
rect 4212 19808 4261 19836
rect 4212 19796 4218 19808
rect 4249 19805 4261 19808
rect 4295 19805 4307 19839
rect 4249 19799 4307 19805
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19805 4951 19839
rect 4893 19799 4951 19805
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19805 5595 19839
rect 6932 19822 6960 19876
rect 7006 19864 7012 19876
rect 7064 19864 7070 19916
rect 8846 19904 8852 19916
rect 7576 19876 8852 19904
rect 7576 19845 7604 19876
rect 8846 19864 8852 19876
rect 8904 19904 8910 19916
rect 9030 19904 9036 19916
rect 8904 19876 9036 19904
rect 8904 19864 8910 19876
rect 9030 19864 9036 19876
rect 9088 19864 9094 19916
rect 9122 19864 9128 19916
rect 9180 19904 9186 19916
rect 10873 19907 10931 19913
rect 10873 19904 10885 19907
rect 9180 19876 10885 19904
rect 9180 19864 9186 19876
rect 10873 19873 10885 19876
rect 10919 19873 10931 19907
rect 10873 19867 10931 19873
rect 11790 19864 11796 19916
rect 11848 19904 11854 19916
rect 11885 19907 11943 19913
rect 11885 19904 11897 19907
rect 11848 19876 11897 19904
rect 11848 19864 11854 19876
rect 11885 19873 11897 19876
rect 11931 19873 11943 19907
rect 11885 19867 11943 19873
rect 12529 19907 12587 19913
rect 12529 19873 12541 19907
rect 12575 19904 12587 19907
rect 12986 19904 12992 19916
rect 12575 19876 12992 19904
rect 12575 19873 12587 19876
rect 12529 19867 12587 19873
rect 12986 19864 12992 19876
rect 13044 19904 13050 19916
rect 16945 19907 17003 19913
rect 16945 19904 16957 19907
rect 13044 19876 16957 19904
rect 13044 19864 13050 19876
rect 16945 19873 16957 19876
rect 16991 19873 17003 19907
rect 17420 19904 17448 19944
rect 18693 19907 18751 19913
rect 18693 19904 18705 19907
rect 17420 19876 18705 19904
rect 16945 19867 17003 19873
rect 18693 19873 18705 19876
rect 18739 19904 18751 19907
rect 19306 19904 19334 20012
rect 29178 20000 29184 20012
rect 29236 20000 29242 20052
rect 20162 19932 20168 19984
rect 20220 19972 20226 19984
rect 21637 19975 21695 19981
rect 20220 19944 21496 19972
rect 20220 19932 20226 19944
rect 21358 19904 21364 19916
rect 18739 19876 19334 19904
rect 19536 19876 21364 19904
rect 18739 19873 18751 19876
rect 18693 19867 18751 19873
rect 7561 19839 7619 19845
rect 5537 19799 5595 19805
rect 7561 19805 7573 19839
rect 7607 19805 7619 19839
rect 7561 19799 7619 19805
rect 1949 19771 2007 19777
rect 1949 19737 1961 19771
rect 1995 19737 2007 19771
rect 1949 19731 2007 19737
rect 1964 19700 1992 19731
rect 2682 19728 2688 19780
rect 2740 19728 2746 19780
rect 4614 19728 4620 19780
rect 4672 19768 4678 19780
rect 5552 19768 5580 19799
rect 8202 19796 8208 19848
rect 8260 19836 8266 19848
rect 8389 19839 8447 19845
rect 8389 19836 8401 19839
rect 8260 19808 8401 19836
rect 8260 19796 8266 19808
rect 8389 19805 8401 19808
rect 8435 19805 8447 19839
rect 8389 19799 8447 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19805 12127 19839
rect 12069 19799 12127 19805
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 14274 19836 14280 19848
rect 13587 19808 14280 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 4672 19740 5580 19768
rect 4672 19728 4678 19740
rect 5718 19728 5724 19780
rect 5776 19768 5782 19780
rect 5813 19771 5871 19777
rect 5813 19768 5825 19771
rect 5776 19740 5825 19768
rect 5776 19728 5782 19740
rect 5813 19737 5825 19740
rect 5859 19737 5871 19771
rect 5813 19731 5871 19737
rect 8754 19728 8760 19780
rect 8812 19768 8818 19780
rect 8812 19740 9430 19768
rect 8812 19728 8818 19740
rect 10318 19728 10324 19780
rect 10376 19768 10382 19780
rect 10597 19771 10655 19777
rect 10597 19768 10609 19771
rect 10376 19740 10609 19768
rect 10376 19728 10382 19740
rect 10597 19737 10609 19740
rect 10643 19737 10655 19771
rect 10597 19731 10655 19737
rect 10870 19728 10876 19780
rect 10928 19768 10934 19780
rect 12084 19768 12112 19799
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 14550 19836 14556 19848
rect 14511 19808 14556 19836
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 14737 19839 14795 19845
rect 14737 19805 14749 19839
rect 14783 19805 14795 19839
rect 14737 19799 14795 19805
rect 14752 19768 14780 19799
rect 17678 19796 17684 19848
rect 17736 19836 17742 19848
rect 19536 19845 19564 19876
rect 21358 19864 21364 19876
rect 21416 19864 21422 19916
rect 18509 19839 18567 19845
rect 18509 19836 18521 19839
rect 17736 19808 18521 19836
rect 17736 19796 17742 19808
rect 18509 19805 18521 19808
rect 18555 19805 18567 19839
rect 18509 19799 18567 19805
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 20162 19796 20168 19848
rect 20220 19836 20226 19848
rect 20349 19839 20407 19845
rect 20349 19836 20361 19839
rect 20220 19808 20361 19836
rect 20220 19796 20226 19808
rect 20349 19805 20361 19808
rect 20395 19805 20407 19839
rect 20990 19836 20996 19848
rect 20951 19808 20996 19836
rect 20349 19799 20407 19805
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 21468 19845 21496 19944
rect 21637 19941 21649 19975
rect 21683 19972 21695 19975
rect 29730 19972 29736 19984
rect 21683 19944 22094 19972
rect 21683 19941 21695 19944
rect 21637 19935 21695 19941
rect 21453 19839 21511 19845
rect 21453 19805 21465 19839
rect 21499 19805 21511 19839
rect 22066 19836 22094 19944
rect 22940 19944 29736 19972
rect 22281 19839 22339 19845
rect 22281 19836 22293 19839
rect 22066 19808 22293 19836
rect 21453 19799 21511 19805
rect 22281 19805 22293 19808
rect 22327 19805 22339 19839
rect 22281 19799 22339 19805
rect 15746 19768 15752 19780
rect 10928 19740 12112 19768
rect 12544 19740 14780 19768
rect 15707 19740 15752 19768
rect 10928 19728 10934 19740
rect 3418 19700 3424 19712
rect 1964 19672 3424 19700
rect 3418 19660 3424 19672
rect 3476 19700 3482 19712
rect 3970 19700 3976 19712
rect 3476 19672 3976 19700
rect 3476 19660 3482 19672
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 4798 19660 4804 19712
rect 4856 19700 4862 19712
rect 5902 19700 5908 19712
rect 4856 19672 5908 19700
rect 4856 19660 4862 19672
rect 5902 19660 5908 19672
rect 5960 19660 5966 19712
rect 7098 19660 7104 19712
rect 7156 19700 7162 19712
rect 8386 19700 8392 19712
rect 7156 19672 8392 19700
rect 7156 19660 7162 19672
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 12544 19700 12572 19740
rect 15746 19728 15752 19740
rect 15804 19728 15810 19780
rect 15838 19728 15844 19780
rect 15896 19768 15902 19780
rect 16390 19768 16396 19780
rect 15896 19740 15941 19768
rect 16351 19740 16396 19768
rect 15896 19728 15902 19740
rect 16390 19728 16396 19740
rect 16448 19728 16454 19780
rect 17034 19768 17040 19780
rect 16995 19740 17040 19768
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 17218 19728 17224 19780
rect 17276 19768 17282 19780
rect 17589 19771 17647 19777
rect 17589 19768 17601 19771
rect 17276 19740 17601 19768
rect 17276 19728 17282 19740
rect 17589 19737 17601 19740
rect 17635 19768 17647 19771
rect 22940 19768 22968 19944
rect 29730 19932 29736 19944
rect 29788 19932 29794 19984
rect 24026 19904 24032 19916
rect 23987 19876 24032 19904
rect 24026 19864 24032 19876
rect 24084 19864 24090 19916
rect 24578 19836 24584 19848
rect 24539 19808 24584 19836
rect 24578 19796 24584 19808
rect 24636 19796 24642 19848
rect 25406 19836 25412 19848
rect 25367 19808 25412 19836
rect 25406 19796 25412 19808
rect 25464 19796 25470 19848
rect 38286 19836 38292 19848
rect 38247 19808 38292 19836
rect 38286 19796 38292 19808
rect 38344 19796 38350 19848
rect 17635 19740 22968 19768
rect 17635 19737 17647 19740
rect 17589 19731 17647 19737
rect 23106 19728 23112 19780
rect 23164 19768 23170 19780
rect 23385 19771 23443 19777
rect 23385 19768 23397 19771
rect 23164 19740 23397 19768
rect 23164 19728 23170 19740
rect 23385 19737 23397 19740
rect 23431 19737 23443 19771
rect 23385 19731 23443 19737
rect 23477 19771 23535 19777
rect 23477 19737 23489 19771
rect 23523 19768 23535 19771
rect 24673 19771 24731 19777
rect 24673 19768 24685 19771
rect 23523 19740 24685 19768
rect 23523 19737 23535 19740
rect 23477 19731 23535 19737
rect 24673 19737 24685 19740
rect 24719 19737 24731 19771
rect 24673 19731 24731 19737
rect 8527 19672 12572 19700
rect 19705 19703 19763 19709
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 20070 19700 20076 19712
rect 19751 19672 20076 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20254 19700 20260 19712
rect 20215 19672 20260 19700
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 20806 19700 20812 19712
rect 20767 19672 20812 19700
rect 20806 19660 20812 19672
rect 20864 19660 20870 19712
rect 22094 19660 22100 19712
rect 22152 19700 22158 19712
rect 25222 19700 25228 19712
rect 22152 19672 22197 19700
rect 25183 19672 25228 19700
rect 22152 19660 22158 19672
rect 25222 19660 25228 19672
rect 25280 19660 25286 19712
rect 35526 19660 35532 19712
rect 35584 19700 35590 19712
rect 38105 19703 38163 19709
rect 38105 19700 38117 19703
rect 35584 19672 38117 19700
rect 35584 19660 35590 19672
rect 38105 19669 38117 19672
rect 38151 19669 38163 19703
rect 38105 19663 38163 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1857 19499 1915 19505
rect 1857 19465 1869 19499
rect 1903 19496 1915 19499
rect 2222 19496 2228 19508
rect 1903 19468 2228 19496
rect 1903 19465 1915 19468
rect 1857 19459 1915 19465
rect 2222 19456 2228 19468
rect 2280 19456 2286 19508
rect 3053 19499 3111 19505
rect 3053 19465 3065 19499
rect 3099 19496 3111 19499
rect 8110 19496 8116 19508
rect 3099 19468 8116 19496
rect 3099 19465 3111 19468
rect 3053 19459 3111 19465
rect 8110 19456 8116 19468
rect 8168 19456 8174 19508
rect 8386 19456 8392 19508
rect 8444 19496 8450 19508
rect 8444 19468 9904 19496
rect 8444 19456 8450 19468
rect 3878 19428 3884 19440
rect 1688 19400 3884 19428
rect 1688 19369 1716 19400
rect 3878 19388 3884 19400
rect 3936 19388 3942 19440
rect 4062 19388 4068 19440
rect 4120 19428 4126 19440
rect 4120 19400 4186 19428
rect 4120 19388 4126 19400
rect 5902 19388 5908 19440
rect 5960 19428 5966 19440
rect 9125 19431 9183 19437
rect 5960 19400 7958 19428
rect 5960 19388 5966 19400
rect 9125 19397 9137 19431
rect 9171 19428 9183 19431
rect 9674 19428 9680 19440
rect 9171 19400 9680 19428
rect 9171 19397 9183 19400
rect 9125 19391 9183 19397
rect 9674 19388 9680 19400
rect 9732 19388 9738 19440
rect 9876 19428 9904 19468
rect 9950 19456 9956 19508
rect 10008 19496 10014 19508
rect 12529 19499 12587 19505
rect 10008 19468 10053 19496
rect 10008 19456 10014 19468
rect 12529 19465 12541 19499
rect 12575 19496 12587 19499
rect 13722 19496 13728 19508
rect 12575 19468 13728 19496
rect 12575 19465 12587 19468
rect 12529 19459 12587 19465
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 14274 19496 14280 19508
rect 14235 19468 14280 19496
rect 14274 19456 14280 19468
rect 14332 19456 14338 19508
rect 14366 19456 14372 19508
rect 14424 19496 14430 19508
rect 15838 19496 15844 19508
rect 14424 19468 15844 19496
rect 14424 19456 14430 19468
rect 15838 19456 15844 19468
rect 15896 19456 15902 19508
rect 18414 19496 18420 19508
rect 15948 19468 18420 19496
rect 9876 19400 12434 19428
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19329 1731 19363
rect 2314 19360 2320 19372
rect 2275 19332 2320 19360
rect 1673 19323 1731 19329
rect 2314 19320 2320 19332
rect 2372 19320 2378 19372
rect 3145 19363 3203 19369
rect 3145 19329 3157 19363
rect 3191 19360 3203 19363
rect 3326 19360 3332 19372
rect 3191 19332 3332 19360
rect 3191 19329 3203 19332
rect 3145 19323 3203 19329
rect 3326 19320 3332 19332
rect 3384 19320 3390 19372
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 3694 19360 3700 19372
rect 3651 19332 3700 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 3694 19320 3700 19332
rect 3752 19320 3758 19372
rect 6917 19363 6975 19369
rect 6917 19329 6929 19363
rect 6963 19360 6975 19363
rect 7282 19360 7288 19372
rect 6963 19332 7288 19360
rect 6963 19329 6975 19332
rect 6917 19323 6975 19329
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 9401 19363 9459 19369
rect 9401 19329 9413 19363
rect 9447 19360 9459 19363
rect 9447 19332 9536 19360
rect 9447 19329 9459 19332
rect 9401 19323 9459 19329
rect 3970 19252 3976 19304
rect 4028 19292 4034 19304
rect 5353 19295 5411 19301
rect 5353 19292 5365 19295
rect 4028 19264 5365 19292
rect 4028 19252 4034 19264
rect 5353 19261 5365 19264
rect 5399 19261 5411 19295
rect 5353 19255 5411 19261
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19292 5687 19295
rect 5718 19292 5724 19304
rect 5675 19264 5724 19292
rect 5675 19261 5687 19264
rect 5629 19255 5687 19261
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 9508 19292 9536 19332
rect 9582 19320 9588 19372
rect 9640 19360 9646 19372
rect 9640 19332 9812 19360
rect 9640 19320 9646 19332
rect 9674 19292 9680 19304
rect 6104 19264 9352 19292
rect 9508 19264 9680 19292
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 6104 19156 6132 19264
rect 9324 19224 9352 19264
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 9784 19292 9812 19332
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 10318 19360 10324 19372
rect 9916 19332 9961 19360
rect 10060 19332 10324 19360
rect 9916 19320 9922 19332
rect 10060 19292 10088 19332
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19360 10563 19363
rect 10962 19360 10968 19372
rect 10551 19332 10968 19360
rect 10551 19329 10563 19332
rect 10505 19323 10563 19329
rect 10962 19320 10968 19332
rect 11020 19320 11026 19372
rect 11882 19360 11888 19372
rect 11843 19332 11888 19360
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 12406 19360 12434 19400
rect 13538 19388 13544 19440
rect 13596 19428 13602 19440
rect 15948 19428 15976 19468
rect 18414 19456 18420 19468
rect 18472 19456 18478 19508
rect 19058 19496 19064 19508
rect 19019 19468 19064 19496
rect 19058 19456 19064 19468
rect 19116 19456 19122 19508
rect 19705 19499 19763 19505
rect 19705 19465 19717 19499
rect 19751 19496 19763 19499
rect 21174 19496 21180 19508
rect 19751 19468 21180 19496
rect 19751 19465 19763 19468
rect 19705 19459 19763 19465
rect 21174 19456 21180 19468
rect 21232 19456 21238 19508
rect 16114 19428 16120 19440
rect 13596 19400 14964 19428
rect 13596 19388 13602 19400
rect 14366 19360 14372 19372
rect 12406 19332 14372 19360
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 14516 19332 14561 19360
rect 14516 19320 14522 19332
rect 14642 19320 14648 19372
rect 14700 19360 14706 19372
rect 14936 19369 14964 19400
rect 15028 19400 15976 19428
rect 16075 19400 16120 19428
rect 14921 19363 14979 19369
rect 14700 19332 14872 19360
rect 14700 19320 14706 19332
rect 9784 19264 10088 19292
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19261 10747 19295
rect 12066 19292 12072 19304
rect 12027 19264 12072 19292
rect 10689 19255 10747 19261
rect 10594 19224 10600 19236
rect 9324 19196 10600 19224
rect 10594 19184 10600 19196
rect 10652 19184 10658 19236
rect 7098 19156 7104 19168
rect 2547 19128 6132 19156
rect 7059 19128 7104 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 7190 19116 7196 19168
rect 7248 19156 7254 19168
rect 7650 19156 7656 19168
rect 7248 19128 7656 19156
rect 7248 19116 7254 19128
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 9582 19116 9588 19168
rect 9640 19156 9646 19168
rect 10705 19156 10733 19255
rect 12066 19252 12072 19264
rect 12124 19252 12130 19304
rect 13262 19252 13268 19304
rect 13320 19292 13326 19304
rect 13449 19295 13507 19301
rect 13449 19292 13461 19295
rect 13320 19264 13461 19292
rect 13320 19252 13326 19264
rect 13449 19261 13461 19264
rect 13495 19261 13507 19295
rect 13630 19292 13636 19304
rect 13591 19264 13636 19292
rect 13449 19255 13507 19261
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 14844 19292 14872 19332
rect 14921 19329 14933 19363
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15028 19292 15056 19400
rect 16114 19388 16120 19400
rect 16172 19388 16178 19440
rect 16209 19431 16267 19437
rect 16209 19397 16221 19431
rect 16255 19428 16267 19431
rect 32122 19428 32128 19440
rect 16255 19400 17908 19428
rect 16255 19397 16267 19400
rect 16209 19391 16267 19397
rect 17310 19360 17316 19372
rect 17271 19332 17316 19360
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 15562 19292 15568 19304
rect 14844 19264 15056 19292
rect 15523 19264 15568 19292
rect 15562 19252 15568 19264
rect 15620 19252 15626 19304
rect 17770 19292 17776 19304
rect 17731 19264 17776 19292
rect 17770 19252 17776 19264
rect 17828 19252 17834 19304
rect 17880 19292 17908 19400
rect 17972 19400 32128 19428
rect 17972 19369 18000 19400
rect 17957 19363 18015 19369
rect 17957 19329 17969 19363
rect 18003 19329 18015 19363
rect 19426 19360 19432 19372
rect 17957 19323 18015 19329
rect 18064 19332 19432 19360
rect 18064 19292 18092 19332
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 20165 19363 20223 19369
rect 20165 19329 20177 19363
rect 20211 19360 20223 19363
rect 20254 19360 20260 19372
rect 20211 19332 20260 19360
rect 20211 19329 20223 19332
rect 20165 19323 20223 19329
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 20346 19320 20352 19372
rect 20404 19360 20410 19372
rect 20809 19363 20867 19369
rect 20404 19332 20449 19360
rect 20404 19320 20410 19332
rect 20809 19329 20821 19363
rect 20855 19360 20867 19363
rect 21174 19360 21180 19372
rect 20855 19332 21180 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 21468 19369 21496 19400
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19329 21511 19363
rect 22186 19360 22192 19372
rect 22147 19332 22192 19360
rect 21453 19323 21511 19329
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 23106 19360 23112 19372
rect 23067 19332 23112 19360
rect 23106 19320 23112 19332
rect 23164 19320 23170 19372
rect 23768 19369 23796 19400
rect 32122 19388 32128 19400
rect 32180 19388 32186 19440
rect 23753 19363 23811 19369
rect 23753 19329 23765 19363
rect 23799 19329 23811 19363
rect 23753 19323 23811 19329
rect 24857 19363 24915 19369
rect 24857 19329 24869 19363
rect 24903 19329 24915 19363
rect 25498 19360 25504 19372
rect 25459 19332 25504 19360
rect 24857 19323 24915 19329
rect 18414 19292 18420 19304
rect 17880 19264 18092 19292
rect 18375 19264 18420 19292
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 18601 19295 18659 19301
rect 18601 19261 18613 19295
rect 18647 19292 18659 19295
rect 18782 19292 18788 19304
rect 18647 19264 18788 19292
rect 18647 19261 18659 19264
rect 18601 19255 18659 19261
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 21269 19295 21327 19301
rect 21269 19261 21281 19295
rect 21315 19261 21327 19295
rect 21269 19255 21327 19261
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19261 23627 19295
rect 23569 19255 23627 19261
rect 24673 19295 24731 19301
rect 24673 19261 24685 19295
rect 24719 19292 24731 19295
rect 24762 19292 24768 19304
rect 24719 19264 24768 19292
rect 24719 19261 24731 19264
rect 24673 19255 24731 19261
rect 15105 19227 15163 19233
rect 15105 19193 15117 19227
rect 15151 19224 15163 19227
rect 15654 19224 15660 19236
rect 15151 19196 15660 19224
rect 15151 19193 15163 19196
rect 15105 19187 15163 19193
rect 15654 19184 15660 19196
rect 15712 19184 15718 19236
rect 21284 19224 21312 19255
rect 22094 19224 22100 19236
rect 21284 19196 22100 19224
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 23584 19224 23612 19255
rect 24762 19252 24768 19264
rect 24820 19252 24826 19304
rect 24872 19292 24900 19323
rect 25498 19320 25504 19332
rect 25556 19320 25562 19372
rect 25038 19292 25044 19304
rect 24872 19264 25044 19292
rect 25038 19252 25044 19264
rect 25096 19292 25102 19304
rect 25866 19292 25872 19304
rect 25096 19264 25872 19292
rect 25096 19252 25102 19264
rect 25866 19252 25872 19264
rect 25924 19252 25930 19304
rect 25222 19224 25228 19236
rect 23584 19196 25228 19224
rect 25222 19184 25228 19196
rect 25280 19184 25286 19236
rect 11054 19156 11060 19168
rect 9640 19128 10733 19156
rect 11015 19128 11060 19156
rect 9640 19116 9646 19128
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12989 19159 13047 19165
rect 12989 19156 13001 19159
rect 12492 19128 13001 19156
rect 12492 19116 12498 19128
rect 12989 19125 13001 19128
rect 13035 19125 13047 19159
rect 12989 19119 13047 19125
rect 21266 19116 21272 19168
rect 21324 19156 21330 19168
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21324 19128 22017 19156
rect 21324 19116 21330 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 22005 19119 22063 19125
rect 24489 19159 24547 19165
rect 24489 19125 24501 19159
rect 24535 19156 24547 19159
rect 24670 19156 24676 19168
rect 24535 19128 24676 19156
rect 24535 19125 24547 19128
rect 24489 19119 24547 19125
rect 24670 19116 24676 19128
rect 24728 19116 24734 19168
rect 24854 19116 24860 19168
rect 24912 19156 24918 19168
rect 25317 19159 25375 19165
rect 25317 19156 25329 19159
rect 24912 19128 25329 19156
rect 24912 19116 24918 19128
rect 25317 19125 25329 19128
rect 25363 19125 25375 19159
rect 25317 19119 25375 19125
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 5064 18955 5122 18961
rect 5064 18921 5076 18955
rect 5110 18952 5122 18955
rect 8573 18955 8631 18961
rect 5110 18924 8524 18952
rect 5110 18921 5122 18924
rect 5064 18915 5122 18921
rect 6086 18844 6092 18896
rect 6144 18884 6150 18896
rect 6362 18884 6368 18896
rect 6144 18856 6368 18884
rect 6144 18844 6150 18856
rect 6362 18844 6368 18856
rect 6420 18884 6426 18896
rect 6549 18887 6607 18893
rect 6549 18884 6561 18887
rect 6420 18856 6561 18884
rect 6420 18844 6426 18856
rect 6549 18853 6561 18856
rect 6595 18853 6607 18887
rect 6549 18847 6607 18853
rect 1946 18776 1952 18828
rect 2004 18776 2010 18828
rect 3421 18819 3479 18825
rect 3421 18785 3433 18819
rect 3467 18816 3479 18819
rect 4614 18816 4620 18828
rect 3467 18788 4620 18816
rect 3467 18785 3479 18788
rect 3421 18779 3479 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 4798 18816 4804 18828
rect 4711 18788 4804 18816
rect 4798 18776 4804 18788
rect 4856 18816 4862 18828
rect 5718 18816 5724 18828
rect 4856 18788 5724 18816
rect 4856 18776 4862 18788
rect 5718 18776 5724 18788
rect 5776 18776 5782 18828
rect 8110 18816 8116 18828
rect 8071 18788 8116 18816
rect 8110 18776 8116 18788
rect 8168 18776 8174 18828
rect 8496 18816 8524 18924
rect 8573 18921 8585 18955
rect 8619 18952 8631 18955
rect 12434 18952 12440 18964
rect 8619 18924 12440 18952
rect 8619 18921 8631 18924
rect 8573 18915 8631 18921
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 12986 18952 12992 18964
rect 12947 18924 12992 18952
rect 12986 18912 12992 18924
rect 13044 18912 13050 18964
rect 13078 18912 13084 18964
rect 13136 18952 13142 18964
rect 14645 18955 14703 18961
rect 14645 18952 14657 18955
rect 13136 18924 14657 18952
rect 13136 18912 13142 18924
rect 14645 18921 14657 18924
rect 14691 18921 14703 18955
rect 19426 18952 19432 18964
rect 19387 18924 19432 18952
rect 14645 18915 14703 18921
rect 19426 18912 19432 18924
rect 19484 18912 19490 18964
rect 20901 18955 20959 18961
rect 20901 18921 20913 18955
rect 20947 18952 20959 18955
rect 20990 18952 20996 18964
rect 20947 18924 20996 18952
rect 20947 18921 20959 18924
rect 20901 18915 20959 18921
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 21361 18955 21419 18961
rect 21361 18921 21373 18955
rect 21407 18952 21419 18955
rect 21450 18952 21456 18964
rect 21407 18924 21456 18952
rect 21407 18921 21419 18924
rect 21361 18915 21419 18921
rect 21450 18912 21456 18924
rect 21508 18912 21514 18964
rect 25406 18912 25412 18964
rect 25464 18952 25470 18964
rect 25777 18955 25835 18961
rect 25777 18952 25789 18955
rect 25464 18924 25789 18952
rect 25464 18912 25470 18924
rect 25777 18921 25789 18924
rect 25823 18921 25835 18955
rect 25777 18915 25835 18921
rect 25866 18912 25872 18964
rect 25924 18952 25930 18964
rect 31021 18955 31079 18961
rect 31021 18952 31033 18955
rect 25924 18924 31033 18952
rect 25924 18912 25930 18924
rect 31021 18921 31033 18924
rect 31067 18921 31079 18955
rect 31021 18915 31079 18921
rect 8662 18844 8668 18896
rect 8720 18884 8726 18896
rect 9125 18887 9183 18893
rect 9125 18884 9137 18887
rect 8720 18856 9137 18884
rect 8720 18844 8726 18856
rect 9125 18853 9137 18856
rect 9171 18853 9183 18887
rect 18233 18887 18291 18893
rect 18233 18884 18245 18887
rect 9125 18847 9183 18853
rect 11072 18856 18245 18884
rect 11072 18828 11100 18856
rect 18233 18853 18245 18856
rect 18279 18853 18291 18887
rect 18233 18847 18291 18853
rect 18322 18844 18328 18896
rect 18380 18884 18386 18896
rect 21542 18884 21548 18896
rect 18380 18856 21548 18884
rect 18380 18844 18386 18856
rect 21542 18844 21548 18856
rect 21600 18844 21606 18896
rect 24762 18844 24768 18896
rect 24820 18884 24826 18896
rect 26421 18887 26479 18893
rect 26421 18884 26433 18887
rect 24820 18856 26433 18884
rect 24820 18844 24826 18856
rect 26421 18853 26433 18856
rect 26467 18853 26479 18887
rect 26421 18847 26479 18853
rect 9214 18816 9220 18828
rect 8496 18788 9220 18816
rect 9214 18776 9220 18788
rect 9272 18776 9278 18828
rect 11054 18816 11060 18828
rect 9416 18788 11060 18816
rect 1964 18748 1992 18776
rect 4341 18751 4399 18757
rect 1964 18720 2070 18748
rect 4341 18717 4353 18751
rect 4387 18748 4399 18751
rect 4430 18748 4436 18760
rect 4387 18720 4436 18748
rect 4387 18717 4399 18720
rect 4341 18711 4399 18717
rect 4430 18708 4436 18720
rect 4488 18708 4494 18760
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 7101 18751 7159 18757
rect 7101 18748 7113 18751
rect 6972 18720 7113 18748
rect 6972 18708 6978 18720
rect 7101 18717 7113 18720
rect 7147 18748 7159 18751
rect 7834 18748 7840 18760
rect 7147 18720 7840 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18748 7987 18751
rect 9416 18748 9444 18788
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11146 18776 11152 18828
rect 11204 18816 11210 18828
rect 13173 18819 13231 18825
rect 11204 18788 13124 18816
rect 11204 18776 11210 18788
rect 7975 18720 9444 18748
rect 7975 18717 7987 18720
rect 7929 18711 7987 18717
rect 9490 18708 9496 18760
rect 9548 18708 9554 18760
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 11609 18751 11667 18757
rect 10928 18720 10973 18748
rect 10928 18708 10934 18720
rect 11609 18717 11621 18751
rect 11655 18717 11667 18751
rect 11790 18748 11796 18760
rect 11751 18720 11796 18748
rect 11609 18711 11667 18717
rect 3050 18640 3056 18692
rect 3108 18680 3114 18692
rect 3145 18683 3203 18689
rect 3145 18680 3157 18683
rect 3108 18652 3157 18680
rect 3108 18640 3114 18652
rect 3145 18649 3157 18652
rect 3191 18649 3203 18683
rect 5166 18680 5172 18692
rect 3145 18643 3203 18649
rect 4172 18652 5172 18680
rect 1673 18615 1731 18621
rect 1673 18581 1685 18615
rect 1719 18612 1731 18615
rect 4172 18612 4200 18652
rect 5166 18640 5172 18652
rect 5224 18640 5230 18692
rect 5626 18640 5632 18692
rect 5684 18640 5690 18692
rect 10594 18680 10600 18692
rect 6472 18652 9352 18680
rect 10555 18652 10600 18680
rect 1719 18584 4200 18612
rect 4249 18615 4307 18621
rect 1719 18581 1731 18584
rect 1673 18575 1731 18581
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 6472 18612 6500 18652
rect 4295 18584 6500 18612
rect 7193 18615 7251 18621
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 7193 18581 7205 18615
rect 7239 18612 7251 18615
rect 8938 18612 8944 18624
rect 7239 18584 8944 18612
rect 7239 18581 7251 18584
rect 7193 18575 7251 18581
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 9324 18612 9352 18652
rect 10594 18640 10600 18652
rect 10652 18640 10658 18692
rect 11624 18680 11652 18711
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 10796 18652 11652 18680
rect 13096 18680 13124 18788
rect 13173 18785 13185 18819
rect 13219 18816 13231 18819
rect 13262 18816 13268 18828
rect 13219 18788 13268 18816
rect 13219 18785 13231 18788
rect 13173 18779 13231 18785
rect 13262 18776 13268 18788
rect 13320 18776 13326 18828
rect 15562 18816 15568 18828
rect 15523 18788 15568 18816
rect 15562 18776 15568 18788
rect 15620 18776 15626 18828
rect 17218 18816 17224 18828
rect 17179 18788 17224 18816
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 18693 18819 18751 18825
rect 18693 18785 18705 18819
rect 18739 18816 18751 18819
rect 19426 18816 19432 18828
rect 18739 18788 19432 18816
rect 18739 18785 18751 18788
rect 18693 18779 18751 18785
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 19889 18819 19947 18825
rect 19889 18785 19901 18819
rect 19935 18816 19947 18819
rect 22097 18819 22155 18825
rect 22097 18816 22109 18819
rect 19935 18788 22109 18816
rect 19935 18785 19947 18788
rect 19889 18779 19947 18785
rect 22097 18785 22109 18788
rect 22143 18785 22155 18819
rect 24026 18816 24032 18828
rect 23987 18788 24032 18816
rect 22097 18779 22155 18785
rect 24026 18776 24032 18788
rect 24084 18776 24090 18828
rect 24670 18816 24676 18828
rect 24631 18788 24676 18816
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 25314 18816 25320 18828
rect 25275 18788 25320 18816
rect 25314 18776 25320 18788
rect 25372 18776 25378 18828
rect 13354 18748 13360 18760
rect 13315 18720 13360 18748
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 14826 18748 14832 18760
rect 13464 18720 14832 18748
rect 13464 18680 13492 18720
rect 14826 18708 14832 18720
rect 14884 18708 14890 18760
rect 18874 18748 18880 18760
rect 18835 18720 18880 18748
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 20073 18751 20131 18757
rect 20073 18748 20085 18751
rect 20036 18720 20085 18748
rect 20036 18708 20042 18720
rect 20073 18717 20085 18720
rect 20119 18717 20131 18751
rect 20073 18711 20131 18717
rect 20717 18751 20775 18757
rect 20717 18717 20729 18751
rect 20763 18748 20775 18751
rect 20898 18748 20904 18760
rect 20763 18720 20904 18748
rect 20763 18717 20775 18720
rect 20717 18711 20775 18717
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 20990 18708 20996 18760
rect 21048 18748 21054 18760
rect 21545 18751 21603 18757
rect 21545 18748 21557 18751
rect 21048 18720 21557 18748
rect 21048 18708 21054 18720
rect 21545 18717 21557 18720
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 22005 18751 22063 18757
rect 22005 18717 22017 18751
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 25961 18751 26019 18757
rect 25961 18717 25973 18751
rect 26007 18717 26019 18751
rect 26602 18748 26608 18760
rect 26563 18720 26608 18748
rect 25961 18711 26019 18717
rect 13096 18652 13492 18680
rect 10796 18624 10824 18652
rect 13814 18640 13820 18692
rect 13872 18680 13878 18692
rect 15841 18683 15899 18689
rect 15841 18680 15853 18683
rect 13872 18652 15853 18680
rect 13872 18640 13878 18652
rect 15841 18649 15853 18652
rect 15887 18649 15899 18683
rect 15841 18643 15899 18649
rect 15933 18683 15991 18689
rect 15933 18649 15945 18683
rect 15979 18649 15991 18683
rect 16574 18680 16580 18692
rect 16535 18652 16580 18680
rect 15933 18643 15991 18649
rect 10686 18612 10692 18624
rect 9324 18584 10692 18612
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 10778 18572 10784 18624
rect 10836 18572 10842 18624
rect 12253 18615 12311 18621
rect 12253 18581 12265 18615
rect 12299 18612 12311 18615
rect 12342 18612 12348 18624
rect 12299 18584 12348 18612
rect 12299 18581 12311 18584
rect 12253 18575 12311 18581
rect 12342 18572 12348 18584
rect 12400 18572 12406 18624
rect 15948 18612 15976 18643
rect 16574 18640 16580 18652
rect 16632 18640 16638 18692
rect 16666 18640 16672 18692
rect 16724 18680 16730 18692
rect 20916 18680 20944 18708
rect 22020 18680 22048 18711
rect 23382 18680 23388 18692
rect 16724 18652 16769 18680
rect 20916 18652 22048 18680
rect 23343 18652 23388 18680
rect 16724 18640 16730 18652
rect 23382 18640 23388 18652
rect 23440 18640 23446 18692
rect 23477 18683 23535 18689
rect 23477 18649 23489 18683
rect 23523 18649 23535 18683
rect 24762 18680 24768 18692
rect 24723 18652 24768 18680
rect 23477 18643 23535 18649
rect 20714 18612 20720 18624
rect 15948 18584 20720 18612
rect 20714 18572 20720 18584
rect 20772 18572 20778 18624
rect 22646 18612 22652 18624
rect 22607 18584 22652 18612
rect 22646 18572 22652 18584
rect 22704 18572 22710 18624
rect 23492 18612 23520 18643
rect 24762 18640 24768 18652
rect 24820 18640 24826 18692
rect 25130 18640 25136 18692
rect 25188 18680 25194 18692
rect 25976 18680 26004 18711
rect 26602 18708 26608 18720
rect 26660 18708 26666 18760
rect 31113 18751 31171 18757
rect 31113 18717 31125 18751
rect 31159 18748 31171 18751
rect 38286 18748 38292 18760
rect 31159 18720 35894 18748
rect 38247 18720 38292 18748
rect 31159 18717 31171 18720
rect 31113 18711 31171 18717
rect 25188 18652 26004 18680
rect 25188 18640 25194 18652
rect 24854 18612 24860 18624
rect 23492 18584 24860 18612
rect 24854 18572 24860 18584
rect 24912 18572 24918 18624
rect 35866 18612 35894 18720
rect 38286 18708 38292 18720
rect 38344 18708 38350 18760
rect 38105 18615 38163 18621
rect 38105 18612 38117 18615
rect 35866 18584 38117 18612
rect 38105 18581 38117 18584
rect 38151 18581 38163 18615
rect 38105 18575 38163 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 3234 18368 3240 18420
rect 3292 18408 3298 18420
rect 3973 18411 4031 18417
rect 3973 18408 3985 18411
rect 3292 18380 3985 18408
rect 3292 18368 3298 18380
rect 3973 18377 3985 18380
rect 4019 18377 4031 18411
rect 3973 18371 4031 18377
rect 4430 18368 4436 18420
rect 4488 18408 4494 18420
rect 7190 18408 7196 18420
rect 4488 18380 7196 18408
rect 4488 18368 4494 18380
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 8294 18368 8300 18420
rect 8352 18408 8358 18420
rect 8754 18408 8760 18420
rect 8352 18380 8760 18408
rect 8352 18368 8358 18380
rect 8754 18368 8760 18380
rect 8812 18368 8818 18420
rect 8849 18411 8907 18417
rect 8849 18377 8861 18411
rect 8895 18408 8907 18411
rect 10226 18408 10232 18420
rect 8895 18380 10232 18408
rect 8895 18377 8907 18380
rect 8849 18371 8907 18377
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 12345 18411 12403 18417
rect 12345 18377 12357 18411
rect 12391 18408 12403 18411
rect 14553 18411 14611 18417
rect 12391 18380 14504 18408
rect 12391 18377 12403 18380
rect 12345 18371 12403 18377
rect 3510 18340 3516 18352
rect 3174 18312 3516 18340
rect 3510 18300 3516 18312
rect 3568 18300 3574 18352
rect 4706 18300 4712 18352
rect 4764 18300 4770 18352
rect 5350 18300 5356 18352
rect 5408 18340 5414 18352
rect 5408 18312 6946 18340
rect 5408 18300 5414 18312
rect 8202 18300 8208 18352
rect 8260 18340 8266 18352
rect 8260 18312 8432 18340
rect 8260 18300 8266 18312
rect 5718 18232 5724 18284
rect 5776 18272 5782 18284
rect 8404 18281 8432 18312
rect 8938 18300 8944 18352
rect 8996 18340 9002 18352
rect 8996 18312 9154 18340
rect 8996 18300 9002 18312
rect 10042 18300 10048 18352
rect 10100 18340 10106 18352
rect 10100 18312 10640 18340
rect 10100 18300 10106 18312
rect 10612 18281 10640 18312
rect 10686 18300 10692 18352
rect 10744 18340 10750 18352
rect 10744 18312 11928 18340
rect 10744 18300 10750 18312
rect 8389 18275 8447 18281
rect 5776 18244 5821 18272
rect 5776 18232 5782 18244
rect 8389 18241 8401 18275
rect 8435 18241 8447 18275
rect 8389 18235 8447 18241
rect 10597 18275 10655 18281
rect 10597 18241 10609 18275
rect 10643 18272 10655 18275
rect 10870 18272 10876 18284
rect 10643 18244 10876 18272
rect 10643 18241 10655 18244
rect 10597 18235 10655 18241
rect 1670 18204 1676 18216
rect 1631 18176 1676 18204
rect 1670 18164 1676 18176
rect 1728 18164 1734 18216
rect 1949 18207 2007 18213
rect 1949 18173 1961 18207
rect 1995 18204 2007 18207
rect 2038 18204 2044 18216
rect 1995 18176 2044 18204
rect 1995 18173 2007 18176
rect 1949 18167 2007 18173
rect 2038 18164 2044 18176
rect 2096 18204 2102 18216
rect 5445 18207 5503 18213
rect 2096 18176 4476 18204
rect 2096 18164 2102 18176
rect 3418 18068 3424 18080
rect 3379 18040 3424 18068
rect 3418 18028 3424 18040
rect 3476 18028 3482 18080
rect 3786 18028 3792 18080
rect 3844 18068 3850 18080
rect 4154 18068 4160 18080
rect 3844 18040 4160 18068
rect 3844 18028 3850 18040
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 4448 18068 4476 18176
rect 5445 18173 5457 18207
rect 5491 18204 5503 18207
rect 6086 18204 6092 18216
rect 5491 18176 6092 18204
rect 5491 18173 5503 18176
rect 5445 18167 5503 18173
rect 6086 18164 6092 18176
rect 6144 18164 6150 18216
rect 6638 18204 6644 18216
rect 6551 18176 6644 18204
rect 6638 18164 6644 18176
rect 6696 18204 6702 18216
rect 7466 18204 7472 18216
rect 6696 18176 7472 18204
rect 6696 18164 6702 18176
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 8110 18204 8116 18216
rect 8071 18176 8116 18204
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 8404 18204 8432 18235
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 11900 18281 11928 18312
rect 12618 18300 12624 18352
rect 12676 18340 12682 18352
rect 13357 18343 13415 18349
rect 13357 18340 13369 18343
rect 12676 18312 13369 18340
rect 12676 18300 12682 18312
rect 13357 18309 13369 18312
rect 13403 18309 13415 18343
rect 13357 18303 13415 18309
rect 13446 18300 13452 18352
rect 13504 18340 13510 18352
rect 14476 18340 14504 18380
rect 14553 18377 14565 18411
rect 14599 18408 14611 18411
rect 15746 18408 15752 18420
rect 14599 18380 15752 18408
rect 14599 18377 14611 18380
rect 14553 18371 14611 18377
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 16301 18411 16359 18417
rect 16301 18377 16313 18411
rect 16347 18408 16359 18411
rect 16574 18408 16580 18420
rect 16347 18380 16580 18408
rect 16347 18377 16359 18380
rect 16301 18371 16359 18377
rect 16574 18368 16580 18380
rect 16632 18408 16638 18420
rect 17497 18411 17555 18417
rect 17497 18408 17509 18411
rect 16632 18380 17509 18408
rect 16632 18368 16638 18380
rect 17497 18377 17509 18380
rect 17543 18377 17555 18411
rect 17497 18371 17555 18377
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19521 18411 19579 18417
rect 19521 18408 19533 18411
rect 19392 18380 19533 18408
rect 19392 18368 19398 18380
rect 19521 18377 19533 18380
rect 19567 18377 19579 18411
rect 19521 18371 19579 18377
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 20036 18380 22094 18408
rect 20036 18368 20042 18380
rect 17310 18340 17316 18352
rect 13504 18312 13549 18340
rect 14476 18312 17316 18340
rect 13504 18300 13510 18312
rect 17310 18300 17316 18312
rect 17368 18300 17374 18352
rect 17586 18300 17592 18352
rect 17644 18340 17650 18352
rect 18325 18343 18383 18349
rect 18325 18340 18337 18343
rect 17644 18312 18337 18340
rect 17644 18300 17650 18312
rect 18325 18309 18337 18312
rect 18371 18309 18383 18343
rect 22066 18340 22094 18380
rect 22370 18368 22376 18420
rect 22428 18408 22434 18420
rect 22649 18411 22707 18417
rect 22649 18408 22661 18411
rect 22428 18380 22661 18408
rect 22428 18368 22434 18380
rect 22649 18377 22661 18380
rect 22695 18408 22707 18411
rect 23382 18408 23388 18420
rect 22695 18380 23388 18408
rect 22695 18377 22707 18380
rect 22649 18371 22707 18377
rect 23382 18368 23388 18380
rect 23440 18368 23446 18420
rect 24305 18411 24363 18417
rect 24305 18377 24317 18411
rect 24351 18408 24363 18411
rect 24670 18408 24676 18420
rect 24351 18380 24676 18408
rect 24351 18377 24363 18380
rect 24305 18371 24363 18377
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 24762 18368 24768 18420
rect 24820 18408 24826 18420
rect 26145 18411 26203 18417
rect 26145 18408 26157 18411
rect 24820 18380 26157 18408
rect 24820 18368 24826 18380
rect 26145 18377 26157 18380
rect 26191 18377 26203 18411
rect 26145 18371 26203 18377
rect 28994 18340 29000 18352
rect 22066 18312 29000 18340
rect 18325 18303 18383 18309
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18241 11943 18275
rect 15013 18275 15071 18281
rect 15013 18272 15025 18275
rect 11885 18235 11943 18241
rect 14844 18244 15025 18272
rect 9674 18204 9680 18216
rect 8404 18176 9680 18204
rect 9674 18164 9680 18176
rect 9732 18204 9738 18216
rect 9950 18204 9956 18216
rect 9732 18176 9956 18204
rect 9732 18164 9738 18176
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 10318 18204 10324 18216
rect 10279 18176 10324 18204
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 11112 18176 11713 18204
rect 11112 18164 11118 18176
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 11701 18167 11759 18173
rect 5644 18108 6776 18136
rect 5644 18068 5672 18108
rect 4448 18040 5672 18068
rect 6748 18068 6776 18108
rect 8404 18108 8984 18136
rect 8404 18068 8432 18108
rect 6748 18040 8432 18068
rect 8956 18068 8984 18108
rect 12802 18096 12808 18148
rect 12860 18136 12866 18148
rect 12897 18139 12955 18145
rect 12897 18136 12909 18139
rect 12860 18108 12909 18136
rect 12860 18096 12866 18108
rect 12897 18105 12909 18108
rect 12943 18105 12955 18139
rect 12897 18099 12955 18105
rect 14844 18068 14872 18244
rect 15013 18241 15025 18244
rect 15059 18272 15071 18275
rect 16758 18272 16764 18284
rect 15059 18244 16764 18272
rect 15059 18241 15071 18244
rect 15013 18235 15071 18241
rect 16758 18232 16764 18244
rect 16816 18272 16822 18284
rect 17862 18272 17868 18284
rect 16816 18244 17868 18272
rect 16816 18232 16822 18244
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20806 18272 20812 18284
rect 20027 18244 20812 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 21266 18272 21272 18284
rect 21227 18244 21272 18272
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 21453 18275 21511 18281
rect 21453 18241 21465 18275
rect 21499 18272 21511 18275
rect 22646 18272 22652 18284
rect 21499 18244 22652 18272
rect 21499 18241 21511 18244
rect 21453 18235 21511 18241
rect 22646 18232 22652 18244
rect 22704 18232 22710 18284
rect 23676 18281 23704 18312
rect 28994 18300 29000 18312
rect 29052 18300 29058 18352
rect 23661 18275 23719 18281
rect 23661 18241 23673 18275
rect 23707 18241 23719 18275
rect 24946 18272 24952 18284
rect 24907 18244 24952 18272
rect 23661 18235 23719 18241
rect 24946 18232 24952 18244
rect 25004 18232 25010 18284
rect 25590 18272 25596 18284
rect 25551 18244 25596 18272
rect 25590 18232 25596 18244
rect 25648 18232 25654 18284
rect 26234 18272 26240 18284
rect 26195 18244 26240 18272
rect 26234 18232 26240 18244
rect 26292 18232 26298 18284
rect 34333 18275 34391 18281
rect 34333 18241 34345 18275
rect 34379 18272 34391 18275
rect 35526 18272 35532 18284
rect 34379 18244 35532 18272
rect 34379 18241 34391 18244
rect 34333 18235 34391 18241
rect 35526 18232 35532 18244
rect 35584 18232 35590 18284
rect 15286 18164 15292 18216
rect 15344 18204 15350 18216
rect 15657 18207 15715 18213
rect 15657 18204 15669 18207
rect 15344 18176 15669 18204
rect 15344 18164 15350 18176
rect 15657 18173 15669 18176
rect 15703 18173 15715 18207
rect 15657 18167 15715 18173
rect 15746 18164 15752 18216
rect 15804 18204 15810 18216
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15804 18176 15853 18204
rect 15804 18164 15810 18176
rect 15841 18173 15853 18176
rect 15887 18173 15899 18207
rect 16850 18204 16856 18216
rect 16811 18176 16856 18204
rect 15841 18167 15899 18173
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 17034 18204 17040 18216
rect 16995 18176 17040 18204
rect 17034 18164 17040 18176
rect 17092 18164 17098 18216
rect 18233 18207 18291 18213
rect 18233 18204 18245 18207
rect 18156 18176 18245 18204
rect 18156 18148 18184 18176
rect 18233 18173 18245 18176
rect 18279 18173 18291 18207
rect 18506 18204 18512 18216
rect 18467 18176 18512 18204
rect 18233 18167 18291 18173
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 18874 18164 18880 18216
rect 18932 18204 18938 18216
rect 20165 18207 20223 18213
rect 20165 18204 20177 18207
rect 18932 18176 20177 18204
rect 18932 18164 18938 18176
rect 20165 18173 20177 18176
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 18138 18096 18144 18148
rect 18196 18096 18202 18148
rect 20180 18136 20208 18167
rect 21358 18164 21364 18216
rect 21416 18204 21422 18216
rect 22005 18207 22063 18213
rect 22005 18204 22017 18207
rect 21416 18176 22017 18204
rect 21416 18164 21422 18176
rect 22005 18173 22017 18176
rect 22051 18173 22063 18207
rect 22005 18167 22063 18173
rect 22189 18207 22247 18213
rect 22189 18173 22201 18207
rect 22235 18204 22247 18207
rect 22278 18204 22284 18216
rect 22235 18176 22284 18204
rect 22235 18173 22247 18176
rect 22189 18167 22247 18173
rect 22278 18164 22284 18176
rect 22336 18164 22342 18216
rect 23845 18207 23903 18213
rect 23845 18173 23857 18207
rect 23891 18204 23903 18207
rect 25501 18207 25559 18213
rect 25501 18204 25513 18207
rect 23891 18176 25513 18204
rect 23891 18173 23903 18176
rect 23845 18167 23903 18173
rect 25501 18173 25513 18176
rect 25547 18173 25559 18207
rect 25501 18167 25559 18173
rect 25038 18136 25044 18148
rect 20180 18108 25044 18136
rect 25038 18096 25044 18108
rect 25096 18096 25102 18148
rect 8956 18040 14872 18068
rect 15105 18071 15163 18077
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 16482 18068 16488 18080
rect 15151 18040 16488 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20809 18071 20867 18077
rect 20809 18068 20821 18071
rect 20772 18040 20821 18068
rect 20772 18028 20778 18040
rect 20809 18037 20821 18040
rect 20855 18037 20867 18071
rect 24762 18068 24768 18080
rect 24723 18040 24768 18068
rect 20809 18031 20867 18037
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 34238 18068 34244 18080
rect 34199 18040 34244 18068
rect 34238 18028 34244 18040
rect 34296 18028 34302 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1581 17867 1639 17873
rect 1581 17833 1593 17867
rect 1627 17864 1639 17867
rect 4065 17867 4123 17873
rect 1627 17836 4016 17864
rect 1627 17833 1639 17836
rect 1581 17827 1639 17833
rect 3988 17796 4016 17836
rect 4065 17833 4077 17867
rect 4111 17864 4123 17867
rect 8570 17864 8576 17876
rect 4111 17836 7788 17864
rect 8531 17836 8576 17864
rect 4111 17833 4123 17836
rect 4065 17827 4123 17833
rect 5350 17796 5356 17808
rect 3988 17768 5356 17796
rect 5350 17756 5356 17768
rect 5408 17756 5414 17808
rect 3329 17731 3387 17737
rect 3329 17697 3341 17731
rect 3375 17728 3387 17731
rect 4798 17728 4804 17740
rect 3375 17700 4804 17728
rect 3375 17697 3387 17700
rect 3329 17691 3387 17697
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 6641 17731 6699 17737
rect 6641 17697 6653 17731
rect 6687 17728 6699 17731
rect 7374 17728 7380 17740
rect 6687 17700 7380 17728
rect 6687 17697 6699 17700
rect 6641 17691 6699 17697
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 7760 17728 7788 17836
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 8662 17824 8668 17876
rect 8720 17864 8726 17876
rect 17497 17867 17555 17873
rect 8720 17836 15608 17864
rect 8720 17824 8726 17836
rect 7834 17756 7840 17808
rect 7892 17796 7898 17808
rect 8754 17796 8760 17808
rect 7892 17768 8760 17796
rect 7892 17756 7898 17768
rect 8754 17756 8760 17768
rect 8812 17796 8818 17808
rect 9125 17799 9183 17805
rect 9125 17796 9137 17799
rect 8812 17768 9137 17796
rect 8812 17756 8818 17768
rect 9125 17765 9137 17768
rect 9171 17765 9183 17799
rect 9125 17759 9183 17765
rect 11256 17768 11560 17796
rect 11256 17728 11284 17768
rect 11422 17728 11428 17740
rect 7760 17700 11284 17728
rect 11383 17700 11428 17728
rect 11422 17688 11428 17700
rect 11480 17688 11486 17740
rect 11532 17728 11560 17768
rect 11698 17756 11704 17808
rect 11756 17796 11762 17808
rect 14277 17799 14335 17805
rect 14277 17796 14289 17799
rect 11756 17768 14289 17796
rect 11756 17756 11762 17768
rect 14277 17765 14289 17768
rect 14323 17765 14335 17799
rect 14277 17759 14335 17765
rect 12618 17728 12624 17740
rect 11532 17700 12624 17728
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 15010 17688 15016 17740
rect 15068 17728 15074 17740
rect 15473 17731 15531 17737
rect 15473 17728 15485 17731
rect 15068 17700 15485 17728
rect 15068 17688 15074 17700
rect 15473 17697 15485 17700
rect 15519 17697 15531 17731
rect 15580 17728 15608 17836
rect 17497 17833 17509 17867
rect 17543 17864 17555 17867
rect 17770 17864 17776 17876
rect 17543 17836 17776 17864
rect 17543 17833 17555 17836
rect 17497 17827 17555 17833
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 22281 17867 22339 17873
rect 22281 17833 22293 17867
rect 22327 17864 22339 17867
rect 22370 17864 22376 17876
rect 22327 17836 22376 17864
rect 22327 17833 22339 17836
rect 22281 17827 22339 17833
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 23106 17864 23112 17876
rect 23067 17836 23112 17864
rect 23106 17824 23112 17836
rect 23164 17824 23170 17876
rect 24765 17867 24823 17873
rect 24765 17833 24777 17867
rect 24811 17864 24823 17867
rect 24946 17864 24952 17876
rect 24811 17836 24952 17864
rect 24811 17833 24823 17836
rect 24765 17827 24823 17833
rect 24946 17824 24952 17836
rect 25004 17824 25010 17876
rect 25409 17867 25467 17873
rect 25409 17833 25421 17867
rect 25455 17864 25467 17867
rect 26602 17864 26608 17876
rect 25455 17836 26608 17864
rect 25455 17833 25467 17836
rect 25409 17827 25467 17833
rect 26602 17824 26608 17836
rect 26660 17824 26666 17876
rect 16025 17799 16083 17805
rect 16025 17765 16037 17799
rect 16071 17796 16083 17799
rect 18506 17796 18512 17808
rect 16071 17768 18512 17796
rect 16071 17765 16083 17768
rect 16025 17759 16083 17765
rect 18506 17756 18512 17768
rect 18564 17796 18570 17808
rect 18564 17768 29776 17796
rect 18564 17756 18570 17768
rect 16761 17731 16819 17737
rect 15580 17700 16160 17728
rect 15473 17691 15531 17697
rect 3418 17620 3424 17672
rect 3476 17660 3482 17672
rect 3970 17660 3976 17672
rect 3476 17632 3976 17660
rect 3476 17620 3482 17632
rect 3970 17620 3976 17632
rect 4028 17620 4034 17672
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 1762 17552 1768 17604
rect 1820 17592 1826 17604
rect 3053 17595 3111 17601
rect 1820 17564 1886 17592
rect 1820 17552 1826 17564
rect 3053 17561 3065 17595
rect 3099 17592 3111 17595
rect 3694 17592 3700 17604
rect 3099 17564 3700 17592
rect 3099 17561 3111 17564
rect 3053 17555 3111 17561
rect 3694 17552 3700 17564
rect 3752 17552 3758 17604
rect 3418 17484 3424 17536
rect 3476 17524 3482 17536
rect 3786 17524 3792 17536
rect 3476 17496 3792 17524
rect 3476 17484 3482 17496
rect 3786 17484 3792 17496
rect 3844 17484 3850 17536
rect 3988 17524 4016 17620
rect 4614 17592 4620 17604
rect 4575 17564 4620 17592
rect 4614 17552 4620 17564
rect 4672 17552 4678 17604
rect 5074 17552 5080 17604
rect 5132 17592 5138 17604
rect 6362 17592 6368 17604
rect 5132 17564 5198 17592
rect 6323 17564 6368 17592
rect 5132 17552 5138 17564
rect 6362 17552 6368 17564
rect 6420 17552 6426 17604
rect 7300 17592 7328 17623
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7524 17632 7941 17660
rect 7524 17620 7530 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8397 17663 8455 17669
rect 8397 17629 8409 17663
rect 8443 17662 8455 17663
rect 8443 17634 8524 17662
rect 8443 17629 8455 17634
rect 8397 17623 8455 17629
rect 6472 17564 7328 17592
rect 7944 17592 7972 17623
rect 8496 17604 8524 17634
rect 10870 17620 10876 17672
rect 10928 17660 10934 17672
rect 10928 17632 10973 17660
rect 10928 17620 10934 17632
rect 14090 17620 14096 17672
rect 14148 17660 14154 17672
rect 14737 17663 14795 17669
rect 14737 17660 14749 17663
rect 14148 17632 14749 17660
rect 14148 17620 14154 17632
rect 14737 17629 14749 17632
rect 14783 17629 14795 17663
rect 14918 17660 14924 17672
rect 14879 17632 14924 17660
rect 14737 17623 14795 17629
rect 14918 17620 14924 17632
rect 14976 17660 14982 17672
rect 15286 17660 15292 17672
rect 14976 17632 15292 17660
rect 14976 17620 14982 17632
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 8294 17592 8300 17604
rect 7944 17564 8300 17592
rect 6472 17524 6500 17564
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 8478 17552 8484 17604
rect 8536 17552 8542 17604
rect 8570 17552 8576 17604
rect 8628 17592 8634 17604
rect 8628 17564 9430 17592
rect 8628 17552 8634 17564
rect 10502 17552 10508 17604
rect 10560 17592 10566 17604
rect 10597 17595 10655 17601
rect 10597 17592 10609 17595
rect 10560 17564 10609 17592
rect 10560 17552 10566 17564
rect 10597 17561 10609 17564
rect 10643 17561 10655 17595
rect 10597 17555 10655 17561
rect 11146 17552 11152 17604
rect 11204 17592 11210 17604
rect 11517 17595 11575 17601
rect 11517 17592 11529 17595
rect 11204 17564 11529 17592
rect 11204 17552 11210 17564
rect 11517 17561 11529 17564
rect 11563 17561 11575 17595
rect 11517 17555 11575 17561
rect 12069 17595 12127 17601
rect 12069 17561 12081 17595
rect 12115 17592 12127 17595
rect 12158 17592 12164 17604
rect 12115 17564 12164 17592
rect 12115 17561 12127 17564
rect 12069 17555 12127 17561
rect 12158 17552 12164 17564
rect 12216 17552 12222 17604
rect 12802 17552 12808 17604
rect 12860 17592 12866 17604
rect 12989 17595 13047 17601
rect 12989 17592 13001 17595
rect 12860 17564 13001 17592
rect 12860 17552 12866 17564
rect 12989 17561 13001 17564
rect 13035 17561 13047 17595
rect 13538 17592 13544 17604
rect 13499 17564 13544 17592
rect 12989 17555 13047 17561
rect 13538 17552 13544 17564
rect 13596 17552 13602 17604
rect 13633 17595 13691 17601
rect 13633 17561 13645 17595
rect 13679 17561 13691 17595
rect 15562 17592 15568 17604
rect 15523 17564 15568 17592
rect 13633 17555 13691 17561
rect 7098 17524 7104 17536
rect 3988 17496 6500 17524
rect 7059 17496 7104 17524
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 7190 17484 7196 17536
rect 7248 17524 7254 17536
rect 7745 17527 7803 17533
rect 7745 17524 7757 17527
rect 7248 17496 7757 17524
rect 7248 17484 7254 17496
rect 7745 17493 7757 17496
rect 7791 17493 7803 17527
rect 7745 17487 7803 17493
rect 7834 17484 7840 17536
rect 7892 17524 7898 17536
rect 10226 17524 10232 17536
rect 7892 17496 10232 17524
rect 7892 17484 7898 17496
rect 10226 17484 10232 17496
rect 10284 17484 10290 17536
rect 13170 17484 13176 17536
rect 13228 17524 13234 17536
rect 13446 17524 13452 17536
rect 13228 17496 13452 17524
rect 13228 17484 13234 17496
rect 13446 17484 13452 17496
rect 13504 17484 13510 17536
rect 13648 17524 13676 17555
rect 15562 17552 15568 17564
rect 15620 17552 15626 17604
rect 16132 17592 16160 17700
rect 16761 17697 16773 17731
rect 16807 17728 16819 17731
rect 18417 17731 18475 17737
rect 18417 17728 18429 17731
rect 16807 17700 18429 17728
rect 16807 17697 16819 17700
rect 16761 17691 16819 17697
rect 18417 17697 18429 17700
rect 18463 17697 18475 17731
rect 18417 17691 18475 17697
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17728 18659 17731
rect 19978 17728 19984 17740
rect 18647 17700 19984 17728
rect 18647 17697 18659 17700
rect 18601 17691 18659 17697
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 20898 17728 20904 17740
rect 20364 17700 20904 17728
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 16942 17660 16948 17672
rect 16715 17632 16948 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 17310 17660 17316 17672
rect 17271 17632 17316 17660
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17660 19855 17663
rect 20364 17660 20392 17700
rect 20898 17688 20904 17700
rect 20956 17688 20962 17740
rect 21177 17731 21235 17737
rect 21177 17697 21189 17731
rect 21223 17728 21235 17731
rect 22370 17728 22376 17740
rect 21223 17700 22376 17728
rect 21223 17697 21235 17700
rect 21177 17691 21235 17697
rect 22370 17688 22376 17700
rect 22428 17688 22434 17740
rect 22465 17731 22523 17737
rect 22465 17697 22477 17731
rect 22511 17728 22523 17731
rect 24762 17728 24768 17740
rect 22511 17700 24768 17728
rect 22511 17697 22523 17700
rect 22465 17691 22523 17697
rect 24762 17688 24768 17700
rect 24820 17688 24826 17740
rect 22646 17660 22652 17672
rect 19843 17632 20392 17660
rect 22607 17632 22652 17660
rect 19843 17629 19855 17632
rect 19797 17623 19855 17629
rect 19812 17592 19840 17623
rect 22646 17620 22652 17632
rect 22704 17620 22710 17672
rect 23566 17660 23572 17672
rect 23527 17632 23572 17660
rect 23566 17620 23572 17632
rect 23624 17620 23630 17672
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17629 23811 17663
rect 23753 17623 23811 17629
rect 20530 17592 20536 17604
rect 16132 17564 19840 17592
rect 20491 17564 20536 17592
rect 20530 17552 20536 17564
rect 20588 17552 20594 17604
rect 20625 17595 20683 17601
rect 20625 17561 20637 17595
rect 20671 17592 20683 17595
rect 21450 17592 21456 17604
rect 20671 17564 21456 17592
rect 20671 17561 20683 17564
rect 20625 17555 20683 17561
rect 21450 17552 21456 17564
rect 21508 17552 21514 17604
rect 23768 17592 23796 17623
rect 23842 17620 23848 17672
rect 23900 17660 23906 17672
rect 24581 17663 24639 17669
rect 24581 17660 24593 17663
rect 23900 17632 24593 17660
rect 23900 17620 23906 17632
rect 24581 17629 24593 17632
rect 24627 17660 24639 17663
rect 25130 17660 25136 17672
rect 24627 17632 25136 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 25130 17620 25136 17632
rect 25188 17620 25194 17672
rect 25225 17663 25283 17669
rect 25225 17629 25237 17663
rect 25271 17660 25283 17663
rect 25590 17660 25596 17672
rect 25271 17632 25596 17660
rect 25271 17629 25283 17632
rect 25225 17623 25283 17629
rect 25590 17620 25596 17632
rect 25648 17660 25654 17672
rect 26142 17660 26148 17672
rect 25648 17632 26148 17660
rect 25648 17620 25654 17632
rect 26142 17620 26148 17632
rect 26200 17620 26206 17672
rect 29748 17669 29776 17768
rect 29733 17663 29791 17669
rect 29733 17629 29745 17663
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 34790 17592 34796 17604
rect 23768 17564 34796 17592
rect 34790 17552 34796 17564
rect 34848 17552 34854 17604
rect 17770 17524 17776 17536
rect 13648 17496 17776 17524
rect 17770 17484 17776 17496
rect 17828 17484 17834 17536
rect 17957 17527 18015 17533
rect 17957 17493 17969 17527
rect 18003 17524 18015 17527
rect 18138 17524 18144 17536
rect 18003 17496 18144 17524
rect 18003 17493 18015 17496
rect 17957 17487 18015 17493
rect 18138 17484 18144 17496
rect 18196 17484 18202 17536
rect 19889 17527 19947 17533
rect 19889 17493 19901 17527
rect 19935 17524 19947 17527
rect 21266 17524 21272 17536
rect 19935 17496 21272 17524
rect 19935 17493 19947 17496
rect 19889 17487 19947 17493
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 25498 17484 25504 17536
rect 25556 17524 25562 17536
rect 25869 17527 25927 17533
rect 25869 17524 25881 17527
rect 25556 17496 25881 17524
rect 25556 17484 25562 17496
rect 25869 17493 25881 17496
rect 25915 17493 25927 17527
rect 25869 17487 25927 17493
rect 29825 17527 29883 17533
rect 29825 17493 29837 17527
rect 29871 17524 29883 17527
rect 33778 17524 33784 17536
rect 29871 17496 33784 17524
rect 29871 17493 29883 17496
rect 29825 17487 29883 17493
rect 33778 17484 33784 17496
rect 33836 17484 33842 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 8662 17320 8668 17332
rect 2148 17292 8668 17320
rect 2148 17264 2176 17292
rect 8662 17280 8668 17292
rect 8720 17280 8726 17332
rect 8938 17280 8944 17332
rect 8996 17320 9002 17332
rect 8996 17292 10088 17320
rect 8996 17280 9002 17292
rect 2130 17252 2136 17264
rect 2091 17224 2136 17252
rect 2130 17212 2136 17224
rect 2188 17212 2194 17264
rect 3142 17212 3148 17264
rect 3200 17212 3206 17264
rect 3786 17212 3792 17264
rect 3844 17252 3850 17264
rect 7006 17252 7012 17264
rect 3844 17224 7012 17252
rect 3844 17212 3850 17224
rect 7006 17212 7012 17224
rect 7064 17212 7070 17264
rect 7650 17212 7656 17264
rect 7708 17252 7714 17264
rect 7708 17224 8142 17252
rect 7708 17212 7714 17224
rect 9398 17212 9404 17264
rect 9456 17252 9462 17264
rect 10060 17261 10088 17292
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10284 17292 22094 17320
rect 10284 17280 10290 17292
rect 9953 17255 10011 17261
rect 9953 17252 9965 17255
rect 9456 17224 9965 17252
rect 9456 17212 9462 17224
rect 9953 17221 9965 17224
rect 9999 17221 10011 17255
rect 9953 17215 10011 17221
rect 10045 17255 10103 17261
rect 10045 17221 10057 17255
rect 10091 17221 10103 17255
rect 11974 17252 11980 17264
rect 11935 17224 11980 17252
rect 10045 17215 10103 17221
rect 11974 17212 11980 17224
rect 12032 17212 12038 17264
rect 14826 17212 14832 17264
rect 14884 17252 14890 17264
rect 14884 17224 16160 17252
rect 14884 17212 14890 17224
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4798 17184 4804 17196
rect 4203 17156 4804 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 4890 17144 4896 17196
rect 4948 17184 4954 17196
rect 5169 17187 5227 17193
rect 5169 17184 5181 17187
rect 4948 17156 5181 17184
rect 4948 17144 4954 17156
rect 5169 17153 5181 17156
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 6638 17184 6644 17196
rect 5859 17156 6644 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 3878 17116 3884 17128
rect 3384 17088 3884 17116
rect 3384 17076 3390 17088
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 5828 17048 5856 17147
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 7190 17184 7196 17196
rect 6779 17156 7196 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 9490 17184 9496 17196
rect 9180 17156 9496 17184
rect 9180 17144 9186 17156
rect 9490 17144 9496 17156
rect 9548 17144 9554 17196
rect 10870 17144 10876 17196
rect 10928 17184 10934 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 10928 17156 11713 17184
rect 10928 17144 10934 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 13078 17144 13084 17196
rect 13136 17144 13142 17196
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13280 17156 14105 17184
rect 7374 17116 7380 17128
rect 7335 17088 7380 17116
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 7653 17119 7711 17125
rect 7653 17116 7665 17119
rect 7484 17088 7665 17116
rect 4080 17020 5856 17048
rect 4080 16992 4108 17020
rect 6546 17008 6552 17060
rect 6604 17048 6610 17060
rect 7484 17048 7512 17088
rect 7653 17085 7665 17088
rect 7699 17085 7711 17119
rect 10594 17116 10600 17128
rect 7653 17079 7711 17085
rect 8680 17088 10600 17116
rect 6604 17020 7512 17048
rect 6604 17008 6610 17020
rect 4062 16940 4068 16992
rect 4120 16940 4126 16992
rect 5350 16980 5356 16992
rect 5311 16952 5356 16980
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 5997 16983 6055 16989
rect 5997 16949 6009 16983
rect 6043 16980 6055 16983
rect 6638 16980 6644 16992
rect 6043 16952 6644 16980
rect 6043 16949 6055 16952
rect 5997 16943 6055 16949
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 6917 16983 6975 16989
rect 6917 16949 6929 16983
rect 6963 16980 6975 16983
rect 8680 16980 8708 17088
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10686 17076 10692 17128
rect 10744 17116 10750 17128
rect 13280 17116 13308 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 15470 17184 15476 17196
rect 15431 17156 15476 17184
rect 14093 17147 14151 17153
rect 15470 17144 15476 17156
rect 15528 17144 15534 17196
rect 16132 17193 16160 17224
rect 16482 17212 16488 17264
rect 16540 17252 16546 17264
rect 16540 17224 18092 17252
rect 16540 17212 16546 17224
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17153 16175 17187
rect 17218 17184 17224 17196
rect 17179 17156 17224 17184
rect 16117 17147 16175 17153
rect 17218 17144 17224 17156
rect 17276 17144 17282 17196
rect 17862 17184 17868 17196
rect 17823 17156 17868 17184
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 18064 17193 18092 17224
rect 20714 17212 20720 17264
rect 20772 17252 20778 17264
rect 20809 17255 20867 17261
rect 20809 17252 20821 17255
rect 20772 17224 20821 17252
rect 20772 17212 20778 17224
rect 20809 17221 20821 17224
rect 20855 17221 20867 17255
rect 20809 17215 20867 17221
rect 20898 17212 20904 17264
rect 20956 17252 20962 17264
rect 22066 17252 22094 17292
rect 22186 17280 22192 17332
rect 22244 17320 22250 17332
rect 22646 17320 22652 17332
rect 22244 17292 22289 17320
rect 22607 17292 22652 17320
rect 22244 17280 22250 17292
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 26234 17320 26240 17332
rect 24964 17292 26240 17320
rect 24964 17252 24992 17292
rect 26234 17280 26240 17292
rect 26292 17280 26298 17332
rect 33965 17323 34023 17329
rect 33965 17289 33977 17323
rect 34011 17320 34023 17323
rect 34011 17292 35894 17320
rect 34011 17289 34023 17292
rect 33965 17283 34023 17289
rect 25130 17252 25136 17264
rect 20956 17224 21404 17252
rect 22066 17224 24992 17252
rect 25091 17224 25136 17252
rect 20956 17212 20962 17224
rect 18049 17187 18107 17193
rect 18049 17153 18061 17187
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20257 17187 20315 17193
rect 20257 17184 20269 17187
rect 20128 17156 20269 17184
rect 20128 17144 20134 17156
rect 20257 17153 20269 17156
rect 20303 17153 20315 17187
rect 21266 17184 21272 17196
rect 21227 17156 21272 17184
rect 20257 17147 20315 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 21376 17184 21404 17224
rect 25130 17212 25136 17224
rect 25188 17212 25194 17264
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21376 17156 22017 17184
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 26142 17184 26148 17196
rect 26103 17156 26148 17184
rect 22005 17147 22063 17153
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 26252 17184 26280 17280
rect 27341 17187 27399 17193
rect 27341 17184 27353 17187
rect 26252 17156 27353 17184
rect 27341 17153 27353 17156
rect 27387 17153 27399 17187
rect 33778 17184 33784 17196
rect 33739 17156 33784 17184
rect 27341 17147 27399 17153
rect 33778 17144 33784 17156
rect 33836 17144 33842 17196
rect 35866 17184 35894 17292
rect 38013 17187 38071 17193
rect 38013 17184 38025 17187
rect 35866 17156 38025 17184
rect 38013 17153 38025 17156
rect 38059 17153 38071 17187
rect 38013 17147 38071 17153
rect 13446 17116 13452 17128
rect 10744 17088 13308 17116
rect 13407 17088 13452 17116
rect 10744 17076 10750 17088
rect 13446 17076 13452 17088
rect 13504 17076 13510 17128
rect 13909 17119 13967 17125
rect 13909 17085 13921 17119
rect 13955 17116 13967 17119
rect 13998 17116 14004 17128
rect 13955 17088 14004 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 13998 17076 14004 17088
rect 14056 17076 14062 17128
rect 15378 17076 15384 17128
rect 15436 17116 15442 17128
rect 15436 17088 17816 17116
rect 15436 17076 15442 17088
rect 10505 17051 10563 17057
rect 10505 17017 10517 17051
rect 10551 17048 10563 17051
rect 11606 17048 11612 17060
rect 10551 17020 11612 17048
rect 10551 17017 10563 17020
rect 10505 17011 10563 17017
rect 11606 17008 11612 17020
rect 11664 17008 11670 17060
rect 14277 17051 14335 17057
rect 14277 17048 14289 17051
rect 13372 17020 14289 17048
rect 9122 16980 9128 16992
rect 6963 16952 8708 16980
rect 9083 16952 9128 16980
rect 6963 16949 6975 16952
rect 6917 16943 6975 16949
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 9214 16940 9220 16992
rect 9272 16980 9278 16992
rect 11974 16980 11980 16992
rect 9272 16952 11980 16980
rect 9272 16940 9278 16952
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12342 16940 12348 16992
rect 12400 16980 12406 16992
rect 13372 16980 13400 17020
rect 14277 17017 14289 17020
rect 14323 17017 14335 17051
rect 14277 17011 14335 17017
rect 16301 17051 16359 17057
rect 16301 17017 16313 17051
rect 16347 17048 16359 17051
rect 17310 17048 17316 17060
rect 16347 17020 17316 17048
rect 16347 17017 16359 17020
rect 16301 17011 16359 17017
rect 17310 17008 17316 17020
rect 17368 17008 17374 17060
rect 17405 17051 17463 17057
rect 17405 17017 17417 17051
rect 17451 17048 17463 17051
rect 17678 17048 17684 17060
rect 17451 17020 17684 17048
rect 17451 17017 17463 17020
rect 17405 17011 17463 17017
rect 17678 17008 17684 17020
rect 17736 17008 17742 17060
rect 12400 16952 13400 16980
rect 15657 16983 15715 16989
rect 12400 16940 12406 16952
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 16666 16980 16672 16992
rect 15703 16952 16672 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 17788 16980 17816 17088
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 18012 17088 18981 17116
rect 18012 17076 18018 17088
rect 18969 17085 18981 17088
rect 19015 17085 19027 17119
rect 19150 17116 19156 17128
rect 19111 17088 19156 17116
rect 18969 17079 19027 17085
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 21453 17119 21511 17125
rect 21453 17085 21465 17119
rect 21499 17116 21511 17119
rect 21726 17116 21732 17128
rect 21499 17088 21732 17116
rect 21499 17085 21511 17088
rect 21453 17079 21511 17085
rect 21726 17076 21732 17088
rect 21784 17076 21790 17128
rect 24305 17119 24363 17125
rect 24305 17085 24317 17119
rect 24351 17085 24363 17119
rect 24486 17116 24492 17128
rect 24447 17088 24492 17116
rect 24305 17079 24363 17085
rect 17862 17008 17868 17060
rect 17920 17048 17926 17060
rect 18233 17051 18291 17057
rect 18233 17048 18245 17051
rect 17920 17020 18245 17048
rect 17920 17008 17926 17020
rect 18233 17017 18245 17020
rect 18279 17048 18291 17051
rect 19337 17051 19395 17057
rect 19337 17048 19349 17051
rect 18279 17020 19349 17048
rect 18279 17017 18291 17020
rect 18233 17011 18291 17017
rect 19337 17017 19349 17020
rect 19383 17017 19395 17051
rect 19337 17011 19395 17017
rect 19426 17008 19432 17060
rect 19484 17048 19490 17060
rect 20073 17051 20131 17057
rect 20073 17048 20085 17051
rect 19484 17020 20085 17048
rect 19484 17008 19490 17020
rect 20073 17017 20085 17020
rect 20119 17017 20131 17051
rect 20073 17011 20131 17017
rect 20990 16980 20996 16992
rect 17788 16952 20996 16980
rect 20990 16940 20996 16952
rect 21048 16980 21054 16992
rect 21818 16980 21824 16992
rect 21048 16952 21824 16980
rect 21048 16940 21054 16952
rect 21818 16940 21824 16952
rect 21876 16940 21882 16992
rect 24118 16980 24124 16992
rect 24079 16952 24124 16980
rect 24118 16940 24124 16952
rect 24176 16940 24182 16992
rect 24320 16980 24348 17079
rect 24486 17076 24492 17088
rect 24544 17076 24550 17128
rect 24578 17076 24584 17128
rect 24636 17116 24642 17128
rect 25041 17119 25099 17125
rect 25041 17116 25053 17119
rect 24636 17088 25053 17116
rect 24636 17076 24642 17088
rect 25041 17085 25053 17088
rect 25087 17085 25099 17119
rect 25314 17116 25320 17128
rect 25275 17088 25320 17116
rect 25041 17079 25099 17085
rect 25314 17076 25320 17088
rect 25372 17076 25378 17128
rect 38194 17048 38200 17060
rect 38155 17020 38200 17048
rect 38194 17008 38200 17020
rect 38252 17008 38258 17060
rect 26237 16983 26295 16989
rect 26237 16980 26249 16983
rect 24320 16952 26249 16980
rect 26237 16949 26249 16952
rect 26283 16949 26295 16983
rect 27154 16980 27160 16992
rect 27115 16952 27160 16980
rect 26237 16943 26295 16949
rect 27154 16940 27160 16952
rect 27212 16940 27218 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 1670 16776 1676 16788
rect 1583 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16776 1734 16788
rect 4420 16779 4478 16785
rect 1728 16748 4200 16776
rect 1728 16736 1734 16748
rect 1688 16649 1716 16736
rect 1673 16643 1731 16649
rect 1673 16609 1685 16643
rect 1719 16609 1731 16643
rect 1673 16603 1731 16609
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16640 2007 16643
rect 4062 16640 4068 16652
rect 1995 16612 4068 16640
rect 1995 16609 2007 16612
rect 1949 16603 2007 16609
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4172 16649 4200 16748
rect 4420 16745 4432 16779
rect 4466 16776 4478 16779
rect 4614 16776 4620 16788
rect 4466 16748 4620 16776
rect 4466 16745 4478 16748
rect 4420 16739 4478 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 9122 16776 9128 16788
rect 4948 16748 9128 16776
rect 4948 16736 4954 16748
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 9490 16736 9496 16788
rect 9548 16776 9554 16788
rect 11698 16776 11704 16788
rect 9548 16748 11704 16776
rect 9548 16736 9554 16748
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 11974 16736 11980 16788
rect 12032 16776 12038 16788
rect 15378 16776 15384 16788
rect 12032 16748 15384 16776
rect 12032 16736 12038 16748
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 15528 16748 16313 16776
rect 15528 16736 15534 16748
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16301 16739 16359 16745
rect 17129 16779 17187 16785
rect 17129 16745 17141 16779
rect 17175 16776 17187 16779
rect 17218 16776 17224 16788
rect 17175 16748 17224 16776
rect 17175 16745 17187 16748
rect 17129 16739 17187 16745
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 23477 16779 23535 16785
rect 23477 16745 23489 16779
rect 23523 16776 23535 16779
rect 23566 16776 23572 16788
rect 23523 16748 23572 16776
rect 23523 16745 23535 16748
rect 23477 16739 23535 16745
rect 23566 16736 23572 16748
rect 23624 16736 23630 16788
rect 24118 16736 24124 16788
rect 24176 16776 24182 16788
rect 24578 16776 24584 16788
rect 24176 16748 24584 16776
rect 24176 16736 24182 16748
rect 24578 16736 24584 16748
rect 24636 16736 24642 16788
rect 25130 16736 25136 16788
rect 25188 16776 25194 16788
rect 25685 16779 25743 16785
rect 25685 16776 25697 16779
rect 25188 16748 25697 16776
rect 25188 16736 25194 16748
rect 25685 16745 25697 16748
rect 25731 16745 25743 16779
rect 25685 16739 25743 16745
rect 7006 16668 7012 16720
rect 7064 16708 7070 16720
rect 8938 16708 8944 16720
rect 7064 16680 8944 16708
rect 7064 16668 7070 16680
rect 8938 16668 8944 16680
rect 8996 16668 9002 16720
rect 9140 16708 9168 16736
rect 9140 16680 9444 16708
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4798 16640 4804 16652
rect 4203 16612 4804 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 9125 16643 9183 16649
rect 9125 16609 9137 16643
rect 9171 16640 9183 16643
rect 9306 16640 9312 16652
rect 9171 16612 9312 16640
rect 9171 16609 9183 16612
rect 9125 16603 9183 16609
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 9416 16640 9444 16680
rect 13998 16668 14004 16720
rect 14056 16708 14062 16720
rect 14366 16708 14372 16720
rect 14056 16680 14372 16708
rect 14056 16668 14062 16680
rect 14366 16668 14372 16680
rect 14424 16668 14430 16720
rect 16390 16708 16396 16720
rect 14936 16680 16396 16708
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 9416 16612 10609 16640
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10870 16640 10876 16652
rect 10831 16612 10876 16640
rect 10597 16603 10655 16609
rect 10870 16600 10876 16612
rect 10928 16640 10934 16652
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 10928 16612 11345 16640
rect 10928 16600 10934 16612
rect 11333 16609 11345 16612
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 11606 16600 11612 16652
rect 11664 16640 11670 16652
rect 14936 16640 14964 16680
rect 16390 16668 16396 16680
rect 16448 16668 16454 16720
rect 21634 16708 21640 16720
rect 18248 16680 21640 16708
rect 18248 16649 18276 16680
rect 21634 16668 21640 16680
rect 21692 16668 21698 16720
rect 34238 16708 34244 16720
rect 22940 16680 34244 16708
rect 18049 16643 18107 16649
rect 18049 16640 18061 16643
rect 11664 16612 14964 16640
rect 15028 16612 18061 16640
rect 11664 16600 11670 16612
rect 6822 16572 6828 16584
rect 6783 16544 6828 16572
rect 6822 16532 6828 16544
rect 6880 16532 6886 16584
rect 8846 16532 8852 16584
rect 8904 16572 8910 16584
rect 9214 16572 9220 16584
rect 8904 16544 9220 16572
rect 8904 16532 8910 16544
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 9490 16532 9496 16584
rect 9548 16532 9554 16584
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16572 13599 16575
rect 14182 16572 14188 16584
rect 13587 16544 14188 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 14182 16532 14188 16544
rect 14240 16532 14246 16584
rect 14461 16575 14519 16581
rect 14461 16541 14473 16575
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16572 14611 16575
rect 15028 16572 15056 16612
rect 18049 16609 18061 16612
rect 18095 16609 18107 16643
rect 18049 16603 18107 16609
rect 18233 16643 18291 16649
rect 18233 16609 18245 16643
rect 18279 16609 18291 16643
rect 18233 16603 18291 16609
rect 18690 16600 18696 16652
rect 18748 16640 18754 16652
rect 18748 16612 18920 16640
rect 18748 16600 18754 16612
rect 14599 16544 15056 16572
rect 15841 16575 15899 16581
rect 14599 16541 14611 16544
rect 14553 16535 14611 16541
rect 15841 16541 15853 16575
rect 15887 16572 15899 16575
rect 15930 16572 15936 16584
rect 15887 16544 15936 16572
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 3602 16504 3608 16516
rect 3174 16476 3608 16504
rect 3602 16464 3608 16476
rect 3660 16464 3666 16516
rect 4522 16504 4528 16516
rect 3988 16476 4528 16504
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3384 16408 3433 16436
rect 3384 16396 3390 16408
rect 3421 16405 3433 16408
rect 3467 16436 3479 16439
rect 3988 16436 4016 16476
rect 4522 16464 4528 16476
rect 4580 16464 4586 16516
rect 5902 16504 5908 16516
rect 5658 16476 5908 16504
rect 5902 16464 5908 16476
rect 5960 16464 5966 16516
rect 6181 16507 6239 16513
rect 6181 16473 6193 16507
rect 6227 16504 6239 16507
rect 10502 16504 10508 16516
rect 6227 16476 9260 16504
rect 6227 16473 6239 16476
rect 6181 16467 6239 16473
rect 3467 16408 4016 16436
rect 3467 16405 3479 16408
rect 3421 16399 3479 16405
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 6196 16436 6224 16467
rect 4120 16408 6224 16436
rect 8113 16439 8171 16445
rect 4120 16396 4126 16408
rect 8113 16405 8125 16439
rect 8159 16436 8171 16439
rect 8202 16436 8208 16448
rect 8159 16408 8208 16436
rect 8159 16405 8171 16408
rect 8113 16399 8171 16405
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 9232 16436 9260 16476
rect 10244 16476 10508 16504
rect 10244 16436 10272 16476
rect 10502 16464 10508 16476
rect 10560 16464 10566 16516
rect 11606 16504 11612 16516
rect 11567 16476 11612 16504
rect 11606 16464 11612 16476
rect 11664 16464 11670 16516
rect 12618 16464 12624 16516
rect 12676 16464 12682 16516
rect 14476 16504 14504 16535
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 16482 16572 16488 16584
rect 16443 16544 16488 16572
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16592 16544 16957 16572
rect 15194 16504 15200 16516
rect 13004 16476 14504 16504
rect 15155 16476 15200 16504
rect 9232 16408 10272 16436
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 13004 16436 13032 16476
rect 10928 16408 13032 16436
rect 10928 16396 10934 16408
rect 13078 16396 13084 16448
rect 13136 16436 13142 16448
rect 13725 16439 13783 16445
rect 13136 16408 13181 16436
rect 13136 16396 13142 16408
rect 13725 16405 13737 16439
rect 13771 16436 13783 16439
rect 13814 16436 13820 16448
rect 13771 16408 13820 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 14476 16436 14504 16476
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 15289 16507 15347 16513
rect 15289 16473 15301 16507
rect 15335 16504 15347 16507
rect 15378 16504 15384 16516
rect 15335 16476 15384 16504
rect 15335 16473 15347 16476
rect 15289 16467 15347 16473
rect 15378 16464 15384 16476
rect 15436 16464 15442 16516
rect 16592 16436 16620 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 18782 16572 18788 16584
rect 18743 16544 18788 16572
rect 16945 16535 17003 16541
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 18892 16581 18920 16612
rect 18966 16600 18972 16652
rect 19024 16640 19030 16652
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 19024 16612 19993 16640
rect 19024 16600 19030 16612
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 22646 16640 22652 16652
rect 20211 16612 22652 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 22940 16649 22968 16680
rect 34238 16668 34244 16680
rect 34296 16668 34302 16720
rect 22741 16643 22799 16649
rect 22741 16609 22753 16643
rect 22787 16640 22799 16643
rect 22925 16643 22983 16649
rect 22787 16612 22876 16640
rect 22787 16609 22799 16612
rect 22741 16603 22799 16609
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16541 18935 16575
rect 21450 16572 21456 16584
rect 21411 16544 21456 16572
rect 18877 16535 18935 16541
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 21542 16532 21548 16584
rect 21600 16572 21606 16584
rect 22848 16572 22876 16612
rect 22925 16609 22937 16643
rect 22971 16609 22983 16643
rect 23750 16640 23756 16652
rect 22925 16603 22983 16609
rect 23032 16612 23756 16640
rect 23032 16572 23060 16612
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 23842 16600 23848 16652
rect 23900 16600 23906 16652
rect 25225 16643 25283 16649
rect 25225 16609 25237 16643
rect 25271 16640 25283 16643
rect 25498 16640 25504 16652
rect 25271 16612 25504 16640
rect 25271 16609 25283 16612
rect 25225 16603 25283 16609
rect 25498 16600 25504 16612
rect 25556 16600 25562 16652
rect 38102 16640 38108 16652
rect 35084 16612 38108 16640
rect 21600 16544 21645 16572
rect 22848 16544 23060 16572
rect 23385 16575 23443 16581
rect 21600 16532 21606 16544
rect 23385 16541 23397 16575
rect 23431 16572 23443 16575
rect 23860 16572 23888 16600
rect 25038 16572 25044 16584
rect 23431 16544 23888 16572
rect 24999 16544 25044 16572
rect 23431 16541 23443 16544
rect 23385 16535 23443 16541
rect 17589 16507 17647 16513
rect 17589 16473 17601 16507
rect 17635 16504 17647 16507
rect 18230 16504 18236 16516
rect 17635 16476 18236 16504
rect 17635 16473 17647 16476
rect 17589 16467 17647 16473
rect 18230 16464 18236 16476
rect 18288 16464 18294 16516
rect 18322 16464 18328 16516
rect 18380 16504 18386 16516
rect 22002 16504 22008 16516
rect 18380 16476 22008 16504
rect 18380 16464 18386 16476
rect 22002 16464 22008 16476
rect 22060 16504 22066 16516
rect 23400 16504 23428 16535
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 25869 16575 25927 16581
rect 25869 16541 25881 16575
rect 25915 16572 25927 16575
rect 27154 16572 27160 16584
rect 25915 16544 27160 16572
rect 25915 16541 25927 16544
rect 25869 16535 25927 16541
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 34790 16532 34796 16584
rect 34848 16572 34854 16584
rect 35084 16581 35112 16612
rect 38102 16600 38108 16612
rect 38160 16600 38166 16652
rect 34977 16575 35035 16581
rect 34977 16572 34989 16575
rect 34848 16544 34989 16572
rect 34848 16532 34854 16544
rect 34977 16541 34989 16544
rect 35023 16541 35035 16575
rect 34977 16535 35035 16541
rect 35069 16575 35127 16581
rect 35069 16541 35081 16575
rect 35115 16574 35127 16575
rect 35115 16546 35149 16574
rect 35115 16541 35127 16546
rect 35069 16535 35127 16541
rect 22060 16476 23428 16504
rect 22060 16464 22066 16476
rect 14476 16408 16620 16436
rect 16942 16396 16948 16448
rect 17000 16436 17006 16448
rect 18874 16436 18880 16448
rect 17000 16408 18880 16436
rect 17000 16396 17006 16408
rect 18874 16396 18880 16408
rect 18932 16396 18938 16448
rect 20622 16436 20628 16448
rect 20583 16408 20628 16436
rect 20622 16396 20628 16408
rect 20680 16396 20686 16448
rect 22281 16439 22339 16445
rect 22281 16405 22293 16439
rect 22327 16436 22339 16439
rect 22646 16436 22652 16448
rect 22327 16408 22652 16436
rect 22327 16405 22339 16408
rect 22281 16399 22339 16405
rect 22646 16396 22652 16408
rect 22704 16396 22710 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 1673 16235 1731 16241
rect 1673 16232 1685 16235
rect 1636 16204 1685 16232
rect 1636 16192 1642 16204
rect 1673 16201 1685 16204
rect 1719 16201 1731 16235
rect 1673 16195 1731 16201
rect 3878 16192 3884 16244
rect 3936 16232 3942 16244
rect 3936 16204 6040 16232
rect 3936 16192 3942 16204
rect 5074 16164 5080 16176
rect 4370 16136 5080 16164
rect 5074 16124 5080 16136
rect 5132 16124 5138 16176
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 1946 16096 1952 16108
rect 1903 16068 1952 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 1946 16056 1952 16068
rect 2004 16056 2010 16108
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 6012 16105 6040 16204
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 12989 16235 13047 16241
rect 12989 16232 13001 16235
rect 6880 16204 13001 16232
rect 6880 16192 6886 16204
rect 12989 16201 13001 16204
rect 13035 16201 13047 16235
rect 12989 16195 13047 16201
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 22646 16232 22652 16244
rect 13780 16204 22094 16232
rect 22607 16204 22652 16232
rect 13780 16192 13786 16204
rect 7834 16164 7840 16176
rect 6656 16136 7840 16164
rect 5997 16099 6055 16105
rect 4580 16068 5948 16096
rect 4580 16056 4586 16068
rect 2866 16028 2872 16040
rect 2827 16000 2872 16028
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 3145 16031 3203 16037
rect 3145 15997 3157 16031
rect 3191 16028 3203 16031
rect 3234 16028 3240 16040
rect 3191 16000 3240 16028
rect 3191 15997 3203 16000
rect 3145 15991 3203 15997
rect 3234 15988 3240 16000
rect 3292 16028 3298 16040
rect 4890 16028 4896 16040
rect 3292 16000 4752 16028
rect 4851 16000 4896 16028
rect 3292 15988 3298 16000
rect 4724 15960 4752 16000
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 5920 16028 5948 16068
rect 5997 16065 6009 16099
rect 6043 16065 6055 16099
rect 5997 16059 6055 16065
rect 6546 16028 6552 16040
rect 5920 16000 6552 16028
rect 6546 15988 6552 16000
rect 6604 15988 6610 16040
rect 6656 15960 6684 16136
rect 7834 16124 7840 16136
rect 7892 16124 7898 16176
rect 8754 16124 8760 16176
rect 8812 16124 8818 16176
rect 9766 16124 9772 16176
rect 9824 16164 9830 16176
rect 10137 16167 10195 16173
rect 10137 16164 10149 16167
rect 9824 16136 10149 16164
rect 9824 16124 9830 16136
rect 10137 16133 10149 16136
rect 10183 16133 10195 16167
rect 10137 16127 10195 16133
rect 10226 16124 10232 16176
rect 10284 16164 10290 16176
rect 11149 16167 11207 16173
rect 10284 16136 10329 16164
rect 10284 16124 10290 16136
rect 11149 16133 11161 16167
rect 11195 16164 11207 16167
rect 11195 16136 15240 16164
rect 11195 16133 11207 16136
rect 11149 16127 11207 16133
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 4724 15932 6684 15960
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 5813 15895 5871 15901
rect 5813 15892 5825 15895
rect 2372 15864 5825 15892
rect 2372 15852 2378 15864
rect 5813 15861 5825 15864
rect 5859 15861 5871 15895
rect 6748 15892 6776 16059
rect 9122 16056 9128 16108
rect 9180 16096 9186 16108
rect 11698 16096 11704 16108
rect 9180 16068 9996 16096
rect 11659 16068 11704 16096
rect 9180 16056 9186 16068
rect 7374 15988 7380 16040
rect 7432 16028 7438 16040
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 7432 16000 7481 16028
rect 7432 15988 7438 16000
rect 7469 15997 7481 16000
rect 7515 15997 7527 16031
rect 7742 16028 7748 16040
rect 7703 16000 7748 16028
rect 7469 15991 7527 15997
rect 6914 15960 6920 15972
rect 6875 15932 6920 15960
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7098 15892 7104 15904
rect 6748 15864 7104 15892
rect 5813 15855 5871 15861
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7484 15892 7512 15991
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 8110 15988 8116 16040
rect 8168 16028 8174 16040
rect 9674 16028 9680 16040
rect 8168 16000 9680 16028
rect 8168 15988 8174 16000
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 9968 16028 9996 16068
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 13722 16028 13728 16040
rect 9968 16000 13728 16028
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 13906 16028 13912 16040
rect 13867 16000 13912 16028
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 13998 15988 14004 16040
rect 14056 16028 14062 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 14056 16000 14105 16028
rect 14056 15988 14062 16000
rect 14093 15997 14105 16000
rect 14139 15997 14151 16031
rect 15212 16028 15240 16136
rect 15930 16124 15936 16176
rect 15988 16164 15994 16176
rect 16117 16167 16175 16173
rect 16117 16164 16129 16167
rect 15988 16136 16129 16164
rect 15988 16124 15994 16136
rect 16117 16133 16129 16136
rect 16163 16133 16175 16167
rect 16117 16127 16175 16133
rect 16390 16124 16396 16176
rect 16448 16164 16454 16176
rect 19981 16167 20039 16173
rect 16448 16136 19656 16164
rect 16448 16124 16454 16136
rect 16666 16056 16672 16108
rect 16724 16096 16730 16108
rect 17129 16099 17187 16105
rect 17129 16096 17141 16099
rect 16724 16068 17141 16096
rect 16724 16056 16730 16068
rect 17129 16065 17141 16068
rect 17175 16065 17187 16099
rect 17129 16059 17187 16065
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16096 17279 16099
rect 19521 16099 19579 16105
rect 19521 16096 19533 16099
rect 17267 16068 19533 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 19521 16065 19533 16068
rect 19567 16065 19579 16099
rect 19521 16059 19579 16065
rect 15933 16031 15991 16037
rect 15933 16028 15945 16031
rect 15212 16000 15945 16028
rect 14093 15991 14151 15997
rect 15933 15997 15945 16000
rect 15979 16028 15991 16031
rect 16022 16028 16028 16040
rect 15979 16000 16028 16028
rect 15979 15997 15991 16000
rect 15933 15991 15991 15997
rect 16022 15988 16028 16000
rect 16080 15988 16086 16040
rect 16206 16028 16212 16040
rect 16167 16000 16212 16028
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 16574 15988 16580 16040
rect 16632 16028 16638 16040
rect 17678 16028 17684 16040
rect 16632 16000 17684 16028
rect 16632 15988 16638 16000
rect 17678 15988 17684 16000
rect 17736 16028 17742 16040
rect 17773 16031 17831 16037
rect 17773 16028 17785 16031
rect 17736 16000 17785 16028
rect 17736 15988 17742 16000
rect 17773 15997 17785 16000
rect 17819 15997 17831 16031
rect 17773 15991 17831 15997
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 15997 18015 16031
rect 17957 15991 18015 15997
rect 10318 15920 10324 15972
rect 10376 15960 10382 15972
rect 10870 15960 10876 15972
rect 10376 15932 10876 15960
rect 10376 15920 10382 15932
rect 10870 15920 10876 15932
rect 10928 15920 10934 15972
rect 11974 15920 11980 15972
rect 12032 15960 12038 15972
rect 12032 15932 14504 15960
rect 12032 15920 12038 15932
rect 8202 15892 8208 15904
rect 7484 15864 8208 15892
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 9122 15852 9128 15904
rect 9180 15892 9186 15904
rect 9217 15895 9275 15901
rect 9217 15892 9229 15895
rect 9180 15864 9229 15892
rect 9180 15852 9186 15864
rect 9217 15861 9229 15864
rect 9263 15861 9275 15895
rect 9217 15855 9275 15861
rect 9398 15852 9404 15904
rect 9456 15892 9462 15904
rect 13538 15892 13544 15904
rect 9456 15864 13544 15892
rect 9456 15852 9462 15864
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 14274 15892 14280 15904
rect 14235 15864 14280 15892
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 14476 15892 14504 15932
rect 14550 15920 14556 15972
rect 14608 15960 14614 15972
rect 17972 15960 18000 15991
rect 18414 15988 18420 16040
rect 18472 16028 18478 16040
rect 19337 16031 19395 16037
rect 19337 16028 19349 16031
rect 18472 16000 19349 16028
rect 18472 15988 18478 16000
rect 19337 15997 19349 16000
rect 19383 15997 19395 16031
rect 19628 16028 19656 16136
rect 19981 16133 19993 16167
rect 20027 16164 20039 16167
rect 20622 16164 20628 16176
rect 20027 16136 20628 16164
rect 20027 16133 20039 16136
rect 19981 16127 20039 16133
rect 20622 16124 20628 16136
rect 20680 16164 20686 16176
rect 20809 16167 20867 16173
rect 20809 16164 20821 16167
rect 20680 16136 20821 16164
rect 20680 16124 20686 16136
rect 20809 16133 20821 16136
rect 20855 16133 20867 16167
rect 20809 16127 20867 16133
rect 20898 16124 20904 16176
rect 20956 16164 20962 16176
rect 22066 16164 22094 16204
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 22738 16192 22744 16244
rect 22796 16232 22802 16244
rect 23109 16235 23167 16241
rect 23109 16232 23121 16235
rect 22796 16204 23121 16232
rect 22796 16192 22802 16204
rect 23109 16201 23121 16204
rect 23155 16201 23167 16235
rect 23750 16232 23756 16244
rect 23711 16204 23756 16232
rect 23109 16195 23167 16201
rect 23750 16192 23756 16204
rect 23808 16192 23814 16244
rect 25038 16232 25044 16244
rect 24999 16204 25044 16232
rect 25038 16192 25044 16204
rect 25096 16192 25102 16244
rect 20956 16136 21001 16164
rect 22066 16136 24624 16164
rect 20956 16124 20962 16136
rect 24596 16108 24624 16136
rect 21542 16056 21548 16108
rect 21600 16096 21606 16108
rect 23293 16099 23351 16105
rect 23293 16096 23305 16099
rect 21600 16068 23305 16096
rect 21600 16056 21606 16068
rect 23293 16065 23305 16068
rect 23339 16065 23351 16099
rect 23293 16059 23351 16065
rect 23937 16099 23995 16105
rect 23937 16065 23949 16099
rect 23983 16096 23995 16099
rect 23983 16068 24440 16096
rect 23983 16065 23995 16068
rect 23937 16059 23995 16065
rect 19628 16000 21588 16028
rect 19337 15991 19395 15997
rect 18138 15960 18144 15972
rect 14608 15932 18000 15960
rect 18099 15932 18144 15960
rect 14608 15920 14614 15932
rect 18138 15920 18144 15932
rect 18196 15920 18202 15972
rect 21361 15963 21419 15969
rect 21361 15929 21373 15963
rect 21407 15960 21419 15963
rect 21450 15960 21456 15972
rect 21407 15932 21456 15960
rect 21407 15929 21419 15932
rect 21361 15923 21419 15929
rect 21450 15920 21456 15932
rect 21508 15920 21514 15972
rect 21560 15960 21588 16000
rect 21910 15988 21916 16040
rect 21968 16028 21974 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 21968 16000 22017 16028
rect 21968 15988 21974 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22186 16028 22192 16040
rect 22147 16000 22192 16028
rect 22005 15991 22063 15997
rect 22186 15988 22192 16000
rect 22244 15988 22250 16040
rect 22462 15988 22468 16040
rect 22520 16028 22526 16040
rect 24302 16028 24308 16040
rect 22520 16000 24308 16028
rect 22520 15988 22526 16000
rect 24302 15988 24308 16000
rect 24360 15988 24366 16040
rect 23750 15960 23756 15972
rect 21560 15932 23756 15960
rect 23750 15920 23756 15932
rect 23808 15920 23814 15972
rect 24412 15969 24440 16068
rect 24578 16056 24584 16108
rect 24636 16096 24642 16108
rect 25225 16099 25283 16105
rect 24636 16068 24729 16096
rect 24636 16056 24642 16068
rect 25225 16065 25237 16099
rect 25271 16096 25283 16099
rect 25869 16099 25927 16105
rect 25271 16068 25728 16096
rect 25271 16065 25283 16068
rect 25225 16059 25283 16065
rect 25700 15969 25728 16068
rect 25869 16065 25881 16099
rect 25915 16096 25927 16099
rect 26142 16096 26148 16108
rect 25915 16068 26148 16096
rect 25915 16065 25927 16068
rect 25869 16059 25927 16065
rect 24397 15963 24455 15969
rect 24397 15929 24409 15963
rect 24443 15929 24455 15963
rect 24397 15923 24455 15929
rect 25685 15963 25743 15969
rect 25685 15929 25697 15963
rect 25731 15929 25743 15963
rect 25685 15923 25743 15929
rect 16482 15892 16488 15904
rect 14476 15864 16488 15892
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 25884 15892 25912 16059
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 22612 15864 25912 15892
rect 22612 15852 22618 15864
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 3292 15660 3341 15688
rect 3292 15648 3298 15660
rect 3329 15657 3341 15660
rect 3375 15657 3387 15691
rect 3329 15651 3387 15657
rect 8573 15691 8631 15697
rect 8573 15657 8585 15691
rect 8619 15688 8631 15691
rect 11606 15688 11612 15700
rect 8619 15660 11612 15688
rect 8619 15657 8631 15660
rect 8573 15651 8631 15657
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 13633 15691 13691 15697
rect 13633 15657 13645 15691
rect 13679 15688 13691 15691
rect 14274 15688 14280 15700
rect 13679 15660 14280 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 14550 15688 14556 15700
rect 14511 15660 14556 15688
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 14642 15648 14648 15700
rect 14700 15688 14706 15700
rect 16574 15688 16580 15700
rect 14700 15660 16580 15688
rect 14700 15648 14706 15660
rect 16574 15648 16580 15660
rect 16632 15648 16638 15700
rect 16945 15691 17003 15697
rect 16945 15657 16957 15691
rect 16991 15688 17003 15691
rect 18322 15688 18328 15700
rect 16991 15660 18328 15688
rect 16991 15657 17003 15660
rect 16945 15651 17003 15657
rect 18322 15648 18328 15660
rect 18380 15648 18386 15700
rect 20070 15688 20076 15700
rect 19983 15660 20076 15688
rect 20070 15648 20076 15660
rect 20128 15688 20134 15700
rect 20530 15688 20536 15700
rect 20128 15660 20536 15688
rect 20128 15648 20134 15660
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 24673 15691 24731 15697
rect 24673 15688 24685 15691
rect 22244 15660 24685 15688
rect 22244 15648 22250 15660
rect 24673 15657 24685 15660
rect 24719 15657 24731 15691
rect 38102 15688 38108 15700
rect 38063 15660 38108 15688
rect 24673 15651 24731 15657
rect 38102 15648 38108 15660
rect 38160 15648 38166 15700
rect 4065 15623 4123 15629
rect 4065 15589 4077 15623
rect 4111 15620 4123 15623
rect 4111 15592 5396 15620
rect 4111 15589 4123 15592
rect 4065 15583 4123 15589
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15552 1639 15555
rect 2866 15552 2872 15564
rect 1627 15524 2872 15552
rect 1627 15521 1639 15524
rect 1581 15515 1639 15521
rect 2866 15512 2872 15524
rect 2924 15552 2930 15564
rect 3602 15552 3608 15564
rect 2924 15524 3608 15552
rect 2924 15512 2930 15524
rect 3602 15512 3608 15524
rect 3660 15552 3666 15564
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 3660 15524 5273 15552
rect 3660 15512 3666 15524
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 5368 15552 5396 15592
rect 6730 15580 6736 15632
rect 6788 15620 6794 15632
rect 8938 15620 8944 15632
rect 6788 15592 8944 15620
rect 6788 15580 6794 15592
rect 8938 15580 8944 15592
rect 8996 15580 9002 15632
rect 10502 15580 10508 15632
rect 10560 15620 10566 15632
rect 22554 15620 22560 15632
rect 10560 15592 22560 15620
rect 10560 15580 10566 15592
rect 22554 15580 22560 15592
rect 22612 15580 22618 15632
rect 27430 15620 27436 15632
rect 22848 15592 27436 15620
rect 22848 15564 22876 15592
rect 27430 15580 27436 15592
rect 27488 15580 27494 15632
rect 12342 15552 12348 15564
rect 5368 15524 11008 15552
rect 12303 15524 12348 15552
rect 5261 15515 5319 15521
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15484 4675 15487
rect 4890 15484 4896 15496
rect 4663 15456 4896 15484
rect 4663 15453 4675 15456
rect 4617 15447 4675 15453
rect 1857 15419 1915 15425
rect 1857 15385 1869 15419
rect 1903 15385 1915 15419
rect 3878 15416 3884 15428
rect 3082 15388 3884 15416
rect 1857 15379 1915 15385
rect 1872 15348 1900 15379
rect 3878 15376 3884 15388
rect 3936 15376 3942 15428
rect 4172 15416 4200 15447
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 6914 15444 6920 15496
rect 6972 15484 6978 15496
rect 6972 15456 7420 15484
rect 6972 15444 6978 15456
rect 5258 15416 5264 15428
rect 4172 15388 5264 15416
rect 5258 15376 5264 15388
rect 5316 15376 5322 15428
rect 5534 15416 5540 15428
rect 5495 15388 5540 15416
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 5994 15376 6000 15428
rect 6052 15376 6058 15428
rect 7282 15416 7288 15428
rect 7243 15388 7288 15416
rect 7282 15376 7288 15388
rect 7340 15376 7346 15428
rect 7392 15416 7420 15456
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 7929 15487 7987 15493
rect 7929 15484 7941 15487
rect 7524 15456 7941 15484
rect 7524 15444 7530 15456
rect 7929 15453 7941 15456
rect 7975 15453 7987 15487
rect 7929 15447 7987 15453
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 8128 15416 8156 15447
rect 8846 15444 8852 15496
rect 8904 15484 8910 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8904 15456 9137 15484
rect 8904 15444 8910 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 7392 15388 8156 15416
rect 8938 15376 8944 15428
rect 8996 15416 9002 15428
rect 9401 15419 9459 15425
rect 9401 15416 9413 15419
rect 8996 15388 9413 15416
rect 8996 15376 9002 15388
rect 9401 15385 9413 15388
rect 9447 15385 9459 15419
rect 9401 15379 9459 15385
rect 10134 15376 10140 15428
rect 10192 15376 10198 15428
rect 4062 15348 4068 15360
rect 1872 15320 4068 15348
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 4801 15351 4859 15357
rect 4801 15317 4813 15351
rect 4847 15348 4859 15351
rect 8386 15348 8392 15360
rect 4847 15320 8392 15348
rect 4847 15317 4859 15320
rect 4801 15311 4859 15317
rect 8386 15308 8392 15320
rect 8444 15308 8450 15360
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 9674 15348 9680 15360
rect 8536 15320 9680 15348
rect 8536 15308 8542 15320
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 10410 15308 10416 15360
rect 10468 15348 10474 15360
rect 10873 15351 10931 15357
rect 10873 15348 10885 15351
rect 10468 15320 10885 15348
rect 10468 15308 10474 15320
rect 10873 15317 10885 15320
rect 10919 15317 10931 15351
rect 10980 15348 11008 15524
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 12989 15555 13047 15561
rect 12989 15521 13001 15555
rect 13035 15552 13047 15555
rect 13814 15552 13820 15564
rect 13035 15524 13820 15552
rect 13035 15521 13047 15524
rect 12989 15515 13047 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 14182 15512 14188 15564
rect 14240 15552 14246 15564
rect 15470 15552 15476 15564
rect 14240 15524 15476 15552
rect 14240 15512 14246 15524
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 15749 15555 15807 15561
rect 15749 15521 15761 15555
rect 15795 15552 15807 15555
rect 16390 15552 16396 15564
rect 15795 15524 16396 15552
rect 15795 15521 15807 15524
rect 15749 15515 15807 15521
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 18877 15555 18935 15561
rect 18877 15521 18889 15555
rect 18923 15552 18935 15555
rect 18966 15552 18972 15564
rect 18923 15524 18972 15552
rect 18923 15521 18935 15524
rect 18877 15515 18935 15521
rect 18966 15512 18972 15524
rect 19024 15512 19030 15564
rect 21174 15552 21180 15564
rect 21135 15524 21180 15552
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 21450 15552 21456 15564
rect 21411 15524 21456 15552
rect 21450 15512 21456 15524
rect 21508 15552 21514 15564
rect 22664 15552 22876 15564
rect 23106 15552 23112 15564
rect 21508 15536 22876 15552
rect 21508 15524 22692 15536
rect 23067 15524 23112 15552
rect 21508 15512 21514 15524
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15453 13231 15487
rect 13173 15447 13231 15453
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15453 14427 15487
rect 16758 15484 16764 15496
rect 16719 15456 16764 15484
rect 14369 15447 14427 15453
rect 11514 15376 11520 15428
rect 11572 15416 11578 15428
rect 11701 15419 11759 15425
rect 11701 15416 11713 15419
rect 11572 15388 11713 15416
rect 11572 15376 11578 15388
rect 11701 15385 11713 15388
rect 11747 15385 11759 15419
rect 11701 15379 11759 15385
rect 12066 15376 12072 15428
rect 12124 15416 12130 15428
rect 12253 15419 12311 15425
rect 12253 15416 12265 15419
rect 12124 15388 12265 15416
rect 12124 15376 12130 15388
rect 12253 15385 12265 15388
rect 12299 15385 12311 15419
rect 12253 15379 12311 15385
rect 13188 15348 13216 15447
rect 10980 15320 13216 15348
rect 14384 15348 14412 15447
rect 16758 15444 16764 15456
rect 16816 15444 16822 15496
rect 20254 15484 20260 15496
rect 20215 15456 20260 15484
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15453 20499 15487
rect 24026 15484 24032 15496
rect 23987 15456 24032 15484
rect 20441 15447 20499 15453
rect 15102 15416 15108 15428
rect 15063 15388 15108 15416
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 15197 15419 15255 15425
rect 15197 15385 15209 15419
rect 15243 15416 15255 15419
rect 15286 15416 15292 15428
rect 15243 15388 15292 15416
rect 15243 15385 15255 15388
rect 15197 15379 15255 15385
rect 15286 15376 15292 15388
rect 15344 15376 15350 15428
rect 17402 15416 17408 15428
rect 17363 15388 17408 15416
rect 17402 15376 17408 15388
rect 17460 15376 17466 15428
rect 17957 15419 18015 15425
rect 17957 15385 17969 15419
rect 18003 15385 18015 15419
rect 17957 15379 18015 15385
rect 18049 15419 18107 15425
rect 18049 15385 18061 15419
rect 18095 15416 18107 15419
rect 20346 15416 20352 15428
rect 18095 15388 20352 15416
rect 18095 15385 18107 15388
rect 18049 15379 18107 15385
rect 17770 15348 17776 15360
rect 14384 15320 17776 15348
rect 10873 15311 10931 15317
rect 17770 15308 17776 15320
rect 17828 15308 17834 15360
rect 17972 15348 18000 15379
rect 20346 15376 20352 15388
rect 20404 15376 20410 15428
rect 18138 15348 18144 15360
rect 17972 15320 18144 15348
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 20456 15348 20484 15447
rect 24026 15444 24032 15456
rect 24084 15444 24090 15496
rect 24578 15484 24584 15496
rect 24539 15456 24584 15484
rect 24578 15444 24584 15456
rect 24636 15444 24642 15496
rect 38286 15484 38292 15496
rect 38247 15456 38292 15484
rect 38286 15444 38292 15456
rect 38344 15444 38350 15496
rect 21266 15376 21272 15428
rect 21324 15416 21330 15428
rect 22738 15416 22744 15428
rect 21324 15388 21369 15416
rect 22699 15388 22744 15416
rect 21324 15376 21330 15388
rect 22738 15376 22744 15388
rect 22796 15376 22802 15428
rect 22833 15419 22891 15425
rect 22833 15385 22845 15419
rect 22879 15416 22891 15419
rect 22879 15388 23060 15416
rect 22879 15385 22891 15388
rect 22833 15379 22891 15385
rect 22462 15348 22468 15360
rect 20456 15320 22468 15348
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 23032 15348 23060 15388
rect 23658 15348 23664 15360
rect 23032 15320 23664 15348
rect 23658 15308 23664 15320
rect 23716 15308 23722 15360
rect 23842 15348 23848 15360
rect 23803 15320 23848 15348
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 1765 15147 1823 15153
rect 1765 15113 1777 15147
rect 1811 15144 1823 15147
rect 2038 15144 2044 15156
rect 1811 15116 2044 15144
rect 1811 15113 1823 15116
rect 1765 15107 1823 15113
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 3694 15104 3700 15156
rect 3752 15144 3758 15156
rect 11698 15144 11704 15156
rect 3752 15116 11704 15144
rect 3752 15104 3758 15116
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 16758 15144 16764 15156
rect 12360 15116 16764 15144
rect 3786 15036 3792 15088
rect 3844 15076 3850 15088
rect 3881 15079 3939 15085
rect 3881 15076 3893 15079
rect 3844 15048 3893 15076
rect 3844 15036 3850 15048
rect 3881 15045 3893 15048
rect 3927 15045 3939 15079
rect 3881 15039 3939 15045
rect 4890 15036 4896 15088
rect 4948 15036 4954 15088
rect 6914 15076 6920 15088
rect 5644 15048 6920 15076
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1762 15008 1768 15020
rect 1719 14980 1768 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 2314 15008 2320 15020
rect 2275 14980 2320 15008
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 14977 3019 15011
rect 3602 15008 3608 15020
rect 3563 14980 3608 15008
rect 2961 14971 3019 14977
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 2774 14804 2780 14816
rect 2455 14776 2780 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 2976 14804 3004 14971
rect 3602 14968 3608 14980
rect 3660 14968 3666 15020
rect 5644 15008 5672 15048
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 9030 15036 9036 15088
rect 9088 15076 9094 15088
rect 9125 15079 9183 15085
rect 9125 15076 9137 15079
rect 9088 15048 9137 15076
rect 9088 15036 9094 15048
rect 9125 15045 9137 15048
rect 9171 15045 9183 15079
rect 10962 15076 10968 15088
rect 10350 15048 10968 15076
rect 9125 15039 9183 15045
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 12250 15076 12256 15088
rect 12211 15048 12256 15076
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 12360 15085 12388 15116
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 17221 15147 17279 15153
rect 17221 15113 17233 15147
rect 17267 15144 17279 15147
rect 17586 15144 17592 15156
rect 17267 15116 17592 15144
rect 17267 15113 17279 15116
rect 17221 15107 17279 15113
rect 17586 15104 17592 15116
rect 17644 15104 17650 15156
rect 19705 15147 19763 15153
rect 17880 15116 19656 15144
rect 12345 15079 12403 15085
rect 12345 15045 12357 15079
rect 12391 15045 12403 15079
rect 14182 15076 14188 15088
rect 12345 15039 12403 15045
rect 12820 15048 14188 15076
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 5552 14980 5672 15008
rect 6380 14980 6561 15008
rect 5552 14940 5580 14980
rect 3160 14912 5580 14940
rect 5629 14943 5687 14949
rect 3160 14881 3188 14912
rect 5629 14909 5641 14943
rect 5675 14909 5687 14943
rect 5629 14903 5687 14909
rect 3145 14875 3203 14881
rect 3145 14841 3157 14875
rect 3191 14841 3203 14875
rect 3145 14835 3203 14841
rect 5258 14832 5264 14884
rect 5316 14872 5322 14884
rect 5644 14872 5672 14903
rect 5316 14844 5672 14872
rect 6380 14872 6408 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 7926 14968 7932 15020
rect 7984 14968 7990 15020
rect 10502 14968 10508 15020
rect 10560 15008 10566 15020
rect 10560 14980 11192 15008
rect 10560 14968 10566 14980
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6512 14912 6837 14940
rect 6512 14900 6518 14912
rect 6825 14909 6837 14912
rect 6871 14940 6883 14943
rect 7834 14940 7840 14952
rect 6871 14912 7840 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 8846 14940 8852 14952
rect 8220 14912 8852 14940
rect 6380 14844 6684 14872
rect 5316 14832 5322 14844
rect 6270 14804 6276 14816
rect 2976 14776 6276 14804
rect 6270 14764 6276 14776
rect 6328 14764 6334 14816
rect 6656 14804 6684 14844
rect 7374 14804 7380 14816
rect 6656 14776 7380 14804
rect 7374 14764 7380 14776
rect 7432 14804 7438 14816
rect 8220 14804 8248 14912
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 9214 14900 9220 14952
rect 9272 14940 9278 14952
rect 11054 14940 11060 14952
rect 9272 14912 11060 14940
rect 9272 14900 9278 14912
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11164 14940 11192 14980
rect 12820 14940 12848 15048
rect 14182 15036 14188 15048
rect 14240 15036 14246 15088
rect 14274 15036 14280 15088
rect 14332 15076 14338 15088
rect 15657 15079 15715 15085
rect 15657 15076 15669 15079
rect 14332 15048 15669 15076
rect 14332 15036 14338 15048
rect 15657 15045 15669 15048
rect 15703 15045 15715 15079
rect 15657 15039 15715 15045
rect 15749 15079 15807 15085
rect 15749 15045 15761 15079
rect 15795 15076 15807 15079
rect 16942 15076 16948 15088
rect 15795 15048 16948 15076
rect 15795 15045 15807 15048
rect 15749 15039 15807 15045
rect 16942 15036 16948 15048
rect 17000 15036 17006 15088
rect 17880 15076 17908 15116
rect 17052 15048 17908 15076
rect 17957 15079 18015 15085
rect 12986 14968 12992 15020
rect 13044 15008 13050 15020
rect 13044 14980 14964 15008
rect 13044 14968 13050 14980
rect 11164 14912 12848 14940
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 13078 14940 13084 14952
rect 12952 14912 12997 14940
rect 13039 14912 13084 14940
rect 12952 14900 12958 14912
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 13872 14912 14473 14940
rect 13872 14900 13878 14912
rect 14461 14909 14473 14912
rect 14507 14940 14519 14943
rect 14550 14940 14556 14952
rect 14507 14912 14556 14940
rect 14507 14909 14519 14912
rect 14461 14903 14519 14909
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14940 14703 14943
rect 14826 14940 14832 14952
rect 14691 14912 14832 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 14826 14900 14832 14912
rect 14884 14900 14890 14952
rect 14936 14940 14964 14980
rect 16666 14968 16672 15020
rect 16724 15008 16730 15020
rect 17052 15008 17080 15048
rect 17957 15045 17969 15079
rect 18003 15076 18015 15079
rect 18046 15076 18052 15088
rect 18003 15048 18052 15076
rect 18003 15045 18015 15048
rect 17957 15039 18015 15045
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 19628 15076 19656 15116
rect 19705 15113 19717 15147
rect 19751 15144 19763 15147
rect 20070 15144 20076 15156
rect 19751 15116 20076 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 20898 15104 20904 15156
rect 20956 15144 20962 15156
rect 22005 15147 22063 15153
rect 22005 15144 22017 15147
rect 20956 15116 22017 15144
rect 20956 15104 20962 15116
rect 22005 15113 22017 15116
rect 22051 15113 22063 15147
rect 23842 15144 23848 15156
rect 22005 15107 22063 15113
rect 22756 15116 23848 15144
rect 20162 15076 20168 15088
rect 19628 15048 20168 15076
rect 20162 15036 20168 15048
rect 20220 15076 20226 15088
rect 20220 15048 21312 15076
rect 20220 15036 20226 15048
rect 16724 14980 17080 15008
rect 17129 15011 17187 15017
rect 16724 14968 16730 14980
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 20625 15011 20683 15017
rect 20625 14977 20637 15011
rect 20671 15008 20683 15011
rect 21174 15008 21180 15020
rect 20671 14980 21180 15008
rect 20671 14977 20683 14980
rect 20625 14971 20683 14977
rect 17144 14940 17172 14971
rect 21174 14968 21180 14980
rect 21232 14968 21238 15020
rect 21284 15017 21312 15048
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 22189 15011 22247 15017
rect 22189 14977 22201 15011
rect 22235 15008 22247 15011
rect 22756 15008 22784 15116
rect 23842 15104 23848 15116
rect 23900 15104 23906 15156
rect 23293 15079 23351 15085
rect 23293 15045 23305 15079
rect 23339 15076 23351 15079
rect 24578 15076 24584 15088
rect 23339 15048 24584 15076
rect 23339 15045 23351 15048
rect 23293 15039 23351 15045
rect 24578 15036 24584 15048
rect 24636 15036 24642 15088
rect 22235 14980 22784 15008
rect 22235 14977 22247 14980
rect 22189 14971 22247 14977
rect 23566 14968 23572 15020
rect 23624 15008 23630 15020
rect 24121 15011 24179 15017
rect 24121 15008 24133 15011
rect 23624 14980 24133 15008
rect 23624 14968 23630 14980
rect 24121 14977 24133 14980
rect 24167 14977 24179 15011
rect 24762 15008 24768 15020
rect 24723 14980 24768 15008
rect 24121 14971 24179 14977
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 29181 15011 29239 15017
rect 29181 14977 29193 15011
rect 29227 14977 29239 15011
rect 29181 14971 29239 14977
rect 17862 14940 17868 14952
rect 14936 14912 17172 14940
rect 17823 14912 17868 14940
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 18230 14900 18236 14952
rect 18288 14940 18294 14952
rect 19058 14940 19064 14952
rect 18288 14912 19064 14940
rect 18288 14900 18294 14912
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 19245 14943 19303 14949
rect 19245 14909 19257 14943
rect 19291 14909 19303 14943
rect 20806 14940 20812 14952
rect 20767 14912 20812 14940
rect 19245 14903 19303 14909
rect 10226 14832 10232 14884
rect 10284 14872 10290 14884
rect 11514 14872 11520 14884
rect 10284 14844 11520 14872
rect 10284 14832 10290 14844
rect 11514 14832 11520 14844
rect 11572 14872 11578 14884
rect 11793 14875 11851 14881
rect 11793 14872 11805 14875
rect 11572 14844 11805 14872
rect 11572 14832 11578 14844
rect 11793 14841 11805 14844
rect 11839 14841 11851 14875
rect 11793 14835 11851 14841
rect 13354 14832 13360 14884
rect 13412 14872 13418 14884
rect 16209 14875 16267 14881
rect 13412 14844 16160 14872
rect 13412 14832 13418 14844
rect 7432 14776 8248 14804
rect 8297 14807 8355 14813
rect 7432 14764 7438 14776
rect 8297 14773 8309 14807
rect 8343 14804 8355 14807
rect 9858 14804 9864 14816
rect 8343 14776 9864 14804
rect 8343 14773 8355 14776
rect 8297 14767 8355 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10502 14764 10508 14816
rect 10560 14804 10566 14816
rect 10597 14807 10655 14813
rect 10597 14804 10609 14807
rect 10560 14776 10609 14804
rect 10560 14764 10566 14776
rect 10597 14773 10609 14776
rect 10643 14804 10655 14807
rect 11054 14804 11060 14816
rect 10643 14776 11060 14804
rect 10643 14773 10655 14776
rect 10597 14767 10655 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 13541 14807 13599 14813
rect 13541 14773 13553 14807
rect 13587 14804 13599 14807
rect 13722 14804 13728 14816
rect 13587 14776 13728 14804
rect 13587 14773 13599 14776
rect 13541 14767 13599 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 15102 14804 15108 14816
rect 15063 14776 15108 14804
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 16132 14804 16160 14844
rect 16209 14841 16221 14875
rect 16255 14872 16267 14875
rect 18417 14875 18475 14881
rect 18417 14872 18429 14875
rect 16255 14844 18429 14872
rect 16255 14841 16267 14844
rect 16209 14835 16267 14841
rect 18417 14841 18429 14844
rect 18463 14872 18475 14875
rect 18782 14872 18788 14884
rect 18463 14844 18788 14872
rect 18463 14841 18475 14844
rect 18417 14835 18475 14841
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 19260 14872 19288 14903
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 23106 14940 23112 14952
rect 23019 14912 23112 14940
rect 23106 14900 23112 14912
rect 23164 14900 23170 14952
rect 23290 14900 23296 14952
rect 23348 14940 23354 14952
rect 23385 14943 23443 14949
rect 23385 14940 23397 14943
rect 23348 14912 23397 14940
rect 23348 14900 23354 14912
rect 23385 14909 23397 14912
rect 23431 14909 23443 14943
rect 23385 14903 23443 14909
rect 23658 14900 23664 14952
rect 23716 14940 23722 14952
rect 24673 14943 24731 14949
rect 24673 14940 24685 14943
rect 23716 14912 24685 14940
rect 23716 14900 23722 14912
rect 24673 14909 24685 14912
rect 24719 14909 24731 14943
rect 24673 14903 24731 14909
rect 23124 14872 23152 14900
rect 29196 14872 29224 14971
rect 19260 14844 22094 14872
rect 23124 14844 29224 14872
rect 19426 14804 19432 14816
rect 16132 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 19978 14764 19984 14816
rect 20036 14804 20042 14816
rect 20165 14807 20223 14813
rect 20165 14804 20177 14807
rect 20036 14776 20177 14804
rect 20036 14764 20042 14776
rect 20165 14773 20177 14776
rect 20211 14773 20223 14807
rect 20165 14767 20223 14773
rect 21453 14807 21511 14813
rect 21453 14773 21465 14807
rect 21499 14804 21511 14807
rect 21542 14804 21548 14816
rect 21499 14776 21548 14804
rect 21499 14773 21511 14776
rect 21453 14767 21511 14773
rect 21542 14764 21548 14776
rect 21600 14764 21606 14816
rect 22066 14804 22094 14844
rect 23937 14807 23995 14813
rect 23937 14804 23949 14807
rect 22066 14776 23949 14804
rect 23937 14773 23949 14776
rect 23983 14773 23995 14807
rect 29270 14804 29276 14816
rect 29231 14776 29276 14804
rect 23937 14767 23995 14773
rect 29270 14764 29276 14776
rect 29328 14764 29334 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 4430 14600 4436 14612
rect 2832 14572 4436 14600
rect 2832 14560 2838 14572
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 4709 14603 4767 14609
rect 4709 14569 4721 14603
rect 4755 14600 4767 14603
rect 10042 14600 10048 14612
rect 4755 14572 10048 14600
rect 4755 14569 4767 14572
rect 4709 14563 4767 14569
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10870 14600 10876 14612
rect 10831 14572 10876 14600
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 12342 14560 12348 14612
rect 12400 14600 12406 14612
rect 14550 14600 14556 14612
rect 12400 14572 14556 14600
rect 12400 14560 12406 14572
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 15102 14560 15108 14612
rect 15160 14600 15166 14612
rect 16117 14603 16175 14609
rect 16117 14600 16129 14603
rect 15160 14572 16129 14600
rect 15160 14560 15166 14572
rect 16117 14569 16129 14572
rect 16163 14569 16175 14603
rect 16117 14563 16175 14569
rect 17770 14560 17776 14612
rect 17828 14600 17834 14612
rect 18693 14603 18751 14609
rect 18693 14600 18705 14603
rect 17828 14572 18705 14600
rect 17828 14560 17834 14572
rect 18693 14569 18705 14572
rect 18739 14569 18751 14603
rect 18693 14563 18751 14569
rect 19521 14603 19579 14609
rect 19521 14569 19533 14603
rect 19567 14600 19579 14603
rect 20254 14600 20260 14612
rect 19567 14572 20260 14600
rect 19567 14569 19579 14572
rect 19521 14563 19579 14569
rect 20254 14560 20260 14572
rect 20312 14560 20318 14612
rect 20349 14603 20407 14609
rect 20349 14569 20361 14603
rect 20395 14600 20407 14603
rect 20438 14600 20444 14612
rect 20395 14572 20444 14600
rect 20395 14569 20407 14572
rect 20349 14563 20407 14569
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 21266 14560 21272 14612
rect 21324 14600 21330 14612
rect 21361 14603 21419 14609
rect 21361 14600 21373 14603
rect 21324 14572 21373 14600
rect 21324 14560 21330 14572
rect 21361 14569 21373 14572
rect 21407 14569 21419 14603
rect 21361 14563 21419 14569
rect 21450 14560 21456 14612
rect 21508 14600 21514 14612
rect 24578 14600 24584 14612
rect 21508 14572 24440 14600
rect 24539 14572 24584 14600
rect 21508 14560 21514 14572
rect 3050 14492 3056 14544
rect 3108 14532 3114 14544
rect 5258 14532 5264 14544
rect 3108 14504 5264 14532
rect 3108 14492 3114 14504
rect 5258 14492 5264 14504
rect 5316 14492 5322 14544
rect 7834 14492 7840 14544
rect 7892 14532 7898 14544
rect 7892 14504 9260 14532
rect 7892 14492 7898 14504
rect 1670 14464 1676 14476
rect 1631 14436 1676 14464
rect 1670 14424 1676 14436
rect 1728 14424 1734 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 7006 14464 7012 14476
rect 4111 14436 7012 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 7374 14424 7380 14476
rect 7432 14464 7438 14476
rect 7653 14467 7711 14473
rect 7653 14464 7665 14467
rect 7432 14436 7665 14464
rect 7432 14424 7438 14436
rect 7653 14433 7665 14436
rect 7699 14464 7711 14467
rect 9030 14464 9036 14476
rect 7699 14436 9036 14464
rect 7699 14433 7711 14436
rect 7653 14427 7711 14433
rect 9030 14424 9036 14436
rect 9088 14464 9094 14476
rect 9125 14467 9183 14473
rect 9125 14464 9137 14467
rect 9088 14436 9137 14464
rect 9088 14424 9094 14436
rect 9125 14433 9137 14436
rect 9171 14433 9183 14467
rect 9232 14464 9260 14504
rect 10428 14504 12434 14532
rect 10428 14464 10456 14504
rect 9232 14436 10456 14464
rect 9125 14427 9183 14433
rect 10594 14424 10600 14476
rect 10652 14464 10658 14476
rect 10870 14464 10876 14476
rect 10652 14436 10876 14464
rect 10652 14424 10658 14436
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11606 14424 11612 14476
rect 11664 14464 11670 14476
rect 11793 14467 11851 14473
rect 11793 14464 11805 14467
rect 11664 14436 11805 14464
rect 11664 14424 11670 14436
rect 11793 14433 11805 14436
rect 11839 14433 11851 14467
rect 12158 14464 12164 14476
rect 12119 14436 12164 14464
rect 11793 14427 11851 14433
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 12406 14464 12434 14504
rect 12618 14492 12624 14544
rect 12676 14532 12682 14544
rect 12894 14532 12900 14544
rect 12676 14504 12900 14532
rect 12676 14492 12682 14504
rect 12894 14492 12900 14504
rect 12952 14532 12958 14544
rect 12952 14504 13492 14532
rect 12952 14492 12958 14504
rect 13354 14464 13360 14476
rect 12406 14436 13360 14464
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 13464 14464 13492 14504
rect 13630 14492 13636 14544
rect 13688 14532 13694 14544
rect 13725 14535 13783 14541
rect 13725 14532 13737 14535
rect 13688 14504 13737 14532
rect 13688 14492 13694 14504
rect 13725 14501 13737 14504
rect 13771 14532 13783 14535
rect 15194 14532 15200 14544
rect 13771 14504 15200 14532
rect 13771 14501 13783 14504
rect 13725 14495 13783 14501
rect 15194 14492 15200 14504
rect 15252 14492 15258 14544
rect 15470 14532 15476 14544
rect 15431 14504 15476 14532
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 16022 14492 16028 14544
rect 16080 14532 16086 14544
rect 17586 14532 17592 14544
rect 16080 14504 17592 14532
rect 16080 14492 16086 14504
rect 17586 14492 17592 14504
rect 17644 14492 17650 14544
rect 18782 14492 18788 14544
rect 18840 14532 18846 14544
rect 24302 14532 24308 14544
rect 18840 14504 24308 14532
rect 18840 14492 18846 14504
rect 24302 14492 24308 14504
rect 24360 14492 24366 14544
rect 24412 14532 24440 14572
rect 24578 14560 24584 14572
rect 24636 14560 24642 14612
rect 25222 14600 25228 14612
rect 25183 14572 25228 14600
rect 25222 14560 25228 14572
rect 25280 14560 25286 14612
rect 26142 14532 26148 14544
rect 24412 14504 26148 14532
rect 26142 14492 26148 14504
rect 26200 14492 26206 14544
rect 14642 14464 14648 14476
rect 13464 14436 14648 14464
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 18414 14424 18420 14476
rect 18472 14464 18478 14476
rect 18472 14436 21496 14464
rect 18472 14424 18478 14436
rect 2958 14356 2964 14408
rect 3016 14396 3022 14408
rect 4157 14399 4215 14405
rect 3016 14368 4108 14396
rect 3016 14356 3022 14368
rect 3234 14288 3240 14340
rect 3292 14328 3298 14340
rect 3421 14331 3479 14337
rect 3421 14328 3433 14331
rect 3292 14300 3433 14328
rect 3292 14288 3298 14300
rect 3421 14297 3433 14300
rect 3467 14297 3479 14331
rect 4080 14328 4108 14368
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4614 14396 4620 14408
rect 4203 14368 4620 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 4798 14396 4804 14408
rect 4759 14368 4804 14396
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 8386 14396 8392 14408
rect 8347 14368 8392 14396
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 13081 14399 13139 14405
rect 13081 14396 13093 14399
rect 12952 14368 13093 14396
rect 12952 14356 12958 14368
rect 13081 14365 13093 14368
rect 13127 14365 13139 14399
rect 13081 14359 13139 14365
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14396 13323 14399
rect 14182 14396 14188 14408
rect 13311 14368 14188 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 15654 14396 15660 14408
rect 15615 14368 15660 14396
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 16574 14396 16580 14408
rect 16535 14368 16580 14396
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 17310 14396 17316 14408
rect 16807 14368 17316 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 18874 14396 18880 14408
rect 18835 14368 18880 14396
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 19426 14396 19432 14408
rect 19387 14368 19432 14396
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 20533 14399 20591 14405
rect 20533 14365 20545 14399
rect 20579 14365 20591 14399
rect 20714 14396 20720 14408
rect 20675 14368 20720 14396
rect 20533 14359 20591 14365
rect 5629 14331 5687 14337
rect 5629 14328 5641 14331
rect 4080 14300 5641 14328
rect 3421 14291 3479 14297
rect 5629 14297 5641 14300
rect 5675 14297 5687 14331
rect 5629 14291 5687 14297
rect 5718 14288 5724 14340
rect 5776 14328 5782 14340
rect 7374 14328 7380 14340
rect 5776 14300 6210 14328
rect 7335 14300 7380 14328
rect 5776 14288 5782 14300
rect 7374 14288 7380 14300
rect 7432 14288 7438 14340
rect 8110 14288 8116 14340
rect 8168 14328 8174 14340
rect 9122 14328 9128 14340
rect 8168 14300 9128 14328
rect 8168 14288 8174 14300
rect 9122 14288 9128 14300
rect 9180 14288 9186 14340
rect 9398 14328 9404 14340
rect 9359 14300 9404 14328
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 9950 14288 9956 14340
rect 10008 14288 10014 14340
rect 11885 14331 11943 14337
rect 11885 14297 11897 14331
rect 11931 14297 11943 14331
rect 11885 14291 11943 14297
rect 8570 14260 8576 14272
rect 8531 14232 8576 14260
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 9582 14220 9588 14272
rect 9640 14260 9646 14272
rect 11514 14260 11520 14272
rect 9640 14232 11520 14260
rect 9640 14220 9646 14232
rect 11514 14220 11520 14232
rect 11572 14220 11578 14272
rect 11893 14260 11921 14291
rect 12158 14288 12164 14340
rect 12216 14328 12222 14340
rect 14369 14331 14427 14337
rect 14369 14328 14381 14331
rect 12216 14300 14381 14328
rect 12216 14288 12222 14300
rect 14369 14297 14381 14300
rect 14415 14297 14427 14331
rect 14369 14291 14427 14297
rect 14461 14331 14519 14337
rect 14461 14297 14473 14331
rect 14507 14297 14519 14331
rect 14461 14291 14519 14297
rect 15013 14331 15071 14337
rect 15013 14297 15025 14331
rect 15059 14328 15071 14331
rect 15194 14328 15200 14340
rect 15059 14300 15200 14328
rect 15059 14297 15071 14300
rect 15013 14291 15071 14297
rect 11974 14260 11980 14272
rect 11893 14232 11980 14260
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14476 14260 14504 14291
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 17402 14288 17408 14340
rect 17460 14328 17466 14340
rect 17497 14331 17555 14337
rect 17497 14328 17509 14331
rect 17460 14300 17509 14328
rect 17460 14288 17466 14300
rect 17497 14297 17509 14300
rect 17543 14297 17555 14331
rect 17497 14291 17555 14297
rect 18049 14331 18107 14337
rect 18049 14297 18061 14331
rect 18095 14297 18107 14331
rect 18049 14291 18107 14297
rect 18141 14331 18199 14337
rect 18141 14297 18153 14331
rect 18187 14328 18199 14331
rect 19978 14328 19984 14340
rect 18187 14300 19984 14328
rect 18187 14297 18199 14300
rect 18141 14291 18199 14297
rect 13872 14232 14504 14260
rect 13872 14220 13878 14232
rect 14550 14220 14556 14272
rect 14608 14260 14614 14272
rect 16390 14260 16396 14272
rect 14608 14232 16396 14260
rect 14608 14220 14614 14232
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 18064 14260 18092 14291
rect 19978 14288 19984 14300
rect 20036 14288 20042 14340
rect 20548 14328 20576 14359
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 21468 14405 21496 14436
rect 21726 14424 21732 14476
rect 21784 14464 21790 14476
rect 33597 14467 33655 14473
rect 33597 14464 33609 14467
rect 21784 14436 33609 14464
rect 21784 14424 21790 14436
rect 33597 14433 33609 14436
rect 33643 14433 33655 14467
rect 33597 14427 33655 14433
rect 21453 14399 21511 14405
rect 21453 14365 21465 14399
rect 21499 14396 21511 14399
rect 21542 14396 21548 14408
rect 21499 14368 21548 14396
rect 21499 14365 21511 14368
rect 21453 14359 21511 14365
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 22462 14396 22468 14408
rect 22423 14368 22468 14396
rect 22462 14356 22468 14368
rect 22520 14356 22526 14408
rect 22646 14396 22652 14408
rect 22607 14368 22652 14396
rect 22646 14356 22652 14368
rect 22704 14356 22710 14408
rect 23290 14396 23296 14408
rect 23251 14368 23296 14396
rect 23290 14356 23296 14368
rect 23348 14356 23354 14408
rect 23474 14356 23480 14408
rect 23532 14396 23538 14408
rect 23753 14399 23811 14405
rect 23753 14396 23765 14399
rect 23532 14368 23765 14396
rect 23532 14356 23538 14368
rect 23753 14365 23765 14368
rect 23799 14365 23811 14399
rect 23753 14359 23811 14365
rect 24765 14399 24823 14405
rect 24765 14365 24777 14399
rect 24811 14396 24823 14399
rect 25222 14396 25228 14408
rect 24811 14368 25228 14396
rect 24811 14365 24823 14368
rect 24765 14359 24823 14365
rect 25222 14356 25228 14368
rect 25280 14356 25286 14408
rect 25409 14399 25467 14405
rect 25409 14365 25421 14399
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 33689 14399 33747 14405
rect 33689 14365 33701 14399
rect 33735 14396 33747 14399
rect 36906 14396 36912 14408
rect 33735 14368 36912 14396
rect 33735 14365 33747 14368
rect 33689 14359 33747 14365
rect 23845 14331 23903 14337
rect 23845 14328 23857 14331
rect 20548 14300 23857 14328
rect 23845 14297 23857 14300
rect 23891 14297 23903 14331
rect 25424 14328 25452 14359
rect 36906 14356 36912 14368
rect 36964 14356 36970 14408
rect 23845 14291 23903 14297
rect 24780 14300 25452 14328
rect 24780 14272 24808 14300
rect 18506 14260 18512 14272
rect 18064 14232 18512 14260
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 18598 14220 18604 14272
rect 18656 14260 18662 14272
rect 19242 14260 19248 14272
rect 18656 14232 19248 14260
rect 18656 14220 18662 14232
rect 19242 14220 19248 14232
rect 19300 14260 19306 14272
rect 21450 14260 21456 14272
rect 19300 14232 21456 14260
rect 19300 14220 19306 14232
rect 21450 14220 21456 14232
rect 21508 14220 21514 14272
rect 22005 14263 22063 14269
rect 22005 14229 22017 14263
rect 22051 14260 22063 14263
rect 22370 14260 22376 14272
rect 22051 14232 22376 14260
rect 22051 14229 22063 14232
rect 22005 14223 22063 14229
rect 22370 14220 22376 14232
rect 22428 14220 22434 14272
rect 24762 14220 24768 14272
rect 24820 14220 24826 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 4706 14056 4712 14068
rect 1728 14028 4108 14056
rect 1728 14016 1734 14028
rect 1302 13948 1308 14000
rect 1360 13988 1366 14000
rect 1360 13960 2346 13988
rect 1360 13948 1366 13960
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 3605 13991 3663 13997
rect 3605 13988 3617 13991
rect 3568 13960 3617 13988
rect 3568 13948 3574 13960
rect 3605 13957 3617 13960
rect 3651 13957 3663 13991
rect 3605 13951 3663 13957
rect 4080 13929 4108 14028
rect 4356 14028 4712 14056
rect 4356 13997 4384 14028
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 6822 14056 6828 14068
rect 6783 14028 6828 14056
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 8570 14016 8576 14068
rect 8628 14056 8634 14068
rect 13630 14056 13636 14068
rect 8628 14028 12434 14056
rect 13591 14028 13636 14056
rect 8628 14016 8634 14028
rect 4341 13991 4399 13997
rect 4341 13957 4353 13991
rect 4387 13957 4399 13991
rect 4341 13951 4399 13957
rect 5350 13948 5356 14000
rect 5408 13948 5414 14000
rect 5810 13948 5816 14000
rect 5868 13988 5874 14000
rect 5868 13960 7130 13988
rect 5868 13948 5874 13960
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 9306 13988 9312 14000
rect 8260 13960 8616 13988
rect 9267 13960 9312 13988
rect 8260 13948 8266 13960
rect 8588 13929 8616 13960
rect 9306 13948 9312 13960
rect 9364 13948 9370 14000
rect 11606 13948 11612 14000
rect 11664 13988 11670 14000
rect 11885 13991 11943 13997
rect 11885 13988 11897 13991
rect 11664 13960 11897 13988
rect 11664 13948 11670 13960
rect 11885 13957 11897 13960
rect 11931 13957 11943 13991
rect 12406 13988 12434 14028
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 16025 14059 16083 14065
rect 16025 14025 16037 14059
rect 16071 14056 16083 14059
rect 16114 14056 16120 14068
rect 16071 14028 16120 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 16850 14056 16856 14068
rect 16811 14028 16856 14056
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 17954 14056 17960 14068
rect 17915 14028 17960 14056
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18601 14059 18659 14065
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 19150 14056 19156 14068
rect 18647 14028 19156 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 19978 14056 19984 14068
rect 19939 14028 19984 14056
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 21453 14059 21511 14065
rect 21453 14025 21465 14059
rect 21499 14056 21511 14059
rect 22370 14056 22376 14068
rect 21499 14028 22376 14056
rect 21499 14025 21511 14028
rect 21453 14019 21511 14025
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 24026 14056 24032 14068
rect 22572 14028 24032 14056
rect 14090 13988 14096 14000
rect 12406 13960 14096 13988
rect 11885 13951 11943 13957
rect 14090 13948 14096 13960
rect 14148 13948 14154 14000
rect 14918 13988 14924 14000
rect 14879 13960 14924 13988
rect 14918 13948 14924 13960
rect 14976 13948 14982 14000
rect 15473 13991 15531 13997
rect 15473 13957 15485 13991
rect 15519 13988 15531 13991
rect 15519 13960 16068 13988
rect 15519 13957 15531 13960
rect 15473 13951 15531 13957
rect 16040 13932 16068 13960
rect 17310 13948 17316 14000
rect 17368 13988 17374 14000
rect 17368 13960 20852 13988
rect 17368 13948 17374 13960
rect 4065 13923 4123 13929
rect 4065 13889 4077 13923
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13889 8631 13923
rect 9030 13920 9036 13932
rect 8991 13892 9036 13920
rect 8573 13883 8631 13889
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 10410 13880 10416 13932
rect 10468 13880 10474 13932
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 12986 13920 12992 13932
rect 12584 13892 12992 13920
rect 12584 13880 12590 13892
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 4430 13812 4436 13864
rect 4488 13852 4494 13864
rect 11146 13852 11152 13864
rect 4488 13824 11152 13852
rect 4488 13812 4494 13824
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 11514 13812 11520 13864
rect 11572 13852 11578 13864
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11572 13824 11805 13852
rect 11572 13812 11578 13824
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 11974 13812 11980 13864
rect 12032 13852 12038 13864
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 12032 13824 12081 13852
rect 12032 13812 12038 13824
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 13630 13852 13636 13864
rect 12768 13824 13636 13852
rect 12768 13812 12774 13824
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 14090 13852 14096 13864
rect 14051 13824 14096 13852
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 14277 13855 14335 13861
rect 14277 13821 14289 13855
rect 14323 13852 14335 13855
rect 14458 13852 14464 13864
rect 14323 13824 14464 13852
rect 14323 13821 14335 13824
rect 14277 13815 14335 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15102 13852 15108 13864
rect 14875 13824 15108 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 5813 13787 5871 13793
rect 5813 13753 5825 13787
rect 5859 13784 5871 13787
rect 6086 13784 6092 13796
rect 5859 13756 6092 13784
rect 5859 13753 5871 13756
rect 5813 13747 5871 13753
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10781 13787 10839 13793
rect 10781 13784 10793 13787
rect 10376 13756 10793 13784
rect 10376 13744 10382 13756
rect 10781 13753 10793 13756
rect 10827 13753 10839 13787
rect 15654 13784 15660 13796
rect 10781 13747 10839 13753
rect 13004 13756 15660 13784
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 1838 13719 1896 13725
rect 1838 13716 1850 13719
rect 1728 13688 1850 13716
rect 1728 13676 1734 13688
rect 1838 13685 1850 13688
rect 1884 13685 1896 13719
rect 1838 13679 1896 13685
rect 6270 13676 6276 13728
rect 6328 13716 6334 13728
rect 8202 13716 8208 13728
rect 6328 13688 8208 13716
rect 6328 13676 6334 13688
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8315 13719 8373 13725
rect 8315 13685 8327 13719
rect 8361 13716 8373 13719
rect 8662 13716 8668 13728
rect 8361 13688 8668 13716
rect 8361 13685 8373 13688
rect 8315 13679 8373 13685
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 13004 13716 13032 13756
rect 15654 13744 15660 13756
rect 15712 13784 15718 13796
rect 15948 13784 15976 13883
rect 16022 13880 16028 13932
rect 16080 13880 16086 13932
rect 18322 13880 18328 13932
rect 18380 13920 18386 13932
rect 18417 13923 18475 13929
rect 18417 13920 18429 13923
rect 18380 13892 18429 13920
rect 18380 13880 18386 13892
rect 18417 13889 18429 13892
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 20824 13929 20852 13960
rect 21542 13948 21548 14000
rect 21600 13988 21606 14000
rect 22572 13988 22600 14028
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 24302 14016 24308 14068
rect 24360 14056 24366 14068
rect 27614 14056 27620 14068
rect 24360 14028 27620 14056
rect 24360 14016 24366 14028
rect 27614 14016 27620 14028
rect 27672 14016 27678 14068
rect 35069 14059 35127 14065
rect 35069 14025 35081 14059
rect 35115 14056 35127 14059
rect 35115 14028 35894 14056
rect 35115 14025 35127 14028
rect 35069 14019 35127 14025
rect 21600 13960 22600 13988
rect 22649 13991 22707 13997
rect 21600 13948 21606 13960
rect 22649 13957 22661 13991
rect 22695 13988 22707 13991
rect 23566 13988 23572 14000
rect 22695 13960 23572 13988
rect 22695 13957 22707 13960
rect 22649 13951 22707 13957
rect 23566 13948 23572 13960
rect 23624 13948 23630 14000
rect 19337 13923 19395 13929
rect 19337 13920 19349 13923
rect 19300 13892 19349 13920
rect 19300 13880 19306 13892
rect 19337 13889 19349 13892
rect 19383 13889 19395 13923
rect 19337 13883 19395 13889
rect 20809 13923 20867 13929
rect 20809 13889 20821 13923
rect 20855 13889 20867 13923
rect 23474 13920 23480 13932
rect 23435 13892 23480 13920
rect 20809 13883 20867 13889
rect 23474 13880 23480 13892
rect 23532 13880 23538 13932
rect 29270 13880 29276 13932
rect 29328 13920 29334 13932
rect 34885 13923 34943 13929
rect 34885 13920 34897 13923
rect 29328 13892 34897 13920
rect 29328 13880 29334 13892
rect 34885 13889 34897 13892
rect 34931 13889 34943 13923
rect 35866 13920 35894 14028
rect 38013 13923 38071 13929
rect 38013 13920 38025 13923
rect 35866 13892 38025 13920
rect 34885 13883 34943 13889
rect 38013 13889 38025 13892
rect 38059 13889 38071 13923
rect 38013 13883 38071 13889
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19484 13824 19533 13852
rect 19484 13812 19490 13824
rect 19521 13821 19533 13824
rect 19567 13821 19579 13855
rect 20990 13852 20996 13864
rect 20951 13824 20996 13852
rect 19521 13815 19579 13821
rect 20990 13812 20996 13824
rect 21048 13812 21054 13864
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13852 22523 13855
rect 22554 13852 22560 13864
rect 22511 13824 22560 13852
rect 22511 13821 22523 13824
rect 22465 13815 22523 13821
rect 22554 13812 22560 13824
rect 22612 13812 22618 13864
rect 22741 13855 22799 13861
rect 22741 13821 22753 13855
rect 22787 13852 22799 13855
rect 23937 13855 23995 13861
rect 23937 13852 23949 13855
rect 22787 13824 23949 13852
rect 22787 13821 22799 13824
rect 22741 13815 22799 13821
rect 23937 13821 23949 13824
rect 23983 13821 23995 13855
rect 23937 13815 23995 13821
rect 15712 13756 15976 13784
rect 15712 13744 15718 13756
rect 13170 13716 13176 13728
rect 9364 13688 13032 13716
rect 13131 13688 13176 13716
rect 9364 13676 9370 13688
rect 13170 13676 13176 13688
rect 13228 13676 13234 13728
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 14366 13716 14372 13728
rect 13412 13688 14372 13716
rect 13412 13676 13418 13688
rect 14366 13676 14372 13688
rect 14424 13676 14430 13728
rect 14642 13676 14648 13728
rect 14700 13716 14706 13728
rect 21910 13716 21916 13728
rect 14700 13688 21916 13716
rect 14700 13676 14706 13688
rect 21910 13676 21916 13688
rect 21968 13676 21974 13728
rect 22278 13676 22284 13728
rect 22336 13716 22342 13728
rect 23293 13719 23351 13725
rect 23293 13716 23305 13719
rect 22336 13688 23305 13716
rect 22336 13676 22342 13688
rect 23293 13685 23305 13688
rect 23339 13685 23351 13719
rect 38194 13716 38200 13728
rect 38155 13688 38200 13716
rect 23293 13679 23351 13685
rect 38194 13676 38200 13688
rect 38252 13676 38258 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2222 13472 2228 13524
rect 2280 13512 2286 13524
rect 7929 13515 7987 13521
rect 2280 13484 7696 13512
rect 2280 13472 2286 13484
rect 7466 13444 7472 13456
rect 7208 13416 7472 13444
rect 1578 13376 1584 13388
rect 1491 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13376 1642 13388
rect 2866 13376 2872 13388
rect 1636 13348 2872 13376
rect 1636 13336 1642 13348
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13376 3387 13379
rect 4706 13376 4712 13388
rect 3375 13348 4712 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 4985 13379 5043 13385
rect 4985 13345 4997 13379
rect 5031 13376 5043 13379
rect 7208 13376 7236 13416
rect 7466 13404 7472 13416
rect 7524 13404 7530 13456
rect 5031 13348 7236 13376
rect 5031 13345 5043 13348
rect 4985 13339 5043 13345
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13308 4307 13311
rect 5442 13308 5448 13320
rect 4295 13280 5448 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 7282 13268 7288 13320
rect 7340 13308 7346 13320
rect 7668 13310 7696 13484
rect 7929 13481 7941 13515
rect 7975 13512 7987 13515
rect 10686 13512 10692 13524
rect 7975 13484 10692 13512
rect 7975 13481 7987 13484
rect 7929 13475 7987 13481
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13512 10931 13515
rect 11882 13512 11888 13524
rect 10919 13484 11888 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 13446 13512 13452 13524
rect 12952 13484 13452 13512
rect 12952 13472 12958 13484
rect 13446 13472 13452 13484
rect 13504 13512 13510 13524
rect 21177 13515 21235 13521
rect 13504 13484 17724 13512
rect 13504 13472 13510 13484
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 13354 13444 13360 13456
rect 8527 13416 9260 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 9088 13348 9137 13376
rect 9088 13336 9094 13348
rect 9125 13345 9137 13348
rect 9171 13345 9183 13379
rect 9232 13376 9260 13416
rect 11348 13416 13360 13444
rect 10778 13376 10784 13388
rect 9232 13348 10784 13376
rect 9125 13339 9183 13345
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 11348 13385 11376 13416
rect 13354 13404 13360 13416
rect 13412 13404 13418 13456
rect 13633 13447 13691 13453
rect 13633 13413 13645 13447
rect 13679 13444 13691 13447
rect 16022 13444 16028 13456
rect 13679 13416 16028 13444
rect 13679 13413 13691 13416
rect 13633 13407 13691 13413
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13376 12035 13379
rect 13722 13376 13728 13388
rect 12023 13348 13728 13376
rect 12023 13345 12035 13348
rect 11977 13339 12035 13345
rect 13722 13336 13728 13348
rect 13780 13376 13786 13388
rect 14553 13379 14611 13385
rect 14553 13376 14565 13379
rect 13780 13348 14565 13376
rect 13780 13336 13786 13348
rect 14553 13345 14565 13348
rect 14599 13345 14611 13379
rect 14553 13339 14611 13345
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15562 13376 15568 13388
rect 15252 13348 15568 13376
rect 15252 13336 15258 13348
rect 15562 13336 15568 13348
rect 15620 13336 15626 13388
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 15896 13348 16313 13376
rect 15896 13336 15902 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16758 13376 16764 13388
rect 16719 13348 16764 13376
rect 16301 13339 16359 13345
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 17696 13385 17724 13484
rect 21177 13481 21189 13515
rect 21223 13512 21235 13515
rect 23382 13512 23388 13524
rect 21223 13484 23388 13512
rect 21223 13481 21235 13484
rect 21177 13475 21235 13481
rect 23382 13472 23388 13484
rect 23440 13472 23446 13524
rect 23477 13515 23535 13521
rect 23477 13481 23489 13515
rect 23523 13512 23535 13515
rect 23566 13512 23572 13524
rect 23523 13484 23572 13512
rect 23523 13481 23535 13484
rect 23477 13475 23535 13481
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 26142 13472 26148 13524
rect 26200 13512 26206 13524
rect 30653 13515 30711 13521
rect 30653 13512 30665 13515
rect 26200 13484 30665 13512
rect 26200 13472 26206 13484
rect 30653 13481 30665 13484
rect 30699 13481 30711 13515
rect 30653 13475 30711 13481
rect 24762 13444 24768 13456
rect 19306 13416 24768 13444
rect 17681 13379 17739 13385
rect 17681 13345 17693 13379
rect 17727 13345 17739 13379
rect 17681 13339 17739 13345
rect 7745 13311 7803 13317
rect 7745 13310 7757 13311
rect 7340 13280 7385 13308
rect 7668 13282 7757 13310
rect 7340 13268 7346 13280
rect 7745 13277 7757 13282
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 8352 13280 8401 13308
rect 8352 13268 8358 13280
rect 8389 13277 8401 13280
rect 8435 13308 8447 13311
rect 8478 13308 8484 13320
rect 8435 13280 8484 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 10744 13280 11529 13308
rect 10744 13268 10750 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 16114 13308 16120 13320
rect 16075 13280 16120 13308
rect 11517 13271 11575 13277
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13308 17923 13311
rect 17954 13308 17960 13320
rect 17911 13280 17960 13308
rect 17911 13277 17923 13280
rect 17865 13271 17923 13277
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 1762 13200 1768 13252
rect 1820 13240 1826 13252
rect 1857 13243 1915 13249
rect 1857 13240 1869 13243
rect 1820 13212 1869 13240
rect 1820 13200 1826 13212
rect 1857 13209 1869 13212
rect 1903 13209 1915 13243
rect 1857 13203 1915 13209
rect 1964 13212 2346 13240
rect 1394 13132 1400 13184
rect 1452 13172 1458 13184
rect 1964 13172 1992 13212
rect 6454 13200 6460 13252
rect 6512 13200 6518 13252
rect 7009 13243 7067 13249
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 8110 13240 8116 13252
rect 7055 13212 8116 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 8110 13200 8116 13212
rect 8168 13200 8174 13252
rect 9306 13200 9312 13252
rect 9364 13240 9370 13252
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 9364 13212 9413 13240
rect 9364 13200 9370 13212
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 9401 13203 9459 13209
rect 10042 13200 10048 13252
rect 10100 13200 10106 13252
rect 12710 13240 12716 13252
rect 10704 13212 12716 13240
rect 4062 13172 4068 13184
rect 1452 13144 1992 13172
rect 4023 13144 4068 13172
rect 1452 13132 1458 13144
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 5537 13175 5595 13181
rect 5537 13141 5549 13175
rect 5583 13172 5595 13175
rect 6086 13172 6092 13184
rect 5583 13144 6092 13172
rect 5583 13141 5595 13144
rect 5537 13135 5595 13141
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 7282 13132 7288 13184
rect 7340 13172 7346 13184
rect 8478 13172 8484 13184
rect 7340 13144 8484 13172
rect 7340 13132 7346 13144
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 8570 13132 8576 13184
rect 8628 13172 8634 13184
rect 10704 13172 10732 13212
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 12894 13200 12900 13252
rect 12952 13240 12958 13252
rect 13081 13243 13139 13249
rect 13081 13240 13093 13243
rect 12952 13212 13093 13240
rect 12952 13200 12958 13212
rect 13081 13209 13093 13212
rect 13127 13209 13139 13243
rect 13081 13203 13139 13209
rect 13173 13243 13231 13249
rect 13173 13209 13185 13243
rect 13219 13240 13231 13243
rect 13354 13240 13360 13252
rect 13219 13212 13360 13240
rect 13219 13209 13231 13212
rect 13173 13203 13231 13209
rect 13354 13200 13360 13212
rect 13412 13200 13418 13252
rect 14642 13200 14648 13252
rect 14700 13240 14706 13252
rect 15197 13243 15255 13249
rect 14700 13212 14745 13240
rect 14700 13200 14706 13212
rect 15197 13209 15209 13243
rect 15243 13240 15255 13243
rect 15654 13240 15660 13252
rect 15243 13212 15660 13240
rect 15243 13209 15255 13212
rect 15197 13203 15255 13209
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 19306 13240 19334 13416
rect 24762 13404 24768 13416
rect 24820 13404 24826 13456
rect 19518 13336 19524 13388
rect 19576 13376 19582 13388
rect 19576 13348 20300 13376
rect 19576 13336 19582 13348
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13308 19947 13311
rect 19978 13308 19984 13320
rect 19935 13280 19984 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13308 20131 13311
rect 20162 13308 20168 13320
rect 20119 13280 20168 13308
rect 20119 13277 20131 13280
rect 20073 13271 20131 13277
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 20272 13308 20300 13348
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 21637 13379 21695 13385
rect 21637 13376 21649 13379
rect 20864 13348 21649 13376
rect 20864 13336 20870 13348
rect 21637 13345 21649 13348
rect 21683 13345 21695 13379
rect 22370 13376 22376 13388
rect 22331 13348 22376 13376
rect 21637 13339 21695 13345
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 22554 13336 22560 13388
rect 22612 13376 22618 13388
rect 22649 13379 22707 13385
rect 22649 13376 22661 13379
rect 22612 13348 22661 13376
rect 22612 13336 22618 13348
rect 22649 13345 22661 13348
rect 22695 13376 22707 13379
rect 23014 13376 23020 13388
rect 22695 13348 23020 13376
rect 22695 13345 22707 13348
rect 22649 13339 22707 13345
rect 23014 13336 23020 13348
rect 23072 13336 23078 13388
rect 20993 13311 21051 13317
rect 20993 13308 21005 13311
rect 20272 13280 21005 13308
rect 20993 13277 21005 13280
rect 21039 13277 21051 13311
rect 23658 13308 23664 13320
rect 23619 13280 23664 13308
rect 20993 13271 21051 13277
rect 23658 13268 23664 13280
rect 23716 13268 23722 13320
rect 30742 13308 30748 13320
rect 30703 13280 30748 13308
rect 30742 13268 30748 13280
rect 30800 13268 30806 13320
rect 15764 13212 19334 13240
rect 22465 13243 22523 13249
rect 8628 13144 10732 13172
rect 8628 13132 8634 13144
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 12158 13172 12164 13184
rect 10836 13144 12164 13172
rect 10836 13132 10842 13144
rect 12158 13132 12164 13144
rect 12216 13132 12222 13184
rect 12342 13132 12348 13184
rect 12400 13172 12406 13184
rect 15764 13172 15792 13212
rect 22465 13209 22477 13243
rect 22511 13240 22523 13243
rect 22830 13240 22836 13252
rect 22511 13212 22836 13240
rect 22511 13209 22523 13212
rect 22465 13203 22523 13209
rect 22830 13200 22836 13212
rect 22888 13200 22894 13252
rect 18322 13172 18328 13184
rect 12400 13144 15792 13172
rect 18283 13144 18328 13172
rect 12400 13132 12406 13144
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 20533 13175 20591 13181
rect 20533 13141 20545 13175
rect 20579 13172 20591 13175
rect 21082 13172 21088 13184
rect 20579 13144 21088 13172
rect 20579 13141 20591 13144
rect 20533 13135 20591 13141
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 8570 12968 8576 12980
rect 7331 12940 8576 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 8570 12928 8576 12940
rect 8628 12928 8634 12980
rect 9030 12928 9036 12980
rect 9088 12968 9094 12980
rect 9125 12971 9183 12977
rect 9125 12968 9137 12971
rect 9088 12940 9137 12968
rect 9088 12928 9094 12940
rect 9125 12937 9137 12940
rect 9171 12937 9183 12971
rect 10594 12968 10600 12980
rect 9125 12931 9183 12937
rect 9416 12940 10600 12968
rect 3326 12900 3332 12912
rect 3287 12872 3332 12900
rect 3326 12860 3332 12872
rect 3384 12860 3390 12912
rect 3694 12860 3700 12912
rect 3752 12900 3758 12912
rect 5629 12903 5687 12909
rect 3752 12872 4462 12900
rect 3752 12860 3758 12872
rect 5629 12869 5641 12903
rect 5675 12900 5687 12903
rect 6270 12900 6276 12912
rect 5675 12872 6276 12900
rect 5675 12869 5687 12872
rect 5629 12863 5687 12869
rect 6270 12860 6276 12872
rect 6328 12860 6334 12912
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 7837 12903 7895 12909
rect 7837 12900 7849 12903
rect 6788 12872 7849 12900
rect 6788 12860 6794 12872
rect 7837 12869 7849 12872
rect 7883 12869 7895 12903
rect 7837 12863 7895 12869
rect 2222 12792 2228 12844
rect 2280 12792 2286 12844
rect 3605 12835 3663 12841
rect 3605 12801 3617 12835
rect 3651 12801 3663 12835
rect 3605 12795 3663 12801
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12832 6607 12835
rect 6822 12832 6828 12844
rect 6595 12804 6828 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 1581 12767 1639 12773
rect 1581 12764 1593 12767
rect 1544 12736 1593 12764
rect 1544 12724 1550 12736
rect 1581 12733 1593 12736
rect 1627 12733 1639 12767
rect 1581 12727 1639 12733
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 3620 12764 3648 12795
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 7156 12804 7205 12832
rect 7156 12792 7162 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 9416 12832 9444 12940
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 10689 12971 10747 12977
rect 10689 12937 10701 12971
rect 10735 12968 10747 12971
rect 11514 12968 11520 12980
rect 10735 12940 11520 12968
rect 10735 12937 10747 12940
rect 10689 12931 10747 12937
rect 11514 12928 11520 12940
rect 11572 12968 11578 12980
rect 11882 12968 11888 12980
rect 11572 12940 11888 12968
rect 11572 12928 11578 12940
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 14829 12971 14887 12977
rect 12216 12940 14780 12968
rect 12216 12928 12222 12940
rect 12618 12900 12624 12912
rect 10060 12872 12624 12900
rect 10060 12841 10088 12872
rect 12618 12860 12624 12872
rect 12676 12860 12682 12912
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 14550 12900 14556 12912
rect 12768 12872 14556 12900
rect 12768 12860 12774 12872
rect 14550 12860 14556 12872
rect 14608 12860 14614 12912
rect 7340 12804 9444 12832
rect 10045 12835 10103 12841
rect 7340 12792 7346 12804
rect 10045 12801 10057 12835
rect 10091 12801 10103 12835
rect 12069 12835 12127 12841
rect 10045 12795 10103 12801
rect 10152 12804 12020 12832
rect 2924 12736 3648 12764
rect 5905 12767 5963 12773
rect 2924 12724 2930 12736
rect 3528 12640 3556 12736
rect 5905 12733 5917 12767
rect 5951 12733 5963 12767
rect 5905 12727 5963 12733
rect 3510 12588 3516 12640
rect 3568 12588 3574 12640
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 4157 12631 4215 12637
rect 4157 12628 4169 12631
rect 4120 12600 4169 12628
rect 4120 12588 4126 12600
rect 4157 12597 4169 12600
rect 4203 12597 4215 12631
rect 4157 12591 4215 12597
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 5920 12628 5948 12727
rect 6086 12724 6092 12776
rect 6144 12764 6150 12776
rect 10152 12764 10180 12804
rect 6144 12736 10180 12764
rect 10229 12767 10287 12773
rect 6144 12724 6150 12736
rect 10229 12733 10241 12767
rect 10275 12764 10287 12767
rect 10410 12764 10416 12776
rect 10275 12736 10416 12764
rect 10275 12733 10287 12736
rect 10229 12727 10287 12733
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 10594 12724 10600 12776
rect 10652 12764 10658 12776
rect 11992 12764 12020 12804
rect 12069 12801 12081 12835
rect 12115 12832 12127 12835
rect 12158 12832 12164 12844
rect 12115 12804 12164 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 13170 12792 13176 12844
rect 13228 12832 13234 12844
rect 14752 12841 14780 12940
rect 14829 12937 14841 12971
rect 14875 12968 14887 12971
rect 15746 12968 15752 12980
rect 14875 12940 15752 12968
rect 14875 12937 14887 12940
rect 14829 12931 14887 12937
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 22005 12971 22063 12977
rect 22005 12968 22017 12971
rect 21232 12940 22017 12968
rect 21232 12928 21238 12940
rect 22005 12937 22017 12940
rect 22051 12937 22063 12971
rect 22005 12931 22063 12937
rect 22462 12928 22468 12980
rect 22520 12968 22526 12980
rect 22649 12971 22707 12977
rect 22649 12968 22661 12971
rect 22520 12940 22661 12968
rect 22520 12928 22526 12940
rect 22649 12937 22661 12940
rect 22695 12937 22707 12971
rect 22649 12931 22707 12937
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 24029 12971 24087 12977
rect 24029 12968 24041 12971
rect 22888 12940 24041 12968
rect 22888 12928 22894 12940
rect 24029 12937 24041 12940
rect 24075 12937 24087 12971
rect 24029 12931 24087 12937
rect 15562 12900 15568 12912
rect 15523 12872 15568 12900
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 15654 12860 15660 12912
rect 15712 12900 15718 12912
rect 16117 12903 16175 12909
rect 16117 12900 16129 12903
rect 15712 12872 16129 12900
rect 15712 12860 15718 12872
rect 16117 12869 16129 12872
rect 16163 12900 16175 12903
rect 18230 12900 18236 12912
rect 16163 12872 18236 12900
rect 16163 12869 16175 12872
rect 16117 12863 16175 12869
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 18325 12903 18383 12909
rect 18325 12869 18337 12903
rect 18371 12900 18383 12903
rect 19242 12900 19248 12912
rect 18371 12872 19248 12900
rect 18371 12869 18383 12872
rect 18325 12863 18383 12869
rect 19242 12860 19248 12872
rect 19300 12860 19306 12912
rect 19518 12900 19524 12912
rect 19479 12872 19524 12900
rect 19518 12860 19524 12872
rect 19576 12860 19582 12912
rect 20898 12900 20904 12912
rect 20859 12872 20904 12900
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 21634 12860 21640 12912
rect 21692 12900 21698 12912
rect 21692 12872 23520 12900
rect 21692 12860 21698 12872
rect 14093 12835 14151 12841
rect 14093 12832 14105 12835
rect 13228 12804 14105 12832
rect 13228 12792 13234 12804
rect 14093 12801 14105 12804
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12832 22247 12835
rect 22278 12832 22284 12844
rect 22235 12804 22284 12832
rect 22235 12801 22247 12804
rect 22189 12795 22247 12801
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 23492 12841 23520 12872
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12832 22891 12835
rect 23477 12835 23535 12841
rect 22879 12804 23336 12832
rect 22879 12801 22891 12804
rect 22833 12795 22891 12801
rect 12342 12764 12348 12776
rect 10652 12736 11921 12764
rect 11992 12736 12348 12764
rect 10652 12724 10658 12736
rect 6733 12699 6791 12705
rect 6733 12665 6745 12699
rect 6779 12696 6791 12699
rect 8938 12696 8944 12708
rect 6779 12668 8944 12696
rect 6779 12665 6791 12668
rect 6733 12659 6791 12665
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 9398 12656 9404 12708
rect 9456 12696 9462 12708
rect 11146 12696 11152 12708
rect 9456 12668 11152 12696
rect 9456 12656 9462 12668
rect 11146 12656 11152 12668
rect 11204 12656 11210 12708
rect 11893 12705 11921 12736
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 12526 12764 12532 12776
rect 12487 12736 12532 12764
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 12710 12764 12716 12776
rect 12671 12736 12716 12764
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 15470 12764 15476 12776
rect 15431 12736 15476 12764
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 17494 12764 17500 12776
rect 17455 12736 17500 12764
rect 17494 12724 17500 12736
rect 17552 12724 17558 12776
rect 17678 12764 17684 12776
rect 17639 12736 17684 12764
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 18233 12767 18291 12773
rect 18233 12733 18245 12767
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 11885 12699 11943 12705
rect 11885 12665 11897 12699
rect 11931 12665 11943 12699
rect 12894 12696 12900 12708
rect 12855 12668 12900 12696
rect 11885 12659 11943 12665
rect 12894 12656 12900 12668
rect 12952 12696 12958 12708
rect 13170 12696 13176 12708
rect 12952 12668 13176 12696
rect 12952 12656 12958 12668
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 14277 12699 14335 12705
rect 14277 12665 14289 12699
rect 14323 12696 14335 12699
rect 15194 12696 15200 12708
rect 14323 12668 15200 12696
rect 14323 12665 14335 12668
rect 14277 12659 14335 12665
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 17310 12696 17316 12708
rect 17223 12668 17316 12696
rect 17310 12656 17316 12668
rect 17368 12696 17374 12708
rect 18248 12696 18276 12727
rect 18322 12724 18328 12776
rect 18380 12764 18386 12776
rect 19429 12767 19487 12773
rect 19429 12764 19441 12767
rect 18380 12736 19441 12764
rect 18380 12724 18386 12736
rect 19429 12733 19441 12736
rect 19475 12733 19487 12767
rect 19429 12727 19487 12733
rect 20622 12724 20628 12776
rect 20680 12764 20686 12776
rect 20809 12767 20867 12773
rect 20809 12764 20821 12767
rect 20680 12736 20821 12764
rect 20680 12724 20686 12736
rect 20809 12733 20821 12736
rect 20855 12764 20867 12767
rect 21082 12764 21088 12776
rect 20855 12736 21088 12764
rect 20855 12733 20867 12736
rect 20809 12727 20867 12733
rect 21082 12724 21088 12736
rect 21140 12724 21146 12776
rect 21453 12767 21511 12773
rect 21453 12733 21465 12767
rect 21499 12764 21511 12767
rect 23106 12764 23112 12776
rect 21499 12736 23112 12764
rect 21499 12733 21511 12736
rect 21453 12727 21511 12733
rect 23106 12724 23112 12736
rect 23164 12724 23170 12776
rect 23308 12705 23336 12804
rect 23477 12801 23489 12835
rect 23523 12801 23535 12835
rect 23477 12795 23535 12801
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 23382 12724 23388 12776
rect 23440 12764 23446 12776
rect 23952 12764 23980 12795
rect 27614 12792 27620 12844
rect 27672 12832 27678 12844
rect 29641 12835 29699 12841
rect 29641 12832 29653 12835
rect 27672 12804 29653 12832
rect 27672 12792 27678 12804
rect 29641 12801 29653 12804
rect 29687 12801 29699 12835
rect 29641 12795 29699 12801
rect 23440 12736 23980 12764
rect 23440 12724 23446 12736
rect 17368 12668 18276 12696
rect 18785 12699 18843 12705
rect 17368 12656 17374 12668
rect 18785 12665 18797 12699
rect 18831 12696 18843 12699
rect 19981 12699 20039 12705
rect 19981 12696 19993 12699
rect 18831 12668 19993 12696
rect 18831 12665 18843 12668
rect 18785 12659 18843 12665
rect 19981 12665 19993 12668
rect 20027 12696 20039 12699
rect 23293 12699 23351 12705
rect 20027 12668 22094 12696
rect 20027 12665 20039 12668
rect 19981 12659 20039 12665
rect 5592 12600 5948 12628
rect 5592 12588 5598 12600
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 6362 12628 6368 12640
rect 6144 12600 6368 12628
rect 6144 12588 6150 12600
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 9306 12628 9312 12640
rect 7984 12600 9312 12628
rect 7984 12588 7990 12600
rect 9306 12588 9312 12600
rect 9364 12628 9370 12640
rect 11698 12628 11704 12640
rect 9364 12600 11704 12628
rect 9364 12588 9370 12600
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 12342 12588 12348 12640
rect 12400 12628 12406 12640
rect 21082 12628 21088 12640
rect 12400 12600 21088 12628
rect 12400 12588 12406 12600
rect 21082 12588 21088 12600
rect 21140 12588 21146 12640
rect 22066 12628 22094 12668
rect 23293 12665 23305 12699
rect 23339 12665 23351 12699
rect 23293 12659 23351 12665
rect 28074 12628 28080 12640
rect 22066 12600 28080 12628
rect 28074 12588 28080 12600
rect 28132 12588 28138 12640
rect 29733 12631 29791 12637
rect 29733 12597 29745 12631
rect 29779 12628 29791 12631
rect 31662 12628 31668 12640
rect 29779 12600 31668 12628
rect 29779 12597 29791 12600
rect 29733 12591 29791 12597
rect 31662 12588 31668 12600
rect 31720 12588 31726 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 3163 12427 3221 12433
rect 3163 12393 3175 12427
rect 3209 12424 3221 12427
rect 6546 12424 6552 12436
rect 3209 12396 6408 12424
rect 6507 12396 6552 12424
rect 3209 12393 3221 12396
rect 3163 12387 3221 12393
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 2832 12260 3433 12288
rect 2832 12248 2838 12260
rect 3421 12257 3433 12260
rect 3467 12288 3479 12291
rect 3510 12288 3516 12300
rect 3467 12260 3516 12288
rect 3467 12257 3479 12260
rect 3421 12251 3479 12257
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 3970 12288 3976 12300
rect 3883 12260 3976 12288
rect 3970 12248 3976 12260
rect 4028 12288 4034 12300
rect 5534 12288 5540 12300
rect 4028 12260 5540 12288
rect 4028 12248 4034 12260
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 3050 12152 3056 12164
rect 2714 12124 3056 12152
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 4246 12152 4252 12164
rect 4207 12124 4252 12152
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 4890 12112 4896 12164
rect 4948 12112 4954 12164
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 5997 12155 6055 12161
rect 5997 12152 6009 12155
rect 5684 12124 6009 12152
rect 5684 12112 5690 12124
rect 5997 12121 6009 12124
rect 6043 12121 6055 12155
rect 5997 12115 6055 12121
rect 1673 12087 1731 12093
rect 1673 12053 1685 12087
rect 1719 12084 1731 12087
rect 1854 12084 1860 12096
rect 1719 12056 1860 12084
rect 1719 12053 1731 12056
rect 1673 12047 1731 12053
rect 1854 12044 1860 12056
rect 1912 12084 1918 12096
rect 5902 12084 5908 12096
rect 1912 12056 5908 12084
rect 1912 12044 1918 12056
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 6380 12084 6408 12396
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 6696 12396 13124 12424
rect 6696 12384 6702 12396
rect 11422 12316 11428 12368
rect 11480 12356 11486 12368
rect 12805 12359 12863 12365
rect 12805 12356 12817 12359
rect 11480 12328 12817 12356
rect 11480 12316 11486 12328
rect 12805 12325 12817 12328
rect 12851 12325 12863 12359
rect 13096 12356 13124 12396
rect 13262 12384 13268 12436
rect 13320 12424 13326 12436
rect 13541 12427 13599 12433
rect 13541 12424 13553 12427
rect 13320 12396 13553 12424
rect 13320 12384 13326 12396
rect 13541 12393 13553 12396
rect 13587 12393 13599 12427
rect 15470 12424 15476 12436
rect 15431 12396 15476 12424
rect 13541 12387 13599 12393
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 16758 12424 16764 12436
rect 16347 12396 16764 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 17310 12384 17316 12436
rect 17368 12424 17374 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 17368 12396 17509 12424
rect 17368 12384 17374 12396
rect 17497 12393 17509 12396
rect 17543 12393 17555 12427
rect 18322 12424 18328 12436
rect 18283 12396 18328 12424
rect 17497 12387 17555 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19613 12427 19671 12433
rect 19613 12424 19625 12427
rect 19484 12396 19625 12424
rect 19484 12384 19490 12396
rect 19613 12393 19625 12396
rect 19659 12393 19671 12427
rect 20714 12424 20720 12436
rect 20675 12396 20720 12424
rect 19613 12387 19671 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 20990 12384 20996 12436
rect 21048 12424 21054 12436
rect 21545 12427 21603 12433
rect 21545 12424 21557 12427
rect 21048 12396 21557 12424
rect 21048 12384 21054 12396
rect 21545 12393 21557 12396
rect 21591 12393 21603 12427
rect 21545 12387 21603 12393
rect 14461 12359 14519 12365
rect 13096 12328 13768 12356
rect 12805 12319 12863 12325
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7650 12288 7656 12300
rect 7064 12260 7656 12288
rect 7064 12248 7070 12260
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 10873 12291 10931 12297
rect 10873 12288 10885 12291
rect 8536 12260 10885 12288
rect 8536 12248 8542 12260
rect 10873 12257 10885 12260
rect 10919 12257 10931 12291
rect 10873 12251 10931 12257
rect 11238 12248 11244 12300
rect 11296 12288 11302 12300
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 11296 12260 11345 12288
rect 11296 12248 11302 12260
rect 11333 12257 11345 12260
rect 11379 12288 11391 12291
rect 11698 12288 11704 12300
rect 11379 12260 11704 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 11977 12291 12035 12297
rect 11977 12288 11989 12291
rect 11940 12260 11989 12288
rect 11940 12248 11946 12260
rect 11977 12257 11989 12260
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12268 12260 12756 12288
rect 6914 12180 6920 12232
rect 6972 12180 6978 12232
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 9030 12220 9036 12232
rect 8343 12192 9036 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 9030 12180 9036 12192
rect 9088 12180 9094 12232
rect 11514 12220 11520 12232
rect 11475 12192 11520 12220
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 7742 12112 7748 12164
rect 7800 12152 7806 12164
rect 7800 12124 9260 12152
rect 7800 12112 7806 12124
rect 8386 12084 8392 12096
rect 6380 12056 8392 12084
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 9125 12087 9183 12093
rect 9125 12084 9137 12087
rect 8904 12056 9137 12084
rect 8904 12044 8910 12056
rect 9125 12053 9137 12056
rect 9171 12053 9183 12087
rect 9232 12084 9260 12124
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 9364 12124 9430 12152
rect 9364 12112 9370 12124
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 10597 12155 10655 12161
rect 10597 12152 10609 12155
rect 10560 12124 10609 12152
rect 10560 12112 10566 12124
rect 10597 12121 10609 12124
rect 10643 12121 10655 12155
rect 10597 12115 10655 12121
rect 12268 12084 12296 12260
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 12618 12220 12624 12232
rect 12579 12192 12624 12220
rect 12437 12183 12495 12189
rect 9232 12056 12296 12084
rect 12452 12084 12480 12183
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 12728 12152 12756 12260
rect 13740 12229 13768 12328
rect 14461 12325 14473 12359
rect 14507 12356 14519 12359
rect 15930 12356 15936 12368
rect 14507 12328 15936 12356
rect 14507 12325 14519 12328
rect 14461 12319 14519 12325
rect 15930 12316 15936 12328
rect 15988 12316 15994 12368
rect 20346 12316 20352 12368
rect 20404 12356 20410 12368
rect 21358 12356 21364 12368
rect 20404 12328 21364 12356
rect 20404 12316 20410 12328
rect 21358 12316 21364 12328
rect 21416 12316 21422 12368
rect 23106 12316 23112 12368
rect 23164 12356 23170 12368
rect 23477 12359 23535 12365
rect 23477 12356 23489 12359
rect 23164 12328 23489 12356
rect 23164 12316 23170 12328
rect 23477 12325 23489 12328
rect 23523 12356 23535 12359
rect 30834 12356 30840 12368
rect 23523 12328 30840 12356
rect 23523 12325 23535 12328
rect 23477 12319 23535 12325
rect 30834 12316 30840 12328
rect 30892 12316 30898 12368
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12288 14979 12291
rect 15746 12288 15752 12300
rect 14967 12260 15752 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15746 12248 15752 12260
rect 15804 12248 15810 12300
rect 22002 12288 22008 12300
rect 19720 12260 22008 12288
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 14274 12220 14280 12232
rect 14235 12192 14280 12220
rect 13725 12183 13783 12189
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 15102 12220 15108 12232
rect 15063 12192 15108 12220
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 16482 12220 16488 12232
rect 16443 12192 16488 12220
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 16666 12220 16672 12232
rect 16627 12192 16672 12220
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 17126 12220 17132 12232
rect 17087 12192 17132 12220
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 17310 12220 17316 12232
rect 17271 12192 17316 12220
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18656 12192 18705 12220
rect 18656 12180 18662 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18874 12220 18880 12232
rect 18835 12192 18880 12220
rect 18693 12183 18751 12189
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 19720 12229 19748 12260
rect 22002 12248 22008 12260
rect 22060 12248 22066 12300
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12189 19763 12223
rect 20346 12220 20352 12232
rect 20307 12192 20352 12220
rect 19705 12183 19763 12189
rect 20346 12180 20352 12192
rect 20404 12180 20410 12232
rect 20438 12180 20444 12232
rect 20496 12220 20502 12232
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 20496 12192 20545 12220
rect 20496 12180 20502 12192
rect 20533 12189 20545 12192
rect 20579 12189 20591 12223
rect 21634 12220 21640 12232
rect 21547 12192 21640 12220
rect 20533 12183 20591 12189
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 21652 12152 21680 12180
rect 12728 12124 21680 12152
rect 22373 12155 22431 12161
rect 22373 12121 22385 12155
rect 22419 12152 22431 12155
rect 22925 12155 22983 12161
rect 22925 12152 22937 12155
rect 22419 12124 22937 12152
rect 22419 12121 22431 12124
rect 22373 12115 22431 12121
rect 22925 12121 22937 12124
rect 22971 12121 22983 12155
rect 22925 12115 22983 12121
rect 23017 12155 23075 12161
rect 23017 12121 23029 12155
rect 23063 12152 23075 12155
rect 23382 12152 23388 12164
rect 23063 12124 23388 12152
rect 23063 12121 23075 12124
rect 23017 12115 23075 12121
rect 23382 12112 23388 12124
rect 23440 12112 23446 12164
rect 12894 12084 12900 12096
rect 12452 12056 12900 12084
rect 9125 12047 9183 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 13630 12044 13636 12096
rect 13688 12084 13694 12096
rect 14550 12084 14556 12096
rect 13688 12056 14556 12084
rect 13688 12044 13694 12056
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 5905 11883 5963 11889
rect 2464 11852 5120 11880
rect 2464 11840 2470 11852
rect 2314 11812 2320 11824
rect 2275 11784 2320 11812
rect 2314 11772 2320 11784
rect 2372 11772 2378 11824
rect 4062 11812 4068 11824
rect 3542 11784 4068 11812
rect 4062 11772 4068 11784
rect 4120 11772 4126 11824
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4764 11716 4813 11744
rect 4764 11704 4770 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 5092 11744 5120 11852
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 5994 11880 6000 11892
rect 5951 11852 6000 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 6825 11883 6883 11889
rect 6825 11849 6837 11883
rect 6871 11880 6883 11883
rect 12345 11883 12403 11889
rect 6871 11852 11928 11880
rect 6871 11849 6883 11852
rect 6825 11843 6883 11849
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 7466 11812 7472 11824
rect 5500 11784 7472 11812
rect 5500 11772 5506 11784
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 8849 11815 8907 11821
rect 8849 11781 8861 11815
rect 8895 11812 8907 11815
rect 10318 11812 10324 11824
rect 8895 11784 10324 11812
rect 8895 11781 8907 11784
rect 8849 11775 8907 11781
rect 10318 11772 10324 11784
rect 10376 11772 10382 11824
rect 5534 11744 5540 11756
rect 5092 11716 5540 11744
rect 4801 11707 4859 11713
rect 5534 11704 5540 11716
rect 5592 11744 5598 11756
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 5592 11716 5825 11744
rect 5592 11704 5598 11716
rect 5813 11713 5825 11716
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 5960 11716 6745 11744
rect 5960 11704 5966 11716
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 7742 11704 7748 11756
rect 7800 11704 7806 11756
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9180 11716 9225 11744
rect 9180 11704 9186 11716
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 9824 11716 10609 11744
rect 9824 11704 9830 11716
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 11900 11753 11928 11852
rect 12345 11849 12357 11883
rect 12391 11880 12403 11883
rect 13170 11880 13176 11892
rect 12391 11852 13176 11880
rect 12391 11849 12403 11852
rect 12345 11843 12403 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 15010 11880 15016 11892
rect 14507 11852 15016 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 15010 11840 15016 11852
rect 15068 11840 15074 11892
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15657 11883 15715 11889
rect 15657 11880 15669 11883
rect 15528 11852 15669 11880
rect 15528 11840 15534 11852
rect 15657 11849 15669 11852
rect 15703 11849 15715 11883
rect 15657 11843 15715 11849
rect 16206 11840 16212 11892
rect 16264 11880 16270 11892
rect 16301 11883 16359 11889
rect 16301 11880 16313 11883
rect 16264 11852 16313 11880
rect 16264 11840 16270 11852
rect 16301 11849 16313 11852
rect 16347 11849 16359 11883
rect 16301 11843 16359 11849
rect 17862 11840 17868 11892
rect 17920 11880 17926 11892
rect 17957 11883 18015 11889
rect 17957 11880 17969 11883
rect 17920 11852 17969 11880
rect 17920 11840 17926 11852
rect 17957 11849 17969 11852
rect 18003 11849 18015 11883
rect 17957 11843 18015 11849
rect 18506 11840 18512 11892
rect 18564 11880 18570 11892
rect 18601 11883 18659 11889
rect 18601 11880 18613 11883
rect 18564 11852 18613 11880
rect 18564 11840 18570 11852
rect 18601 11849 18613 11852
rect 18647 11849 18659 11883
rect 18601 11843 18659 11849
rect 19705 11883 19763 11889
rect 19705 11849 19717 11883
rect 19751 11880 19763 11883
rect 20162 11880 20168 11892
rect 19751 11852 20168 11880
rect 19751 11849 19763 11852
rect 19705 11843 19763 11849
rect 20162 11840 20168 11852
rect 20220 11840 20226 11892
rect 20438 11880 20444 11892
rect 20399 11852 20444 11880
rect 20438 11840 20444 11852
rect 20496 11840 20502 11892
rect 20898 11840 20904 11892
rect 20956 11880 20962 11892
rect 21085 11883 21143 11889
rect 21085 11880 21097 11883
rect 20956 11852 21097 11880
rect 20956 11840 20962 11852
rect 21085 11849 21097 11852
rect 21131 11849 21143 11883
rect 23382 11880 23388 11892
rect 23343 11852 23388 11880
rect 21085 11843 21143 11849
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 36906 11840 36912 11892
rect 36964 11880 36970 11892
rect 38105 11883 38163 11889
rect 38105 11880 38117 11883
rect 36964 11852 38117 11880
rect 36964 11840 36970 11852
rect 38105 11849 38117 11852
rect 38151 11849 38163 11883
rect 38105 11843 38163 11849
rect 17405 11815 17463 11821
rect 11992 11784 13676 11812
rect 11885 11747 11943 11753
rect 10928 11716 11836 11744
rect 10928 11704 10934 11716
rect 2038 11676 2044 11688
rect 1999 11648 2044 11676
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 4154 11676 4160 11688
rect 4111 11648 4160 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 3602 11568 3608 11620
rect 3660 11608 3666 11620
rect 4080 11608 4108 11639
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 4816 11648 9076 11676
rect 4706 11608 4712 11620
rect 3660 11580 4712 11608
rect 3660 11568 3666 11580
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 1670 11500 1676 11552
rect 1728 11540 1734 11552
rect 4816 11540 4844 11648
rect 4893 11611 4951 11617
rect 4893 11577 4905 11611
rect 4939 11608 4951 11611
rect 7834 11608 7840 11620
rect 4939 11580 7840 11608
rect 4939 11577 4951 11580
rect 4893 11571 4951 11577
rect 7834 11568 7840 11580
rect 7892 11568 7898 11620
rect 9048 11608 9076 11648
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 10008 11648 10425 11676
rect 10008 11636 10014 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 10686 11636 10692 11688
rect 10744 11676 10750 11688
rect 10744 11648 11008 11676
rect 10744 11636 10750 11648
rect 10980 11608 11008 11648
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11112 11648 11713 11676
rect 11112 11636 11118 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11808 11676 11836 11716
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 11992 11676 12020 11784
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 13648 11753 13676 11784
rect 17405 11781 17417 11815
rect 17451 11812 17463 11815
rect 18138 11812 18144 11824
rect 17451 11784 18144 11812
rect 17451 11781 17463 11784
rect 17405 11775 17463 11781
rect 18138 11772 18144 11784
rect 18196 11772 18202 11824
rect 36814 11812 36820 11824
rect 18248 11784 36820 11812
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 12492 11716 12817 11744
rect 12492 11704 12498 11716
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 17126 11704 17132 11756
rect 17184 11744 17190 11756
rect 17313 11747 17371 11753
rect 17313 11744 17325 11747
rect 17184 11716 17325 11744
rect 17184 11704 17190 11716
rect 17313 11713 17325 11716
rect 17359 11713 17371 11747
rect 17313 11707 17371 11713
rect 17586 11704 17592 11756
rect 17644 11744 17650 11756
rect 18248 11744 18276 11784
rect 36814 11772 36820 11784
rect 36872 11772 36878 11824
rect 17644 11716 18276 11744
rect 17644 11704 17650 11716
rect 18690 11704 18696 11756
rect 18748 11744 18754 11756
rect 18785 11747 18843 11753
rect 18785 11744 18797 11747
rect 18748 11716 18797 11744
rect 18748 11704 18754 11716
rect 18785 11713 18797 11716
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11713 19671 11747
rect 19613 11707 19671 11713
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11744 20315 11747
rect 20438 11744 20444 11756
rect 20303 11716 20444 11744
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 15010 11676 15016 11688
rect 11808 11648 12020 11676
rect 14971 11648 15016 11676
rect 11701 11639 11759 11645
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 15194 11676 15200 11688
rect 15155 11648 15200 11676
rect 15194 11636 15200 11648
rect 15252 11636 15258 11688
rect 11146 11608 11152 11620
rect 9048 11580 10916 11608
rect 10980 11580 11152 11608
rect 10888 11552 10916 11580
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 12897 11611 12955 11617
rect 12897 11577 12909 11611
rect 12943 11608 12955 11611
rect 14274 11608 14280 11620
rect 12943 11580 14280 11608
rect 12943 11577 12955 11580
rect 12897 11571 12955 11577
rect 14274 11568 14280 11580
rect 14332 11568 14338 11620
rect 14734 11568 14740 11620
rect 14792 11608 14798 11620
rect 19628 11608 19656 11707
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 21082 11704 21088 11756
rect 21140 11744 21146 11756
rect 21177 11747 21235 11753
rect 21177 11744 21189 11747
rect 21140 11716 21189 11744
rect 21140 11704 21146 11716
rect 21177 11713 21189 11716
rect 21223 11744 21235 11747
rect 22097 11747 22155 11753
rect 22097 11744 22109 11747
rect 21223 11716 22109 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 22097 11713 22109 11716
rect 22143 11713 22155 11747
rect 22738 11744 22744 11756
rect 22699 11716 22744 11744
rect 22097 11707 22155 11713
rect 22738 11704 22744 11716
rect 22796 11744 22802 11756
rect 23290 11744 23296 11756
rect 22796 11716 23296 11744
rect 22796 11704 22802 11716
rect 23290 11704 23296 11716
rect 23348 11704 23354 11756
rect 23569 11747 23627 11753
rect 23569 11713 23581 11747
rect 23615 11713 23627 11747
rect 27430 11744 27436 11756
rect 27391 11716 27436 11744
rect 23569 11707 23627 11713
rect 23584 11676 23612 11707
rect 27430 11704 27436 11716
rect 27488 11704 27494 11756
rect 31662 11704 31668 11756
rect 31720 11744 31726 11756
rect 34149 11747 34207 11753
rect 34149 11744 34161 11747
rect 31720 11716 34161 11744
rect 31720 11704 31726 11716
rect 34149 11713 34161 11716
rect 34195 11713 34207 11747
rect 38286 11744 38292 11756
rect 38247 11716 38292 11744
rect 34149 11707 34207 11713
rect 38286 11704 38292 11716
rect 38344 11704 38350 11756
rect 22296 11648 23612 11676
rect 20254 11608 20260 11620
rect 14792 11580 20260 11608
rect 14792 11568 14798 11580
rect 20254 11568 20260 11580
rect 20312 11568 20318 11620
rect 22296 11617 22324 11648
rect 22281 11611 22339 11617
rect 22281 11577 22293 11611
rect 22327 11577 22339 11611
rect 22281 11571 22339 11577
rect 22925 11611 22983 11617
rect 22925 11577 22937 11611
rect 22971 11608 22983 11611
rect 23658 11608 23664 11620
rect 22971 11580 23664 11608
rect 22971 11577 22983 11580
rect 22925 11571 22983 11577
rect 23658 11568 23664 11580
rect 23716 11568 23722 11620
rect 1728 11512 4844 11540
rect 7377 11543 7435 11549
rect 1728 11500 1734 11512
rect 7377 11509 7389 11543
rect 7423 11540 7435 11543
rect 8294 11540 8300 11552
rect 7423 11512 8300 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 10410 11540 10416 11552
rect 8444 11512 10416 11540
rect 8444 11500 8450 11512
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 10744 11512 10793 11540
rect 10744 11500 10750 11512
rect 10781 11509 10793 11512
rect 10827 11509 10839 11543
rect 10781 11503 10839 11509
rect 10870 11500 10876 11552
rect 10928 11500 10934 11552
rect 13817 11543 13875 11549
rect 13817 11509 13829 11543
rect 13863 11540 13875 11543
rect 14366 11540 14372 11552
rect 13863 11512 14372 11540
rect 13863 11509 13875 11512
rect 13817 11503 13875 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 27525 11543 27583 11549
rect 27525 11509 27537 11543
rect 27571 11540 27583 11543
rect 32858 11540 32864 11552
rect 27571 11512 32864 11540
rect 27571 11509 27583 11512
rect 27525 11503 27583 11509
rect 32858 11500 32864 11512
rect 32916 11500 32922 11552
rect 34333 11543 34391 11549
rect 34333 11509 34345 11543
rect 34379 11540 34391 11543
rect 35342 11540 35348 11552
rect 34379 11512 35348 11540
rect 34379 11509 34391 11512
rect 34333 11503 34391 11509
rect 35342 11500 35348 11512
rect 35400 11500 35406 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 3510 11336 3516 11348
rect 3108 11308 3516 11336
rect 3108 11296 3114 11308
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 4249 11339 4307 11345
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 9769 11339 9827 11345
rect 4295 11308 9720 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 9692 11268 9720 11308
rect 9769 11305 9781 11339
rect 9815 11336 9827 11339
rect 10594 11336 10600 11348
rect 9815 11308 10600 11336
rect 9815 11305 9827 11308
rect 9769 11299 9827 11305
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 10965 11339 11023 11345
rect 10965 11305 10977 11339
rect 11011 11336 11023 11339
rect 11146 11336 11152 11348
rect 11011 11308 11152 11336
rect 11011 11305 11023 11308
rect 10965 11299 11023 11305
rect 11146 11296 11152 11308
rect 11204 11296 11210 11348
rect 11790 11336 11796 11348
rect 11751 11308 11796 11336
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 13173 11339 13231 11345
rect 13173 11305 13185 11339
rect 13219 11336 13231 11339
rect 13998 11336 14004 11348
rect 13219 11308 14004 11336
rect 13219 11305 13231 11308
rect 13173 11299 13231 11305
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14553 11339 14611 11345
rect 14553 11305 14565 11339
rect 14599 11336 14611 11339
rect 15286 11336 15292 11348
rect 14599 11308 15292 11336
rect 14599 11305 14611 11308
rect 14553 11299 14611 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 15378 11296 15384 11348
rect 15436 11336 15442 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 15436 11308 15485 11336
rect 15436 11296 15442 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 16942 11336 16948 11348
rect 16715 11308 16948 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17865 11339 17923 11345
rect 17865 11305 17877 11339
rect 17911 11336 17923 11339
rect 18046 11336 18052 11348
rect 17911 11308 18052 11336
rect 17911 11305 17923 11308
rect 17865 11299 17923 11305
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 19484 11308 19625 11336
rect 19484 11296 19490 11308
rect 19613 11305 19625 11308
rect 19659 11305 19671 11339
rect 20438 11336 20444 11348
rect 20399 11308 20444 11336
rect 19613 11299 19671 11305
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 11422 11268 11428 11280
rect 9416 11240 9628 11268
rect 9692 11240 11428 11268
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 2832 11172 6009 11200
rect 2832 11160 2838 11172
rect 5997 11169 6009 11172
rect 6043 11169 6055 11203
rect 5997 11163 6055 11169
rect 6270 11160 6276 11212
rect 6328 11200 6334 11212
rect 6825 11203 6883 11209
rect 6825 11200 6837 11203
rect 6328 11172 6837 11200
rect 6328 11160 6334 11172
rect 6825 11169 6837 11172
rect 6871 11200 6883 11203
rect 7650 11200 7656 11212
rect 6871 11172 7656 11200
rect 6871 11169 6883 11172
rect 6825 11163 6883 11169
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 8294 11200 8300 11212
rect 8255 11172 8300 11200
rect 8294 11160 8300 11172
rect 8352 11200 8358 11212
rect 9416 11200 9444 11240
rect 8352 11172 9444 11200
rect 9600 11200 9628 11240
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 12437 11271 12495 11277
rect 12437 11237 12449 11271
rect 12483 11268 12495 11271
rect 13906 11268 13912 11280
rect 12483 11240 13912 11268
rect 12483 11237 12495 11240
rect 12437 11231 12495 11237
rect 13906 11228 13912 11240
rect 13964 11228 13970 11280
rect 17313 11271 17371 11277
rect 17313 11237 17325 11271
rect 17359 11268 17371 11271
rect 19058 11268 19064 11280
rect 17359 11240 19064 11268
rect 17359 11237 17371 11240
rect 17313 11231 17371 11237
rect 19058 11228 19064 11240
rect 19116 11228 19122 11280
rect 17862 11200 17868 11212
rect 9600 11172 17868 11200
rect 8352 11160 8358 11172
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 3970 11132 3976 11144
rect 3467 11104 3976 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 9398 11132 9404 11144
rect 8628 11104 9404 11132
rect 8628 11092 8634 11104
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 9490 11092 9496 11144
rect 9548 11132 9554 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9548 11104 9689 11132
rect 9548 11092 9554 11104
rect 9677 11101 9689 11104
rect 9723 11132 9735 11135
rect 10226 11132 10232 11144
rect 9723 11104 10232 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 10505 11135 10563 11141
rect 10376 11104 10421 11132
rect 10376 11092 10382 11104
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 10505 11095 10563 11101
rect 2682 11024 2688 11076
rect 2740 11024 2746 11076
rect 3145 11067 3203 11073
rect 3145 11033 3157 11067
rect 3191 11064 3203 11067
rect 3786 11064 3792 11076
rect 3191 11036 3792 11064
rect 3191 11033 3203 11036
rect 3145 11027 3203 11033
rect 3786 11024 3792 11036
rect 3844 11024 3850 11076
rect 3988 11064 4016 11092
rect 3988 11036 4384 11064
rect 4356 10996 4384 11036
rect 5166 11024 5172 11076
rect 5224 11024 5230 11076
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 5721 11067 5779 11073
rect 5721 11064 5733 11067
rect 5684 11036 5733 11064
rect 5684 11024 5690 11036
rect 5721 11033 5733 11036
rect 5767 11064 5779 11067
rect 5767 11036 6408 11064
rect 5767 11033 5779 11036
rect 5721 11027 5779 11033
rect 4706 10996 4712 11008
rect 4356 10968 4712 10996
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 6380 10996 6408 11036
rect 6454 11024 6460 11076
rect 6512 11064 6518 11076
rect 8662 11064 8668 11076
rect 6512 11036 7130 11064
rect 7944 11036 8668 11064
rect 6512 11024 6518 11036
rect 7944 10996 7972 11036
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 8846 11024 8852 11076
rect 8904 11064 8910 11076
rect 8904 11036 9674 11064
rect 8904 11024 8910 11036
rect 6380 10968 7972 10996
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 9490 10996 9496 11008
rect 8536 10968 9496 10996
rect 8536 10956 8542 10968
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 9646 10996 9674 11036
rect 10042 11024 10048 11076
rect 10100 11064 10106 11076
rect 10520 11064 10548 11095
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12342 11132 12348 11144
rect 12303 11104 12348 11132
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12986 11132 12992 11144
rect 12947 11104 12992 11132
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 14366 11132 14372 11144
rect 14327 11104 14372 11132
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 16776 11141 16804 11172
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 15381 11135 15439 11141
rect 15381 11132 15393 11135
rect 14608 11104 15393 11132
rect 14608 11092 14614 11104
rect 15381 11101 15393 11104
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 16761 11135 16819 11141
rect 16761 11101 16773 11135
rect 16807 11101 16819 11135
rect 16761 11095 16819 11101
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 17221 11135 17279 11141
rect 17221 11132 17233 11135
rect 17000 11104 17233 11132
rect 17000 11092 17006 11104
rect 17221 11101 17233 11104
rect 17267 11101 17279 11135
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 17221 11095 17279 11101
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18509 11135 18567 11141
rect 18509 11101 18521 11135
rect 18555 11101 18567 11135
rect 18509 11095 18567 11101
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11132 19855 11135
rect 19978 11132 19984 11144
rect 19843 11104 19984 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 10100 11036 10548 11064
rect 10100 11024 10106 11036
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 17126 11064 17132 11076
rect 10928 11036 17132 11064
rect 10928 11024 10934 11036
rect 17126 11024 17132 11036
rect 17184 11064 17190 11076
rect 18524 11064 18552 11095
rect 19978 11092 19984 11104
rect 20036 11092 20042 11144
rect 20254 11132 20260 11144
rect 20215 11104 20260 11132
rect 20254 11092 20260 11104
rect 20312 11092 20318 11144
rect 17184 11036 18552 11064
rect 17184 11024 17190 11036
rect 10962 10996 10968 11008
rect 9646 10968 10968 10996
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 12066 10996 12072 11008
rect 11204 10968 12072 10996
rect 11204 10956 11210 10968
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 2774 10792 2780 10804
rect 1688 10764 2780 10792
rect 1688 10665 1716 10764
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 2866 10752 2872 10804
rect 2924 10792 2930 10804
rect 3421 10795 3479 10801
rect 3421 10792 3433 10795
rect 2924 10764 3433 10792
rect 2924 10752 2930 10764
rect 3421 10761 3433 10764
rect 3467 10761 3479 10795
rect 6638 10792 6644 10804
rect 3421 10755 3479 10761
rect 4448 10764 6500 10792
rect 6599 10764 6644 10792
rect 1946 10724 1952 10736
rect 1907 10696 1952 10724
rect 1946 10684 1952 10696
rect 2004 10684 2010 10736
rect 4448 10724 4476 10764
rect 3174 10696 4476 10724
rect 5721 10727 5779 10733
rect 5721 10693 5733 10727
rect 5767 10724 5779 10727
rect 6270 10724 6276 10736
rect 5767 10696 6276 10724
rect 5767 10693 5779 10696
rect 5721 10687 5779 10693
rect 6270 10684 6276 10696
rect 6328 10684 6334 10736
rect 6472 10724 6500 10764
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 6822 10752 6828 10804
rect 6880 10792 6886 10804
rect 7653 10795 7711 10801
rect 7653 10792 7665 10795
rect 6880 10764 7665 10792
rect 6880 10752 6886 10764
rect 7653 10761 7665 10764
rect 7699 10761 7711 10795
rect 10137 10795 10195 10801
rect 7653 10755 7711 10761
rect 7852 10764 10088 10792
rect 7282 10724 7288 10736
rect 6472 10696 7288 10724
rect 7282 10684 7288 10696
rect 7340 10684 7346 10736
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 4632 10520 4660 10642
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6052 10628 6097 10656
rect 6288 10628 6561 10656
rect 6052 10616 6058 10628
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5316 10560 5948 10588
rect 5316 10548 5322 10560
rect 3344 10492 4660 10520
rect 5920 10520 5948 10560
rect 6288 10520 6316 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 7852 10656 7880 10764
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 9674 10724 9680 10736
rect 9171 10696 9680 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 10060 10724 10088 10764
rect 10137 10761 10149 10795
rect 10183 10792 10195 10795
rect 11514 10792 11520 10804
rect 10183 10764 11520 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 11882 10752 11888 10804
rect 11940 10792 11946 10804
rect 12805 10795 12863 10801
rect 11940 10764 12572 10792
rect 11940 10752 11946 10764
rect 10689 10727 10747 10733
rect 10060 10696 10640 10724
rect 6696 10628 7880 10656
rect 6696 10616 6702 10628
rect 8018 10616 8024 10668
rect 8076 10616 8082 10668
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9953 10659 10011 10665
rect 9456 10628 9501 10656
rect 9456 10616 9462 10628
rect 9953 10625 9965 10659
rect 9999 10656 10011 10659
rect 10502 10656 10508 10668
rect 9999 10628 10508 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 10612 10665 10640 10696
rect 10689 10693 10701 10727
rect 10735 10724 10747 10727
rect 11146 10724 11152 10736
rect 10735 10696 11152 10724
rect 10735 10693 10747 10696
rect 10689 10687 10747 10693
rect 11146 10684 11152 10696
rect 11204 10684 11210 10736
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 11296 10696 11652 10724
rect 11296 10684 11302 10696
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10656 10655 10659
rect 11514 10656 11520 10668
rect 10643 10628 11520 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 11624 10656 11652 10696
rect 11790 10684 11796 10736
rect 11848 10724 11854 10736
rect 12544 10724 12572 10764
rect 12805 10761 12817 10795
rect 12851 10792 12863 10795
rect 12986 10792 12992 10804
rect 12851 10764 12992 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 13541 10795 13599 10801
rect 13541 10761 13553 10795
rect 13587 10792 13599 10795
rect 14090 10792 14096 10804
rect 13587 10764 14096 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 14826 10792 14832 10804
rect 14787 10764 14832 10792
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 15657 10795 15715 10801
rect 15657 10761 15669 10795
rect 15703 10792 15715 10795
rect 16114 10792 16120 10804
rect 15703 10764 16120 10792
rect 15703 10761 15715 10764
rect 15657 10755 15715 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 16301 10795 16359 10801
rect 16301 10761 16313 10795
rect 16347 10792 16359 10795
rect 16574 10792 16580 10804
rect 16347 10764 16580 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 17313 10795 17371 10801
rect 17313 10761 17325 10795
rect 17359 10792 17371 10795
rect 17494 10792 17500 10804
rect 17359 10764 17500 10792
rect 17359 10761 17371 10764
rect 17313 10755 17371 10761
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 18046 10792 18052 10804
rect 18007 10764 18052 10792
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 18874 10792 18880 10804
rect 18835 10764 18880 10792
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 19705 10795 19763 10801
rect 19705 10761 19717 10795
rect 19751 10792 19763 10795
rect 19978 10792 19984 10804
rect 19751 10764 19984 10792
rect 19751 10761 19763 10764
rect 19705 10755 19763 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 15930 10724 15936 10736
rect 11848 10696 12434 10724
rect 12544 10696 15936 10724
rect 11848 10684 11854 10696
rect 11882 10656 11888 10668
rect 11624 10628 11888 10656
rect 11882 10616 11888 10628
rect 11940 10656 11946 10668
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 11940 10628 11989 10656
rect 11940 10616 11946 10628
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 12406 10656 12434 10696
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 12406 10628 12633 10656
rect 11977 10619 12035 10625
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10656 13507 10659
rect 13906 10656 13912 10668
rect 13495 10628 13912 10656
rect 13495 10625 13507 10628
rect 13449 10619 13507 10625
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 14274 10656 14280 10668
rect 14235 10628 14280 10656
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14608 10628 14933 10656
rect 14608 10616 14614 10628
rect 14921 10625 14933 10628
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 16117 10659 16175 10665
rect 16117 10625 16129 10659
rect 16163 10656 16175 10659
rect 16390 10656 16396 10668
rect 16163 10628 16396 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 16390 10616 16396 10628
rect 16448 10616 16454 10668
rect 17221 10659 17279 10665
rect 17221 10625 17233 10659
rect 17267 10625 17279 10659
rect 17862 10656 17868 10668
rect 17823 10628 17868 10656
rect 17221 10619 17279 10625
rect 17236 10588 17264 10619
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 19518 10656 19524 10668
rect 19479 10628 19524 10656
rect 19518 10616 19524 10628
rect 19576 10616 19582 10668
rect 20349 10659 20407 10665
rect 20349 10625 20361 10659
rect 20395 10625 20407 10659
rect 20349 10619 20407 10625
rect 17678 10588 17684 10600
rect 5920 10492 6316 10520
rect 9324 10560 17684 10588
rect 2406 10412 2412 10464
rect 2464 10452 2470 10464
rect 3344 10452 3372 10492
rect 2464 10424 3372 10452
rect 4249 10455 4307 10461
rect 2464 10412 2470 10424
rect 4249 10421 4261 10455
rect 4295 10452 4307 10455
rect 5626 10452 5632 10464
rect 4295 10424 5632 10452
rect 4295 10421 4307 10424
rect 4249 10415 4307 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 6086 10412 6092 10464
rect 6144 10452 6150 10464
rect 9324 10452 9352 10560
rect 17678 10548 17684 10560
rect 17736 10588 17742 10600
rect 20364 10588 20392 10619
rect 28074 10616 28080 10668
rect 28132 10656 28138 10668
rect 30009 10659 30067 10665
rect 30009 10656 30021 10659
rect 28132 10628 30021 10656
rect 28132 10616 28138 10628
rect 30009 10625 30021 10628
rect 30055 10625 30067 10659
rect 30009 10619 30067 10625
rect 35342 10616 35348 10668
rect 35400 10656 35406 10668
rect 38013 10659 38071 10665
rect 38013 10656 38025 10659
rect 35400 10628 38025 10656
rect 35400 10616 35406 10628
rect 38013 10625 38025 10628
rect 38059 10625 38071 10659
rect 38013 10619 38071 10625
rect 17736 10560 20392 10588
rect 17736 10548 17742 10560
rect 10410 10480 10416 10532
rect 10468 10520 10474 10532
rect 11790 10520 11796 10532
rect 10468 10492 11796 10520
rect 10468 10480 10474 10492
rect 11790 10480 11796 10492
rect 11848 10480 11854 10532
rect 14093 10523 14151 10529
rect 14093 10520 14105 10523
rect 12084 10492 14105 10520
rect 6144 10424 9352 10452
rect 6144 10412 6150 10424
rect 9490 10412 9496 10464
rect 9548 10452 9554 10464
rect 12084 10452 12112 10492
rect 14093 10489 14105 10492
rect 14139 10489 14151 10523
rect 14093 10483 14151 10489
rect 9548 10424 12112 10452
rect 12161 10455 12219 10461
rect 9548 10412 9554 10424
rect 12161 10421 12173 10455
rect 12207 10452 12219 10455
rect 13262 10452 13268 10464
rect 12207 10424 13268 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 13262 10412 13268 10424
rect 13320 10412 13326 10464
rect 18874 10412 18880 10464
rect 18932 10452 18938 10464
rect 20165 10455 20223 10461
rect 20165 10452 20177 10455
rect 18932 10424 20177 10452
rect 18932 10412 18938 10424
rect 20165 10421 20177 10424
rect 20211 10421 20223 10455
rect 30098 10452 30104 10464
rect 30059 10424 30104 10452
rect 20165 10415 20223 10421
rect 30098 10412 30104 10424
rect 30156 10412 30162 10464
rect 38194 10452 38200 10464
rect 38155 10424 38200 10452
rect 38194 10412 38200 10424
rect 38252 10412 38258 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 6086 10248 6092 10260
rect 1544 10220 6092 10248
rect 1544 10208 1550 10220
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 6178 10208 6184 10260
rect 6236 10248 6242 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6236 10220 6837 10248
rect 6236 10208 6242 10220
rect 6825 10217 6837 10220
rect 6871 10217 6883 10251
rect 6825 10211 6883 10217
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8309 10251 8367 10257
rect 8309 10248 8321 10251
rect 8168 10220 8321 10248
rect 8168 10208 8174 10220
rect 8309 10217 8321 10220
rect 8355 10248 8367 10251
rect 9674 10248 9680 10260
rect 8355 10220 9680 10248
rect 8355 10217 8367 10220
rect 8309 10211 8367 10217
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10502 10248 10508 10260
rect 9968 10220 10180 10248
rect 10463 10220 10508 10248
rect 4065 10183 4123 10189
rect 4065 10149 4077 10183
rect 4111 10180 4123 10183
rect 6362 10180 6368 10192
rect 4111 10152 4752 10180
rect 6323 10152 6368 10180
rect 4111 10149 4123 10152
rect 4065 10143 4123 10149
rect 2038 10072 2044 10124
rect 2096 10112 2102 10124
rect 4614 10112 4620 10124
rect 2096 10084 2774 10112
rect 4575 10084 4620 10112
rect 2096 10072 2102 10084
rect 2746 10044 2774 10084
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 4724 10112 4752 10152
rect 6362 10140 6368 10152
rect 6420 10180 6426 10192
rect 6638 10180 6644 10192
rect 6420 10152 6644 10180
rect 6420 10140 6426 10152
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 9309 10183 9367 10189
rect 9309 10149 9321 10183
rect 9355 10180 9367 10183
rect 9968 10180 9996 10220
rect 9355 10152 9996 10180
rect 10152 10180 10180 10220
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 11330 10248 11336 10260
rect 11291 10220 11336 10248
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 11977 10251 12035 10257
rect 11977 10217 11989 10251
rect 12023 10248 12035 10251
rect 12250 10248 12256 10260
rect 12023 10220 12256 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 13078 10248 13084 10260
rect 13039 10220 13084 10248
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14240 10220 14749 10248
rect 14240 10208 14246 10220
rect 14737 10217 14749 10220
rect 14783 10217 14795 10251
rect 14737 10211 14795 10217
rect 15749 10251 15807 10257
rect 15749 10217 15761 10251
rect 15795 10248 15807 10251
rect 15838 10248 15844 10260
rect 15795 10220 15844 10248
rect 15795 10217 15807 10220
rect 15749 10211 15807 10217
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 16390 10248 16396 10260
rect 16351 10220 16396 10248
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 17221 10251 17279 10257
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 17310 10248 17316 10260
rect 17267 10220 17316 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17954 10248 17960 10260
rect 17915 10220 17960 10248
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 18693 10251 18751 10257
rect 18693 10248 18705 10251
rect 18656 10220 18705 10248
rect 18656 10208 18662 10220
rect 18693 10217 18705 10220
rect 18739 10217 18751 10251
rect 18693 10211 18751 10217
rect 19242 10208 19248 10260
rect 19300 10248 19306 10260
rect 19521 10251 19579 10257
rect 19521 10248 19533 10251
rect 19300 10220 19533 10248
rect 19300 10208 19306 10220
rect 19521 10217 19533 10220
rect 19567 10217 19579 10251
rect 19521 10211 19579 10217
rect 21910 10208 21916 10260
rect 21968 10248 21974 10260
rect 25317 10251 25375 10257
rect 25317 10248 25329 10251
rect 21968 10220 25329 10248
rect 21968 10208 21974 10220
rect 25317 10217 25329 10220
rect 25363 10217 25375 10251
rect 25317 10211 25375 10217
rect 12618 10180 12624 10192
rect 10152 10152 12624 10180
rect 9355 10149 9367 10152
rect 9309 10143 9367 10149
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 17770 10140 17776 10192
rect 17828 10180 17834 10192
rect 20165 10183 20223 10189
rect 20165 10180 20177 10183
rect 17828 10152 20177 10180
rect 17828 10140 17834 10152
rect 20165 10149 20177 10152
rect 20211 10149 20223 10183
rect 20165 10143 20223 10149
rect 7006 10112 7012 10124
rect 4724 10084 7012 10112
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 8570 10112 8576 10124
rect 8352 10084 8576 10112
rect 8352 10072 8358 10084
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 10468 10084 11192 10112
rect 10468 10072 10474 10084
rect 3973 10047 4031 10053
rect 3973 10044 3985 10047
rect 2746 10016 3985 10044
rect 3973 10013 3985 10016
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10044 9275 10047
rect 10045 10047 10103 10053
rect 9263 10038 9674 10044
rect 10045 10038 10057 10047
rect 9263 10016 10057 10038
rect 9263 10013 9275 10016
rect 9217 10007 9275 10013
rect 9646 10013 10057 10016
rect 10091 10013 10103 10047
rect 9646 10010 10103 10013
rect 10045 10007 10103 10010
rect 3234 9936 3240 9988
rect 3292 9976 3298 9988
rect 3418 9976 3424 9988
rect 3292 9948 3424 9976
rect 3292 9936 3298 9948
rect 3418 9936 3424 9948
rect 3476 9936 3482 9988
rect 3602 9936 3608 9988
rect 3660 9976 3666 9988
rect 4893 9979 4951 9985
rect 4893 9976 4905 9979
rect 3660 9948 4905 9976
rect 3660 9936 3666 9948
rect 4893 9945 4905 9948
rect 4939 9945 4951 9979
rect 6118 9948 6960 9976
rect 4893 9939 4951 9945
rect 2130 9908 2136 9920
rect 2091 9880 2136 9908
rect 2130 9868 2136 9880
rect 2188 9868 2194 9920
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 5258 9908 5264 9920
rect 3844 9880 5264 9908
rect 3844 9868 3850 9880
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 6932 9908 6960 9948
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 7064 9948 7130 9976
rect 7064 9936 7070 9948
rect 8202 9936 8208 9988
rect 8260 9976 8266 9988
rect 10060 9976 10088 10007
rect 10226 10004 10232 10056
rect 10284 10044 10290 10056
rect 11164 10053 11192 10084
rect 11238 10072 11244 10124
rect 11296 10112 11302 10124
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 11296 10084 12541 10112
rect 11296 10072 11302 10084
rect 12529 10081 12541 10084
rect 12575 10081 12587 10115
rect 16850 10112 16856 10124
rect 12529 10075 12587 10081
rect 15580 10084 16856 10112
rect 10689 10047 10747 10053
rect 10689 10044 10701 10047
rect 10284 10016 10701 10044
rect 10284 10004 10290 10016
rect 10689 10013 10701 10016
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10013 11207 10047
rect 11790 10044 11796 10056
rect 11751 10016 11796 10044
rect 11149 10007 11207 10013
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 12802 10044 12808 10056
rect 12667 10016 12808 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13262 10044 13268 10056
rect 13223 10016 13268 10044
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 14918 10044 14924 10056
rect 14879 10016 14924 10044
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 15580 10053 15608 10084
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17034 10072 17040 10124
rect 17092 10112 17098 10124
rect 17092 10084 22094 10112
rect 17092 10072 17098 10084
rect 15565 10047 15623 10053
rect 15565 10013 15577 10047
rect 15611 10013 15623 10047
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 15565 10007 15623 10013
rect 15764 10016 16221 10044
rect 10594 9976 10600 9988
rect 8260 9948 9812 9976
rect 10060 9948 10600 9976
rect 8260 9936 8266 9948
rect 8478 9908 8484 9920
rect 6932 9880 8484 9908
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 9674 9908 9680 9920
rect 8720 9880 9680 9908
rect 8720 9868 8726 9880
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9784 9908 9812 9948
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 9861 9911 9919 9917
rect 9861 9908 9873 9911
rect 9784 9880 9873 9908
rect 9861 9877 9873 9880
rect 9907 9877 9919 9911
rect 9861 9871 9919 9877
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 15764 9908 15792 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 17402 10044 17408 10056
rect 17363 10016 17408 10044
rect 16209 10007 16267 10013
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 17678 10004 17684 10056
rect 17736 10044 17742 10056
rect 18049 10047 18107 10053
rect 18049 10044 18061 10047
rect 17736 10016 18061 10044
rect 17736 10004 17742 10016
rect 18049 10013 18061 10016
rect 18095 10013 18107 10047
rect 18874 10044 18880 10056
rect 18835 10016 18880 10044
rect 18049 10007 18107 10013
rect 18874 10004 18880 10016
rect 18932 10004 18938 10056
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10044 19487 10047
rect 19518 10044 19524 10056
rect 19475 10016 19524 10044
rect 19475 10013 19487 10016
rect 19429 10007 19487 10013
rect 19518 10004 19524 10016
rect 19576 10004 19582 10056
rect 20257 10047 20315 10053
rect 20257 10013 20269 10047
rect 20303 10044 20315 10047
rect 20438 10044 20444 10056
rect 20303 10016 20444 10044
rect 20303 10013 20315 10016
rect 20257 10007 20315 10013
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 22066 9976 22094 10084
rect 23750 10004 23756 10056
rect 23808 10044 23814 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 23808 10016 24593 10044
rect 23808 10004 23814 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 25406 10044 25412 10056
rect 25367 10016 25412 10044
rect 24581 10007 24639 10013
rect 25406 10004 25412 10016
rect 25464 10004 25470 10056
rect 30098 10004 30104 10056
rect 30156 10044 30162 10056
rect 34885 10047 34943 10053
rect 34885 10044 34897 10047
rect 30156 10016 34897 10044
rect 30156 10004 30162 10016
rect 34885 10013 34897 10016
rect 34931 10013 34943 10047
rect 34885 10007 34943 10013
rect 22738 9976 22744 9988
rect 22066 9948 22744 9976
rect 22738 9936 22744 9948
rect 22796 9936 22802 9988
rect 24673 9979 24731 9985
rect 24673 9945 24685 9979
rect 24719 9976 24731 9979
rect 25590 9976 25596 9988
rect 24719 9948 25596 9976
rect 24719 9945 24731 9948
rect 24673 9939 24731 9945
rect 25590 9936 25596 9948
rect 25648 9936 25654 9988
rect 14608 9880 15792 9908
rect 35069 9911 35127 9917
rect 14608 9868 14614 9880
rect 35069 9877 35081 9911
rect 35115 9908 35127 9911
rect 38010 9908 38016 9920
rect 35115 9880 38016 9908
rect 35115 9877 35127 9880
rect 35069 9871 35127 9877
rect 38010 9868 38016 9880
rect 38068 9868 38074 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4706 9704 4712 9716
rect 4580 9676 4712 9704
rect 4580 9664 4586 9676
rect 4706 9664 4712 9676
rect 4764 9704 4770 9716
rect 8294 9704 8300 9716
rect 4764 9676 7972 9704
rect 8255 9676 8300 9704
rect 4764 9664 4770 9676
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 2832 9608 2877 9636
rect 2832 9596 2838 9608
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 4341 9639 4399 9645
rect 4341 9636 4353 9639
rect 3476 9608 4353 9636
rect 3476 9596 3482 9608
rect 4341 9605 4353 9608
rect 4387 9636 4399 9639
rect 6730 9636 6736 9648
rect 4387 9608 6736 9636
rect 4387 9605 4399 9608
rect 4341 9599 4399 9605
rect 6730 9596 6736 9608
rect 6788 9636 6794 9648
rect 7098 9636 7104 9648
rect 6788 9608 7104 9636
rect 6788 9596 6794 9608
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 7282 9636 7288 9648
rect 7243 9608 7288 9636
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 2038 9568 2044 9580
rect 1719 9540 2044 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5258 9568 5264 9580
rect 4847 9540 5264 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 5859 9540 6561 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 6549 9537 6561 9540
rect 6595 9568 6607 9571
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 6595 9540 7389 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 7377 9537 7389 9540
rect 7423 9568 7435 9571
rect 7466 9568 7472 9580
rect 7423 9540 7472 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 1762 9500 1768 9512
rect 1723 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2056 9500 2084 9528
rect 5828 9500 5856 9531
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 7944 9568 7972 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 11238 9704 11244 9716
rect 8444 9676 11244 9704
rect 8444 9664 8450 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 12526 9704 12532 9716
rect 12483 9676 12532 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 14829 9707 14887 9713
rect 14829 9673 14841 9707
rect 14875 9704 14887 9707
rect 14918 9704 14924 9716
rect 14875 9676 14924 9704
rect 14875 9673 14887 9676
rect 14829 9667 14887 9673
rect 14918 9664 14924 9676
rect 14976 9664 14982 9716
rect 16850 9704 16856 9716
rect 16811 9676 16856 9704
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 17402 9664 17408 9716
rect 17460 9704 17466 9716
rect 17681 9707 17739 9713
rect 17681 9704 17693 9707
rect 17460 9676 17693 9704
rect 17460 9664 17466 9676
rect 17681 9673 17693 9676
rect 17727 9673 17739 9707
rect 17681 9667 17739 9673
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 9585 9639 9643 9645
rect 9585 9636 9597 9639
rect 8168 9608 9597 9636
rect 8168 9596 8174 9608
rect 9585 9605 9597 9608
rect 9631 9605 9643 9639
rect 10594 9636 10600 9648
rect 10555 9608 10600 9636
rect 9585 9599 9643 9605
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 11146 9636 11152 9648
rect 11059 9608 11152 9636
rect 11146 9596 11152 9608
rect 11204 9636 11210 9648
rect 11974 9636 11980 9648
rect 11204 9608 11980 9636
rect 11204 9596 11210 9608
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 12066 9596 12072 9648
rect 12124 9636 12130 9648
rect 13633 9639 13691 9645
rect 12124 9608 13584 9636
rect 12124 9596 12130 9608
rect 9674 9568 9680 9580
rect 7944 9540 9680 9568
rect 9674 9528 9680 9540
rect 9732 9568 9738 9580
rect 10226 9568 10232 9580
rect 9732 9540 10232 9568
rect 9732 9528 9738 9540
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 12894 9568 12900 9580
rect 12855 9540 12900 9568
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 13556 9577 13584 9608
rect 13633 9605 13645 9639
rect 13679 9636 13691 9639
rect 13814 9636 13820 9648
rect 13679 9608 13820 9636
rect 13679 9605 13691 9608
rect 13633 9599 13691 9605
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 16209 9639 16267 9645
rect 13964 9608 15056 9636
rect 13964 9596 13970 9608
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9537 13599 9571
rect 14182 9568 14188 9580
rect 14143 9540 14188 9568
rect 13541 9531 13599 9537
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 14826 9568 14832 9580
rect 14323 9540 14832 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 15028 9577 15056 9608
rect 16209 9605 16221 9639
rect 16255 9636 16267 9639
rect 16482 9636 16488 9648
rect 16255 9608 16488 9636
rect 16255 9605 16267 9608
rect 16209 9599 16267 9605
rect 16482 9596 16488 9608
rect 16540 9596 16546 9648
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15654 9568 15660 9580
rect 15615 9540 15660 9568
rect 15013 9531 15071 9537
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 16301 9571 16359 9577
rect 16301 9568 16313 9571
rect 15988 9540 16313 9568
rect 15988 9528 15994 9540
rect 16301 9537 16313 9540
rect 16347 9568 16359 9571
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16347 9540 17049 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17736 9540 17877 9568
rect 17736 9528 17742 9540
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 34701 9571 34759 9577
rect 34701 9537 34713 9571
rect 34747 9568 34759 9571
rect 38102 9568 38108 9580
rect 34747 9540 38108 9568
rect 34747 9537 34759 9540
rect 34701 9531 34759 9537
rect 38102 9528 38108 9540
rect 38160 9528 38166 9580
rect 2056 9472 5856 9500
rect 5905 9503 5963 9509
rect 5905 9469 5917 9503
rect 5951 9500 5963 9503
rect 6178 9500 6184 9512
rect 5951 9472 6184 9500
rect 5951 9469 5963 9472
rect 5905 9463 5963 9469
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 8754 9500 8760 9512
rect 6687 9472 8760 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9500 10563 9503
rect 10686 9500 10692 9512
rect 10551 9472 10692 9500
rect 10551 9469 10563 9472
rect 10505 9463 10563 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 7558 9432 7564 9444
rect 2746 9404 7564 9432
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 2746 9364 2774 9404
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 13081 9435 13139 9441
rect 13081 9401 13093 9435
rect 13127 9432 13139 9435
rect 13354 9432 13360 9444
rect 13127 9404 13360 9432
rect 13127 9401 13139 9404
rect 13081 9395 13139 9401
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 15473 9435 15531 9441
rect 15473 9401 15485 9435
rect 15519 9432 15531 9435
rect 15562 9432 15568 9444
rect 15519 9404 15568 9432
rect 15519 9401 15531 9404
rect 15473 9395 15531 9401
rect 15562 9392 15568 9404
rect 15620 9392 15626 9444
rect 1728 9336 2774 9364
rect 4893 9367 4951 9373
rect 1728 9324 1734 9336
rect 4893 9333 4905 9367
rect 4939 9364 4951 9367
rect 7834 9364 7840 9376
rect 4939 9336 7840 9364
rect 4939 9333 4951 9336
rect 4893 9327 4951 9333
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 13538 9364 13544 9376
rect 8260 9336 13544 9364
rect 8260 9324 8266 9336
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 17586 9324 17592 9376
rect 17644 9364 17650 9376
rect 34609 9367 34667 9373
rect 34609 9364 34621 9367
rect 17644 9336 34621 9364
rect 17644 9324 17650 9336
rect 34609 9333 34621 9336
rect 34655 9333 34667 9367
rect 34609 9327 34667 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 3163 9163 3221 9169
rect 3163 9129 3175 9163
rect 3209 9160 3221 9163
rect 3970 9160 3976 9172
rect 3209 9132 3976 9160
rect 3209 9129 3221 9132
rect 3163 9123 3221 9129
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 5074 9160 5080 9172
rect 5035 9132 5080 9160
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 7926 9160 7932 9172
rect 5767 9132 7932 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 8478 9160 8484 9172
rect 8439 9132 8484 9160
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 9766 9160 9772 9172
rect 9727 9132 9772 9160
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 11333 9163 11391 9169
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 11606 9160 11612 9172
rect 11379 9132 11612 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 11848 9132 12081 9160
rect 11848 9120 11854 9132
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 12069 9123 12127 9129
rect 12710 9120 12716 9172
rect 12768 9160 12774 9172
rect 12805 9163 12863 9169
rect 12805 9160 12817 9163
rect 12768 9132 12817 9160
rect 12768 9120 12774 9132
rect 12805 9129 12817 9132
rect 12851 9129 12863 9163
rect 12805 9123 12863 9129
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 12952 9132 13553 9160
rect 12952 9120 12958 9132
rect 13541 9129 13553 9132
rect 13587 9129 13599 9163
rect 13541 9123 13599 9129
rect 14461 9163 14519 9169
rect 14461 9129 14473 9163
rect 14507 9160 14519 9163
rect 14642 9160 14648 9172
rect 14507 9132 14648 9160
rect 14507 9129 14519 9132
rect 14461 9123 14519 9129
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 15654 9160 15660 9172
rect 15615 9132 15660 9160
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 4065 9095 4123 9101
rect 4065 9061 4077 9095
rect 4111 9092 4123 9095
rect 5350 9092 5356 9104
rect 4111 9064 5356 9092
rect 4111 9061 4123 9064
rect 4065 9055 4123 9061
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 10134 9092 10140 9104
rect 7392 9064 10140 9092
rect 2130 8984 2136 9036
rect 2188 9024 2194 9036
rect 3421 9027 3479 9033
rect 3421 9024 3433 9027
rect 2188 8996 3433 9024
rect 2188 8984 2194 8996
rect 3421 8993 3433 8996
rect 3467 9024 3479 9027
rect 4614 9024 4620 9036
rect 3467 8996 4620 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 4614 8984 4620 8996
rect 4672 9024 4678 9036
rect 5074 9024 5080 9036
rect 4672 8996 5080 9024
rect 4672 8984 4678 8996
rect 5074 8984 5080 8996
rect 5132 9024 5138 9036
rect 5994 9024 6000 9036
rect 5132 8996 6000 9024
rect 5132 8984 5138 8996
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 7392 9024 7420 9064
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 6236 8996 7420 9024
rect 7469 9027 7527 9033
rect 6236 8984 6242 8996
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 8294 9024 8300 9036
rect 7515 8996 8300 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 14182 9024 14188 9036
rect 8536 8996 14188 9024
rect 8536 8984 8542 8996
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8956 4031 8959
rect 4154 8956 4160 8968
rect 4019 8928 4160 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 4154 8916 4160 8928
rect 4212 8956 4218 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 4212 8928 5181 8956
rect 4212 8916 4218 8928
rect 5169 8925 5181 8928
rect 5215 8956 5227 8959
rect 5442 8956 5448 8968
rect 5215 8928 5448 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 7484 8928 8401 8956
rect 1762 8848 1768 8900
rect 1820 8888 1826 8900
rect 1820 8860 1978 8888
rect 1820 8848 1826 8860
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 7193 8891 7251 8897
rect 5592 8860 6026 8888
rect 5592 8848 5598 8860
rect 7193 8857 7205 8891
rect 7239 8857 7251 8891
rect 7193 8851 7251 8857
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 5626 8820 5632 8832
rect 4120 8792 5632 8820
rect 4120 8780 4126 8792
rect 5626 8780 5632 8792
rect 5684 8780 5690 8832
rect 7208 8820 7236 8851
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 7484 8888 7512 8928
rect 8389 8925 8401 8928
rect 8435 8925 8447 8959
rect 9674 8956 9680 8968
rect 9635 8928 9680 8956
rect 8389 8919 8447 8925
rect 9674 8916 9680 8928
rect 9732 8956 9738 8968
rect 10962 8956 10968 8968
rect 9732 8928 10968 8956
rect 9732 8916 9738 8928
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11238 8956 11244 8968
rect 11199 8928 11244 8956
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11572 8928 11897 8956
rect 11572 8916 11578 8928
rect 11885 8925 11897 8928
rect 11931 8925 11943 8959
rect 12618 8956 12624 8968
rect 12579 8928 12624 8956
rect 11885 8919 11943 8925
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 13740 8965 13768 8996
rect 14182 8984 14188 8996
rect 14240 8984 14246 9036
rect 15010 9024 15016 9036
rect 14971 8996 15016 9024
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 14369 8959 14427 8965
rect 14369 8925 14381 8959
rect 14415 8956 14427 8959
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 14415 8928 15853 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 16482 8956 16488 8968
rect 16443 8928 16488 8956
rect 15841 8919 15899 8925
rect 7340 8860 7512 8888
rect 7340 8848 7346 8860
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 14384 8888 14412 8919
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 18601 8959 18659 8965
rect 18601 8956 18613 8959
rect 18288 8928 18613 8956
rect 18288 8916 18294 8928
rect 18601 8925 18613 8928
rect 18647 8925 18659 8959
rect 18601 8919 18659 8925
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 25133 8959 25191 8965
rect 25133 8956 25145 8959
rect 23072 8928 25145 8956
rect 23072 8916 23078 8928
rect 25133 8925 25145 8928
rect 25179 8925 25191 8959
rect 30834 8956 30840 8968
rect 30795 8928 30840 8956
rect 25133 8919 25191 8925
rect 30834 8916 30840 8928
rect 30892 8916 30898 8968
rect 38010 8956 38016 8968
rect 37971 8928 38016 8956
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 20346 8888 20352 8900
rect 7616 8860 14412 8888
rect 15396 8860 20352 8888
rect 7616 8848 7622 8860
rect 8846 8820 8852 8832
rect 7208 8792 8852 8820
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 10318 8820 10324 8832
rect 10279 8792 10324 8820
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 10410 8780 10416 8832
rect 10468 8820 10474 8832
rect 13354 8820 13360 8832
rect 10468 8792 13360 8820
rect 10468 8780 10474 8792
rect 13354 8780 13360 8792
rect 13412 8820 13418 8832
rect 15396 8820 15424 8860
rect 20346 8848 20352 8860
rect 20404 8848 20410 8900
rect 13412 8792 15424 8820
rect 13412 8780 13418 8792
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 15528 8792 16313 8820
rect 15528 8780 15534 8792
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 16301 8783 16359 8789
rect 18693 8823 18751 8829
rect 18693 8789 18705 8823
rect 18739 8820 18751 8823
rect 20162 8820 20168 8832
rect 18739 8792 20168 8820
rect 18739 8789 18751 8792
rect 18693 8783 18751 8789
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 25225 8823 25283 8829
rect 25225 8789 25237 8823
rect 25271 8820 25283 8823
rect 25498 8820 25504 8832
rect 25271 8792 25504 8820
rect 25271 8789 25283 8792
rect 25225 8783 25283 8789
rect 25498 8780 25504 8792
rect 25556 8780 25562 8832
rect 30929 8823 30987 8829
rect 30929 8789 30941 8823
rect 30975 8820 30987 8823
rect 33042 8820 33048 8832
rect 30975 8792 33048 8820
rect 30975 8789 30987 8792
rect 30929 8783 30987 8789
rect 33042 8780 33048 8792
rect 33100 8780 33106 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 5626 8576 5632 8628
rect 5684 8616 5690 8628
rect 6641 8619 6699 8625
rect 6641 8616 6653 8619
rect 5684 8588 6653 8616
rect 5684 8576 5690 8588
rect 6641 8585 6653 8588
rect 6687 8585 6699 8619
rect 6641 8579 6699 8585
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 7193 8619 7251 8625
rect 7193 8616 7205 8619
rect 6880 8588 7205 8616
rect 6880 8576 6886 8588
rect 7193 8585 7205 8588
rect 7239 8585 7251 8619
rect 7193 8579 7251 8585
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 7929 8619 7987 8625
rect 7340 8588 7788 8616
rect 7340 8576 7346 8588
rect 1946 8548 1952 8560
rect 1907 8520 1952 8548
rect 1946 8508 1952 8520
rect 2004 8508 2010 8560
rect 3694 8508 3700 8560
rect 3752 8548 3758 8560
rect 3752 8520 4554 8548
rect 3752 8508 3758 8520
rect 3050 8440 3056 8492
rect 3108 8440 3114 8492
rect 5994 8440 6000 8492
rect 6052 8480 6058 8492
rect 6052 8452 6097 8480
rect 6052 8440 6058 8452
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 6420 8452 6745 8480
rect 6420 8440 6426 8452
rect 6733 8449 6745 8452
rect 6779 8480 6791 8483
rect 7282 8480 7288 8492
rect 6779 8452 7288 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8480 7435 8483
rect 7466 8480 7472 8492
rect 7423 8452 7472 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7760 8480 7788 8588
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8018 8616 8024 8628
rect 7975 8588 8024 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8665 8619 8723 8625
rect 8665 8585 8677 8619
rect 8711 8616 8723 8619
rect 9214 8616 9220 8628
rect 8711 8588 9220 8616
rect 8711 8585 8723 8588
rect 8665 8579 8723 8585
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 10042 8616 10048 8628
rect 9447 8588 10048 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 10410 8616 10416 8628
rect 10371 8588 10416 8616
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11756 8588 11805 8616
rect 11756 8576 11762 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 12618 8616 12624 8628
rect 12579 8588 12624 8616
rect 11793 8579 11851 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 14737 8619 14795 8625
rect 14737 8585 14749 8619
rect 14783 8616 14795 8619
rect 15102 8616 15108 8628
rect 14783 8588 15108 8616
rect 14783 8585 14795 8588
rect 14737 8579 14795 8585
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15194 8576 15200 8628
rect 15252 8616 15258 8628
rect 15289 8619 15347 8625
rect 15289 8616 15301 8619
rect 15252 8588 15301 8616
rect 15252 8576 15258 8588
rect 15289 8585 15301 8588
rect 15335 8585 15347 8619
rect 15289 8579 15347 8585
rect 8110 8508 8116 8560
rect 8168 8548 8174 8560
rect 8168 8520 11836 8548
rect 8168 8508 8174 8520
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7760 8452 7849 8480
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 2038 8412 2044 8424
rect 1719 8384 2044 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 3326 8372 3332 8424
rect 3384 8412 3390 8424
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3384 8384 3433 8412
rect 3384 8372 3390 8384
rect 3421 8381 3433 8384
rect 3467 8412 3479 8415
rect 5626 8412 5632 8424
rect 3467 8384 5632 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 8202 8412 8208 8424
rect 5767 8384 8208 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 1578 8304 1584 8356
rect 1636 8304 1642 8356
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 8588 8344 8616 8443
rect 9232 8412 9260 8443
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 10321 8483 10379 8489
rect 10321 8480 10333 8483
rect 9916 8452 10333 8480
rect 9916 8440 9922 8452
rect 10321 8449 10333 8452
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 11020 8452 11161 8480
rect 11020 8440 11026 8452
rect 11149 8449 11161 8452
rect 11195 8449 11207 8483
rect 11698 8480 11704 8492
rect 11659 8452 11704 8480
rect 11149 8443 11207 8449
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11808 8480 11836 8520
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 16482 8548 16488 8560
rect 11940 8520 16488 8548
rect 11940 8508 11946 8520
rect 12805 8483 12863 8489
rect 12805 8480 12817 8483
rect 11808 8452 12817 8480
rect 12805 8449 12817 8452
rect 12851 8480 12863 8483
rect 14550 8480 14556 8492
rect 12851 8452 14556 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14660 8489 14688 8520
rect 16482 8508 16488 8520
rect 16540 8508 16546 8560
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 15470 8480 15476 8492
rect 15431 8452 15476 8480
rect 14645 8443 14703 8449
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 16022 8480 16028 8492
rect 15983 8452 16028 8480
rect 16022 8440 16028 8452
rect 16080 8440 16086 8492
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16356 8452 16865 8480
rect 16356 8440 16362 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 9232 8384 11008 8412
rect 10980 8353 11008 8384
rect 6972 8316 8616 8344
rect 10965 8347 11023 8353
rect 6972 8304 6978 8316
rect 10965 8313 10977 8347
rect 11011 8313 11023 8347
rect 10965 8307 11023 8313
rect 16117 8347 16175 8353
rect 16117 8313 16129 8347
rect 16163 8344 16175 8347
rect 16758 8344 16764 8356
rect 16163 8316 16764 8344
rect 16163 8313 16175 8316
rect 16117 8307 16175 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 16850 8304 16856 8356
rect 16908 8344 16914 8356
rect 16945 8347 17003 8353
rect 16945 8344 16957 8347
rect 16908 8316 16957 8344
rect 16908 8304 16914 8316
rect 16945 8313 16957 8316
rect 16991 8313 17003 8347
rect 16945 8307 17003 8313
rect 1596 8276 1624 8304
rect 1946 8276 1952 8288
rect 1596 8248 1952 8276
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 4249 8279 4307 8285
rect 4249 8245 4261 8279
rect 4295 8276 4307 8279
rect 4614 8276 4620 8288
rect 4295 8248 4620 8276
rect 4295 8245 4307 8248
rect 4249 8239 4307 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 11238 8276 11244 8288
rect 7432 8248 11244 8276
rect 7432 8236 7438 8248
rect 11238 8236 11244 8248
rect 11296 8276 11302 8288
rect 11606 8276 11612 8288
rect 11296 8248 11612 8276
rect 11296 8236 11302 8248
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2004 8044 4200 8072
rect 2004 8032 2010 8044
rect 3418 8004 3424 8016
rect 3379 7976 3424 8004
rect 3418 7964 3424 7976
rect 3476 7964 3482 8016
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 2038 7936 2044 7948
rect 1719 7908 2044 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 4172 7868 4200 8044
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 6825 8075 6883 8081
rect 4396 8044 6408 8072
rect 4396 8032 4402 8044
rect 4706 7964 4712 8016
rect 4764 8004 4770 8016
rect 6380 8004 6408 8044
rect 6825 8041 6837 8075
rect 6871 8072 6883 8075
rect 7374 8072 7380 8084
rect 6871 8044 7380 8072
rect 6871 8041 6883 8044
rect 6825 8035 6883 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 10594 8072 10600 8084
rect 9907 8044 10600 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 9766 8004 9772 8016
rect 4764 7976 5212 8004
rect 6380 7976 9772 8004
rect 4764 7964 4770 7976
rect 4246 7896 4252 7948
rect 4304 7936 4310 7948
rect 5074 7936 5080 7948
rect 4304 7908 5080 7936
rect 4304 7896 4310 7908
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5184 7936 5212 7976
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 5184 7908 5365 7936
rect 5353 7905 5365 7908
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6638 7936 6644 7948
rect 5868 7908 6644 7936
rect 5868 7896 5874 7908
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7936 7435 7939
rect 7423 7908 12434 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 4172 7840 4353 7868
rect 4341 7837 4353 7840
rect 4387 7868 4399 7871
rect 7282 7868 7288 7880
rect 4387 7840 4568 7868
rect 7243 7840 7288 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 1486 7760 1492 7812
rect 1544 7800 1550 7812
rect 1949 7803 2007 7809
rect 1949 7800 1961 7803
rect 1544 7772 1961 7800
rect 1544 7760 1550 7772
rect 1949 7769 1961 7772
rect 1995 7769 2007 7803
rect 1949 7763 2007 7769
rect 2958 7760 2964 7812
rect 3016 7760 3022 7812
rect 4430 7800 4436 7812
rect 4391 7772 4436 7800
rect 4430 7760 4436 7772
rect 4488 7760 4494 7812
rect 4540 7800 4568 7840
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 11606 7868 11612 7880
rect 9723 7840 11468 7868
rect 11567 7840 11612 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 5258 7800 5264 7812
rect 4540 7772 5264 7800
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 5810 7760 5816 7812
rect 5868 7760 5874 7812
rect 8588 7800 8616 7831
rect 11146 7800 11152 7812
rect 8588 7772 11152 7800
rect 11146 7760 11152 7772
rect 11204 7760 11210 7812
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 4982 7732 4988 7744
rect 4764 7704 4988 7732
rect 4764 7692 4770 7704
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 8478 7732 8484 7744
rect 8439 7704 8484 7732
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 11440 7741 11468 7840
rect 11606 7828 11612 7840
rect 11664 7828 11670 7880
rect 12406 7800 12434 7908
rect 33042 7828 33048 7880
rect 33100 7868 33106 7880
rect 35345 7871 35403 7877
rect 35345 7868 35357 7871
rect 33100 7840 35357 7868
rect 33100 7828 33106 7840
rect 35345 7837 35357 7840
rect 35391 7837 35403 7871
rect 35345 7831 35403 7837
rect 14734 7800 14740 7812
rect 12406 7772 14740 7800
rect 14734 7760 14740 7772
rect 14792 7760 14798 7812
rect 11425 7735 11483 7741
rect 11425 7701 11437 7735
rect 11471 7701 11483 7735
rect 11425 7695 11483 7701
rect 35529 7735 35587 7741
rect 35529 7701 35541 7735
rect 35575 7732 35587 7735
rect 38010 7732 38016 7744
rect 35575 7704 38016 7732
rect 35575 7701 35587 7704
rect 35529 7695 35587 7701
rect 38010 7692 38016 7704
rect 38068 7692 38074 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 1673 7531 1731 7537
rect 1673 7528 1685 7531
rect 1636 7500 1685 7528
rect 1636 7488 1642 7500
rect 1673 7497 1685 7500
rect 1719 7497 1731 7531
rect 1673 7491 1731 7497
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3142 7528 3148 7540
rect 3099 7500 3148 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 3697 7531 3755 7537
rect 3697 7497 3709 7531
rect 3743 7528 3755 7531
rect 5166 7528 5172 7540
rect 3743 7500 5172 7528
rect 3743 7497 3755 7500
rect 3697 7491 3755 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 6638 7528 6644 7540
rect 5500 7500 5856 7528
rect 6599 7500 6644 7528
rect 5500 7488 5506 7500
rect 4154 7460 4160 7472
rect 3620 7432 4160 7460
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 1872 7188 1900 7355
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 3620 7401 3648 7432
rect 4154 7420 4160 7432
rect 4212 7420 4218 7472
rect 4982 7420 4988 7472
rect 5040 7420 5046 7472
rect 2317 7395 2375 7401
rect 2317 7392 2329 7395
rect 2004 7364 2329 7392
rect 2004 7352 2010 7364
rect 2317 7361 2329 7364
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 4246 7392 4252 7404
rect 4207 7364 4252 7392
rect 3605 7355 3663 7361
rect 2409 7327 2467 7333
rect 2409 7293 2421 7327
rect 2455 7324 2467 7327
rect 3160 7324 3188 7355
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 5828 7392 5856 7500
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 9214 7528 9220 7540
rect 9175 7500 9220 7528
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 24394 7488 24400 7540
rect 24452 7528 24458 7540
rect 24581 7531 24639 7537
rect 24581 7528 24593 7531
rect 24452 7500 24593 7528
rect 24452 7488 24458 7500
rect 24581 7497 24593 7500
rect 24627 7497 24639 7531
rect 38102 7528 38108 7540
rect 38063 7500 38108 7528
rect 24581 7491 24639 7497
rect 38102 7488 38108 7500
rect 38160 7488 38166 7540
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5828 7364 6561 7392
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 9125 7395 9183 7401
rect 9125 7392 9137 7395
rect 6696 7364 9137 7392
rect 6696 7352 6702 7364
rect 9125 7361 9137 7364
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 24673 7395 24731 7401
rect 24673 7361 24685 7395
rect 24719 7392 24731 7395
rect 29730 7392 29736 7404
rect 24719 7364 29736 7392
rect 24719 7361 24731 7364
rect 24673 7355 24731 7361
rect 29730 7352 29736 7364
rect 29788 7352 29794 7404
rect 34330 7352 34336 7404
rect 34388 7392 34394 7404
rect 34425 7395 34483 7401
rect 34425 7392 34437 7395
rect 34388 7364 34437 7392
rect 34388 7352 34394 7364
rect 34425 7361 34437 7364
rect 34471 7361 34483 7395
rect 38286 7392 38292 7404
rect 38247 7364 38292 7392
rect 34425 7355 34483 7361
rect 38286 7352 38292 7364
rect 38344 7352 38350 7404
rect 3786 7324 3792 7336
rect 2455 7296 2774 7324
rect 3160 7296 3792 7324
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 2746 7256 2774 7296
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7324 4583 7327
rect 4614 7324 4620 7336
rect 4571 7296 4620 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 4614 7284 4620 7296
rect 4672 7324 4678 7336
rect 5074 7324 5080 7336
rect 4672 7296 5080 7324
rect 4672 7284 4678 7296
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 4246 7256 4252 7268
rect 2746 7228 4252 7256
rect 4246 7216 4252 7228
rect 4304 7216 4310 7268
rect 5997 7259 6055 7265
rect 5997 7225 6009 7259
rect 6043 7256 6055 7259
rect 12066 7256 12072 7268
rect 6043 7228 12072 7256
rect 6043 7225 6055 7228
rect 5997 7219 6055 7225
rect 12066 7216 12072 7228
rect 12124 7216 12130 7268
rect 22646 7216 22652 7268
rect 22704 7256 22710 7268
rect 34333 7259 34391 7265
rect 34333 7256 34345 7259
rect 22704 7228 34345 7256
rect 22704 7216 22710 7228
rect 34333 7225 34345 7228
rect 34379 7225 34391 7259
rect 34333 7219 34391 7225
rect 4614 7188 4620 7200
rect 1872 7160 4620 7188
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 5905 6987 5963 6993
rect 5905 6984 5917 6987
rect 2280 6956 5917 6984
rect 2280 6944 2286 6956
rect 5905 6953 5917 6956
rect 5951 6953 5963 6987
rect 5905 6947 5963 6953
rect 4617 6919 4675 6925
rect 3068 6888 3832 6916
rect 2682 6848 2688 6860
rect 2643 6820 2688 6848
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 2866 6780 2872 6792
rect 2639 6752 2872 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 2866 6740 2872 6752
rect 2924 6780 2930 6792
rect 3068 6780 3096 6888
rect 3694 6848 3700 6860
rect 2924 6752 3096 6780
rect 3160 6820 3700 6848
rect 2924 6740 2930 6752
rect 2041 6715 2099 6721
rect 2041 6681 2053 6715
rect 2087 6712 2099 6715
rect 3160 6712 3188 6820
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 3804 6848 3832 6888
rect 4617 6885 4629 6919
rect 4663 6916 4675 6919
rect 4663 6888 5856 6916
rect 4663 6885 4675 6888
rect 4617 6879 4675 6885
rect 5261 6851 5319 6857
rect 3804 6820 4660 6848
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 2087 6684 3188 6712
rect 2087 6681 2099 6684
rect 2041 6675 2099 6681
rect 3252 6644 3280 6743
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 4533 6785 4591 6791
rect 3384 6752 3429 6780
rect 3384 6740 3390 6752
rect 4533 6751 4545 6785
rect 4579 6782 4591 6785
rect 4632 6782 4660 6820
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5718 6848 5724 6860
rect 5307 6820 5724 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 5828 6848 5856 6888
rect 5994 6876 6000 6928
rect 6052 6916 6058 6928
rect 7190 6916 7196 6928
rect 6052 6888 7196 6916
rect 6052 6876 6058 6888
rect 7190 6876 7196 6888
rect 7248 6876 7254 6928
rect 9508 6888 9812 6916
rect 9508 6848 9536 6888
rect 5828 6820 9536 6848
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9640 6820 9689 6848
rect 9640 6808 9646 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9784 6848 9812 6888
rect 10778 6848 10784 6860
rect 9784 6820 10784 6848
rect 9677 6811 9735 6817
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 14369 6851 14427 6857
rect 14369 6817 14381 6851
rect 14415 6848 14427 6851
rect 14458 6848 14464 6860
rect 14415 6820 14464 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 21269 6851 21327 6857
rect 21269 6817 21281 6851
rect 21315 6848 21327 6851
rect 21542 6848 21548 6860
rect 21315 6820 21548 6848
rect 21315 6817 21327 6820
rect 21269 6811 21327 6817
rect 21542 6808 21548 6820
rect 21600 6808 21606 6860
rect 35161 6851 35219 6857
rect 35161 6848 35173 6851
rect 23492 6820 35173 6848
rect 4579 6780 4660 6782
rect 4706 6780 4712 6792
rect 4579 6754 4712 6780
rect 4579 6751 4591 6754
rect 4632 6752 4712 6754
rect 4533 6745 4591 6751
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 3786 6672 3792 6724
rect 3844 6712 3850 6724
rect 5184 6712 5212 6743
rect 5442 6740 5448 6792
rect 5500 6780 5506 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5500 6752 6009 6780
rect 5500 6740 5506 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6749 6515 6783
rect 14274 6780 14280 6792
rect 14235 6752 14280 6780
rect 6457 6743 6515 6749
rect 3844 6684 5212 6712
rect 3844 6672 3850 6684
rect 3326 6644 3332 6656
rect 3252 6616 3332 6644
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 6472 6644 6500 6743
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6780 21419 6783
rect 23382 6780 23388 6792
rect 21407 6752 23388 6780
rect 21407 6749 21419 6752
rect 21361 6743 21419 6749
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 9217 6715 9275 6721
rect 9217 6712 9229 6715
rect 8812 6684 9229 6712
rect 8812 6672 8818 6684
rect 9217 6681 9229 6684
rect 9263 6681 9275 6715
rect 9217 6675 9275 6681
rect 9306 6672 9312 6724
rect 9364 6712 9370 6724
rect 9364 6684 9409 6712
rect 9364 6672 9370 6684
rect 20806 6672 20812 6724
rect 20864 6712 20870 6724
rect 23492 6712 23520 6820
rect 35161 6817 35173 6820
rect 35207 6817 35219 6851
rect 35161 6811 35219 6817
rect 29917 6783 29975 6789
rect 29917 6749 29929 6783
rect 29963 6780 29975 6783
rect 30558 6780 30564 6792
rect 29963 6752 30564 6780
rect 29963 6749 29975 6752
rect 29917 6743 29975 6749
rect 30558 6740 30564 6752
rect 30616 6740 30622 6792
rect 30745 6783 30803 6789
rect 30745 6749 30757 6783
rect 30791 6780 30803 6783
rect 33042 6780 33048 6792
rect 30791 6752 33048 6780
rect 30791 6749 30803 6752
rect 30745 6743 30803 6749
rect 33042 6740 33048 6752
rect 33100 6740 33106 6792
rect 35253 6783 35311 6789
rect 35253 6749 35265 6783
rect 35299 6780 35311 6783
rect 35618 6780 35624 6792
rect 35299 6752 35624 6780
rect 35299 6749 35311 6752
rect 35253 6743 35311 6749
rect 35618 6740 35624 6752
rect 35676 6740 35682 6792
rect 30653 6715 30711 6721
rect 30653 6712 30665 6715
rect 20864 6684 23520 6712
rect 23584 6684 30665 6712
rect 20864 6672 20870 6684
rect 4764 6616 6500 6644
rect 6549 6647 6607 6653
rect 4764 6604 4770 6616
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 12802 6644 12808 6656
rect 6595 6616 12808 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 20070 6604 20076 6656
rect 20128 6644 20134 6656
rect 23584 6644 23612 6684
rect 30653 6681 30665 6684
rect 30699 6681 30711 6715
rect 30653 6675 30711 6681
rect 20128 6616 23612 6644
rect 20128 6604 20134 6616
rect 24486 6604 24492 6656
rect 24544 6644 24550 6656
rect 29825 6647 29883 6653
rect 29825 6644 29837 6647
rect 24544 6616 29837 6644
rect 24544 6604 24550 6616
rect 29825 6613 29837 6616
rect 29871 6613 29883 6647
rect 29825 6607 29883 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 2590 6440 2596 6452
rect 1596 6412 2596 6440
rect 1596 6313 1624 6412
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 2685 6443 2743 6449
rect 2685 6409 2697 6443
rect 2731 6440 2743 6443
rect 2958 6440 2964 6452
rect 2731 6412 2964 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3329 6443 3387 6449
rect 3329 6409 3341 6443
rect 3375 6440 3387 6443
rect 3510 6440 3516 6452
rect 3375 6412 3516 6440
rect 3375 6409 3387 6412
rect 3329 6403 3387 6409
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 3878 6400 3884 6452
rect 3936 6440 3942 6452
rect 4065 6443 4123 6449
rect 4065 6440 4077 6443
rect 3936 6412 4077 6440
rect 3936 6400 3942 6412
rect 4065 6409 4077 6412
rect 4111 6409 4123 6443
rect 4065 6403 4123 6409
rect 4709 6443 4767 6449
rect 4709 6409 4721 6443
rect 4755 6440 4767 6443
rect 4798 6440 4804 6452
rect 4755 6412 4804 6440
rect 4755 6409 4767 6412
rect 4709 6403 4767 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 5353 6443 5411 6449
rect 5353 6409 5365 6443
rect 5399 6440 5411 6443
rect 8754 6440 8760 6452
rect 5399 6412 8760 6440
rect 5399 6409 5411 6412
rect 5353 6403 5411 6409
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 8849 6443 8907 6449
rect 8849 6409 8861 6443
rect 8895 6440 8907 6443
rect 9306 6440 9312 6452
rect 8895 6412 9312 6440
rect 8895 6409 8907 6412
rect 8849 6403 8907 6409
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 6362 6372 6368 6384
rect 2608 6344 4200 6372
rect 2608 6313 2636 6344
rect 4172 6316 4200 6344
rect 4632 6344 6368 6372
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 2958 6264 2964 6316
rect 3016 6304 3022 6316
rect 3326 6304 3332 6316
rect 3016 6276 3332 6304
rect 3016 6264 3022 6276
rect 3326 6264 3332 6276
rect 3384 6304 3390 6316
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 3384 6276 3433 6304
rect 3384 6264 3390 6276
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 4154 6304 4160 6316
rect 4115 6276 4160 6304
rect 3421 6267 3479 6273
rect 3436 6236 3464 6267
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 4632 6313 4660 6344
rect 6362 6332 6368 6344
rect 6420 6332 6426 6384
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 5258 6304 5264 6316
rect 5219 6276 5264 6304
rect 4617 6267 4675 6273
rect 4632 6236 4660 6267
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 6730 6304 6736 6316
rect 6691 6276 6736 6304
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 8021 6307 8079 6313
rect 8021 6273 8033 6307
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 3436 6208 4660 6236
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 8036 6236 8064 6267
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8628 6276 8677 6304
rect 8628 6264 8634 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8772 6304 8800 6400
rect 13446 6304 13452 6316
rect 8772 6276 13452 6304
rect 8665 6267 8723 6273
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 28169 6307 28227 6313
rect 28169 6273 28181 6307
rect 28215 6304 28227 6307
rect 30282 6304 30288 6316
rect 28215 6276 30288 6304
rect 28215 6273 28227 6276
rect 28169 6267 28227 6273
rect 30282 6264 30288 6276
rect 30340 6264 30346 6316
rect 4856 6208 8064 6236
rect 8113 6239 8171 6245
rect 4856 6196 4862 6208
rect 8113 6205 8125 6239
rect 8159 6236 8171 6239
rect 11054 6236 11060 6248
rect 8159 6208 11060 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 11698 6168 11704 6180
rect 1811 6140 11704 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 11698 6128 11704 6140
rect 11756 6128 11762 6180
rect 6362 6060 6368 6112
rect 6420 6100 6426 6112
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 6420 6072 6653 6100
rect 6420 6060 6426 6072
rect 6641 6069 6653 6072
rect 6687 6069 6699 6103
rect 6641 6063 6699 6069
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 28077 6103 28135 6109
rect 28077 6100 28089 6103
rect 16724 6072 28089 6100
rect 16724 6060 16730 6072
rect 28077 6069 28089 6072
rect 28123 6069 28135 6103
rect 28077 6063 28135 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5896 2743 5899
rect 3050 5896 3056 5908
rect 2731 5868 3056 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 4890 5896 4896 5908
rect 4479 5868 4896 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 5074 5856 5080 5908
rect 5132 5896 5138 5908
rect 6730 5896 6736 5908
rect 5132 5868 6736 5896
rect 5132 5856 5138 5868
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9950 5896 9956 5908
rect 9911 5868 9956 5896
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 15565 5899 15623 5905
rect 15565 5865 15577 5899
rect 15611 5896 15623 5899
rect 15746 5896 15752 5908
rect 15611 5868 15752 5896
rect 15611 5865 15623 5868
rect 15565 5859 15623 5865
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 3234 5828 3240 5840
rect 2746 5800 3240 5828
rect 2746 5760 2774 5800
rect 3234 5788 3240 5800
rect 3292 5788 3298 5840
rect 3329 5831 3387 5837
rect 3329 5797 3341 5831
rect 3375 5828 3387 5831
rect 6825 5831 6883 5837
rect 3375 5800 6316 5828
rect 3375 5797 3387 5800
rect 3329 5791 3387 5797
rect 6288 5769 6316 5800
rect 6825 5797 6837 5831
rect 6871 5828 6883 5831
rect 9582 5828 9588 5840
rect 6871 5800 9588 5828
rect 6871 5797 6883 5800
rect 6825 5791 6883 5797
rect 9582 5788 9588 5800
rect 9640 5788 9646 5840
rect 1596 5732 2774 5760
rect 6273 5763 6331 5769
rect 1596 5701 1624 5732
rect 6273 5729 6285 5763
rect 6319 5729 6331 5763
rect 6273 5723 6331 5729
rect 6730 5720 6736 5772
rect 6788 5760 6794 5772
rect 6788 5732 8432 5760
rect 6788 5720 6794 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2958 5692 2964 5704
rect 2639 5664 2964 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3234 5692 3240 5704
rect 3195 5664 3240 5692
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 4120 5664 4353 5692
rect 4120 5652 4126 5664
rect 4341 5661 4353 5664
rect 4387 5661 4399 5695
rect 4341 5655 4399 5661
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5692 5779 5695
rect 5902 5692 5908 5704
rect 5767 5664 5908 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 7926 5692 7932 5704
rect 7887 5664 7932 5692
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8404 5701 8432 5732
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 8389 5655 8447 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 15470 5692 15476 5704
rect 15431 5664 15476 5692
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 32858 5692 32864 5704
rect 32819 5664 32864 5692
rect 32858 5652 32864 5664
rect 32916 5652 32922 5704
rect 36814 5692 36820 5704
rect 36775 5664 36820 5692
rect 36814 5652 36820 5664
rect 36872 5652 36878 5704
rect 38010 5692 38016 5704
rect 37971 5664 38016 5692
rect 38010 5652 38016 5664
rect 38068 5652 38074 5704
rect 5994 5624 6000 5636
rect 2746 5596 6000 5624
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5556 1823 5559
rect 2746 5556 2774 5596
rect 5994 5584 6000 5596
rect 6052 5584 6058 5636
rect 6362 5584 6368 5636
rect 6420 5624 6426 5636
rect 6420 5596 6465 5624
rect 6420 5584 6426 5596
rect 7558 5584 7564 5636
rect 7616 5624 7622 5636
rect 7653 5627 7711 5633
rect 7653 5624 7665 5627
rect 7616 5596 7665 5624
rect 7616 5584 7622 5596
rect 7653 5593 7665 5596
rect 7699 5593 7711 5627
rect 7653 5587 7711 5593
rect 5626 5556 5632 5568
rect 1811 5528 2774 5556
rect 5587 5528 5632 5556
rect 1811 5525 1823 5528
rect 1765 5519 1823 5525
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 33045 5559 33103 5565
rect 33045 5525 33057 5559
rect 33091 5556 33103 5559
rect 34422 5556 34428 5568
rect 33091 5528 34428 5556
rect 33091 5525 33103 5528
rect 33045 5519 33103 5525
rect 34422 5516 34428 5528
rect 34480 5516 34486 5568
rect 36909 5559 36967 5565
rect 36909 5525 36921 5559
rect 36955 5556 36967 5559
rect 37458 5556 37464 5568
rect 36955 5528 37464 5556
rect 36955 5525 36967 5528
rect 36909 5519 36967 5525
rect 37458 5516 37464 5528
rect 37516 5516 37522 5568
rect 38194 5556 38200 5568
rect 38155 5528 38200 5556
rect 38194 5516 38200 5528
rect 38252 5516 38258 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4614 5352 4620 5364
rect 4295 5324 4620 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 4982 5352 4988 5364
rect 4943 5324 4988 5352
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 8478 5284 8484 5296
rect 4448 5256 8484 5284
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 2866 5216 2872 5228
rect 2731 5188 2872 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 1670 5012 1676 5024
rect 1631 4984 1676 5012
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 1872 5012 1900 5179
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 4338 5216 4344 5228
rect 3375 5188 4344 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 4448 5225 4476 5256
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4890 5216 4896 5228
rect 4803 5188 4896 5216
rect 4433 5179 4491 5185
rect 4890 5176 4896 5188
rect 4948 5216 4954 5228
rect 5350 5216 5356 5228
rect 4948 5188 5356 5216
rect 4948 5176 4954 5188
rect 5350 5176 5356 5188
rect 5408 5216 5414 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 5408 5188 7665 5216
rect 5408 5176 5414 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 7926 5216 7932 5228
rect 7887 5188 7932 5216
rect 7653 5179 7711 5185
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 16850 5216 16856 5228
rect 16811 5188 16856 5216
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 20162 5216 20168 5228
rect 20123 5188 20168 5216
rect 20162 5176 20168 5188
rect 20220 5176 20226 5228
rect 25498 5216 25504 5228
rect 25459 5188 25504 5216
rect 25498 5176 25504 5188
rect 25556 5176 25562 5228
rect 25590 5176 25596 5228
rect 25648 5216 25654 5228
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 25648 5188 27169 5216
rect 25648 5176 25654 5188
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 37458 5216 37464 5228
rect 37419 5188 37464 5216
rect 27157 5179 27215 5185
rect 37458 5176 37464 5188
rect 37516 5176 37522 5228
rect 2777 5151 2835 5157
rect 2777 5117 2789 5151
rect 2823 5148 2835 5151
rect 7006 5148 7012 5160
rect 2823 5120 7012 5148
rect 2823 5117 2835 5120
rect 2777 5111 2835 5117
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 6822 5080 6828 5092
rect 2746 5052 6828 5080
rect 2746 5012 2774 5052
rect 6822 5040 6828 5052
rect 6880 5040 6886 5092
rect 25685 5083 25743 5089
rect 25685 5049 25697 5083
rect 25731 5080 25743 5083
rect 27798 5080 27804 5092
rect 25731 5052 27804 5080
rect 25731 5049 25743 5052
rect 25685 5043 25743 5049
rect 27798 5040 27804 5052
rect 27856 5040 27862 5092
rect 3418 5012 3424 5024
rect 1872 4984 2774 5012
rect 3379 4984 3424 5012
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 4338 4972 4344 5024
rect 4396 5012 4402 5024
rect 7558 5012 7564 5024
rect 4396 4984 7564 5012
rect 4396 4972 4402 4984
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 17037 5015 17095 5021
rect 17037 4981 17049 5015
rect 17083 5012 17095 5015
rect 20070 5012 20076 5024
rect 17083 4984 20076 5012
rect 17083 4981 17095 4984
rect 17037 4975 17095 4981
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 20349 5015 20407 5021
rect 20349 4981 20361 5015
rect 20395 5012 20407 5015
rect 23290 5012 23296 5024
rect 20395 4984 23296 5012
rect 20395 4981 20407 4984
rect 20349 4975 20407 4981
rect 23290 4972 23296 4984
rect 23348 4972 23354 5024
rect 27341 5015 27399 5021
rect 27341 4981 27353 5015
rect 27387 5012 27399 5015
rect 30006 5012 30012 5024
rect 27387 4984 30012 5012
rect 27387 4981 27399 4984
rect 27341 4975 27399 4981
rect 30006 4972 30012 4984
rect 30064 4972 30070 5024
rect 37645 5015 37703 5021
rect 37645 4981 37657 5015
rect 37691 5012 37703 5015
rect 38010 5012 38016 5024
rect 37691 4984 38016 5012
rect 37691 4981 37703 4984
rect 37645 4975 37703 4981
rect 38010 4972 38016 4984
rect 38068 4972 38074 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 1762 4808 1768 4820
rect 1719 4780 1768 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 2961 4811 3019 4817
rect 2961 4777 2973 4811
rect 3007 4808 3019 4811
rect 3602 4808 3608 4820
rect 3007 4780 3608 4808
rect 3007 4777 3019 4780
rect 2961 4771 3019 4777
rect 3602 4768 3608 4780
rect 3660 4768 3666 4820
rect 4065 4811 4123 4817
rect 4065 4777 4077 4811
rect 4111 4808 4123 4811
rect 6454 4808 6460 4820
rect 4111 4780 6460 4808
rect 4111 4777 4123 4780
rect 4065 4771 4123 4777
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 2317 4743 2375 4749
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 5810 4740 5816 4752
rect 2363 4712 5816 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 5810 4700 5816 4712
rect 5868 4700 5874 4752
rect 3418 4632 3424 4684
rect 3476 4672 3482 4684
rect 6546 4672 6552 4684
rect 3476 4644 6552 4672
rect 3476 4632 3482 4644
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 7650 4632 7656 4684
rect 7708 4672 7714 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 7708 4644 9321 4672
rect 7708 4632 7714 4644
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1728 4576 1777 4604
rect 1728 4564 1734 4576
rect 1765 4573 1777 4576
rect 1811 4604 1823 4607
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 1811 4576 2237 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 2225 4573 2237 4576
rect 2271 4604 2283 4607
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2271 4576 2881 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 2869 4573 2881 4576
rect 2915 4604 2927 4607
rect 3786 4604 3792 4616
rect 2915 4576 3792 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 5626 4604 5632 4616
rect 4847 4576 5632 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 2958 4496 2964 4548
rect 3016 4536 3022 4548
rect 3988 4536 4016 4567
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 7926 4604 7932 4616
rect 7839 4576 7932 4604
rect 7926 4564 7932 4576
rect 7984 4604 7990 4616
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 7984 4576 9597 4604
rect 7984 4564 7990 4576
rect 9585 4573 9597 4576
rect 9631 4604 9643 4607
rect 12618 4604 12624 4616
rect 9631 4576 12624 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 16758 4564 16764 4616
rect 16816 4604 16822 4616
rect 16945 4607 17003 4613
rect 16945 4604 16957 4607
rect 16816 4576 16957 4604
rect 16816 4564 16822 4576
rect 16945 4573 16957 4576
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 7653 4539 7711 4545
rect 7653 4536 7665 4539
rect 3016 4508 7665 4536
rect 3016 4496 3022 4508
rect 7653 4505 7665 4508
rect 7699 4505 7711 4539
rect 7653 4499 7711 4505
rect 4614 4468 4620 4480
rect 4575 4440 4620 4468
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 17129 4471 17187 4477
rect 17129 4437 17141 4471
rect 17175 4468 17187 4471
rect 18598 4468 18604 4480
rect 17175 4440 18604 4468
rect 17175 4437 17187 4440
rect 17129 4431 17187 4437
rect 18598 4428 18604 4440
rect 18656 4428 18662 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1670 4128 1676 4140
rect 1631 4100 1676 4128
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 2222 4088 2228 4140
rect 2280 4128 2286 4140
rect 2777 4131 2835 4137
rect 2777 4128 2789 4131
rect 2280 4100 2789 4128
rect 2280 4088 2286 4100
rect 2777 4097 2789 4100
rect 2823 4128 2835 4131
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 2823 4100 3433 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 3421 4097 3433 4100
rect 3467 4128 3479 4131
rect 4890 4128 4896 4140
rect 3467 4100 4896 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4128 9827 4131
rect 17310 4128 17316 4140
rect 9815 4100 17316 4128
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 1394 4020 1400 4072
rect 1452 4060 1458 4072
rect 1765 4063 1823 4069
rect 1765 4060 1777 4063
rect 1452 4032 1777 4060
rect 1452 4020 1458 4032
rect 1765 4029 1777 4032
rect 1811 4029 1823 4063
rect 1765 4023 1823 4029
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 9214 4060 9220 4072
rect 2915 4032 9220 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 3510 3992 3516 4004
rect 3471 3964 3516 3992
rect 3510 3952 3516 3964
rect 3568 3952 3574 4004
rect 9582 3884 9588 3936
rect 9640 3924 9646 3936
rect 9677 3927 9735 3933
rect 9677 3924 9689 3927
rect 9640 3896 9689 3924
rect 9640 3884 9646 3896
rect 9677 3893 9689 3896
rect 9723 3893 9735 3927
rect 9677 3887 9735 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2225 3723 2283 3729
rect 2225 3689 2237 3723
rect 2271 3720 2283 3723
rect 2406 3720 2412 3732
rect 2271 3692 2412 3720
rect 2271 3689 2283 3692
rect 2225 3683 2283 3689
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 4157 3723 4215 3729
rect 4157 3689 4169 3723
rect 4203 3720 4215 3723
rect 4706 3720 4712 3732
rect 4203 3692 4712 3720
rect 4203 3689 4215 3692
rect 4157 3683 4215 3689
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 30742 3680 30748 3732
rect 30800 3720 30806 3732
rect 38105 3723 38163 3729
rect 38105 3720 38117 3723
rect 30800 3692 38117 3720
rect 30800 3680 30806 3692
rect 38105 3689 38117 3692
rect 38151 3689 38163 3723
rect 38105 3683 38163 3689
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 7742 3652 7748 3664
rect 2915 3624 7748 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 7742 3612 7748 3624
rect 7800 3612 7806 3664
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3516 2375 3519
rect 2777 3519 2835 3525
rect 2777 3516 2789 3519
rect 2363 3488 2789 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 2777 3485 2789 3488
rect 2823 3516 2835 3519
rect 2958 3516 2964 3528
rect 2823 3488 2964 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 38286 3516 38292 3528
rect 38247 3488 38292 3516
rect 38286 3476 38292 3488
rect 38344 3476 38350 3528
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3176 2375 3179
rect 3053 3179 3111 3185
rect 2363 3148 3004 3176
rect 2363 3145 2375 3148
rect 2317 3139 2375 3145
rect 2774 3108 2780 3120
rect 2148 3080 2780 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 2148 3040 2176 3080
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 2976 3108 3004 3148
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 5258 3176 5264 3188
rect 3099 3148 5264 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 35618 3136 35624 3188
rect 35676 3176 35682 3188
rect 36725 3179 36783 3185
rect 36725 3176 36737 3179
rect 35676 3148 36737 3176
rect 35676 3136 35682 3148
rect 36725 3145 36737 3148
rect 36771 3145 36783 3179
rect 36725 3139 36783 3145
rect 5534 3108 5540 3120
rect 2976 3080 5540 3108
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 1627 3012 2176 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2222 3000 2228 3052
rect 2280 3040 2286 3052
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2280 3012 2325 3040
rect 2746 3012 2881 3040
rect 2280 3000 2286 3012
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 2746 2972 2774 3012
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 3510 3040 3516 3052
rect 3471 3012 3516 3040
rect 2869 3003 2927 3009
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 9582 3040 9588 3052
rect 9543 3012 9588 3040
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 36909 3043 36967 3049
rect 36909 3009 36921 3043
rect 36955 3040 36967 3043
rect 37274 3040 37280 3052
rect 36955 3012 37280 3040
rect 36955 3009 36967 3012
rect 36909 3003 36967 3009
rect 37274 3000 37280 3012
rect 37332 3000 37338 3052
rect 38010 3040 38016 3052
rect 37971 3012 38016 3040
rect 38010 3000 38016 3012
rect 38068 3000 38074 3052
rect 1360 2944 2774 2972
rect 1360 2932 1366 2944
rect 3697 2907 3755 2913
rect 3697 2873 3709 2907
rect 3743 2904 3755 2907
rect 6914 2904 6920 2916
rect 3743 2876 6920 2904
rect 3743 2873 3755 2876
rect 3697 2867 3755 2873
rect 6914 2864 6920 2876
rect 6972 2864 6978 2916
rect 1765 2839 1823 2845
rect 1765 2805 1777 2839
rect 1811 2836 1823 2839
rect 6638 2836 6644 2848
rect 1811 2808 6644 2836
rect 1811 2805 1823 2808
rect 1765 2799 1823 2805
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 9398 2836 9404 2848
rect 9359 2808 9404 2836
rect 9398 2796 9404 2808
rect 9456 2796 9462 2848
rect 38194 2836 38200 2848
rect 38155 2808 38200 2836
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 3234 2632 3240 2644
rect 2915 2604 3240 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 4798 2632 4804 2644
rect 4759 2604 4804 2632
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 6733 2635 6791 2641
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 7282 2632 7288 2644
rect 6779 2604 7288 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 9858 2632 9864 2644
rect 8067 2604 9864 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 10100 2604 10425 2632
rect 10100 2592 10106 2604
rect 10413 2601 10425 2604
rect 10459 2601 10471 2635
rect 10413 2595 10471 2601
rect 14274 2592 14280 2644
rect 14332 2632 14338 2644
rect 14461 2635 14519 2641
rect 14461 2632 14473 2635
rect 14332 2604 14473 2632
rect 14332 2592 14338 2604
rect 14461 2601 14473 2604
rect 14507 2601 14519 2635
rect 14461 2595 14519 2601
rect 15470 2592 15476 2644
rect 15528 2632 15534 2644
rect 15565 2635 15623 2641
rect 15565 2632 15577 2635
rect 15528 2604 15577 2632
rect 15528 2592 15534 2604
rect 15565 2601 15577 2604
rect 15611 2601 15623 2635
rect 15565 2595 15623 2601
rect 16942 2592 16948 2644
rect 17000 2632 17006 2644
rect 17037 2635 17095 2641
rect 17037 2632 17049 2635
rect 17000 2604 17049 2632
rect 17000 2592 17006 2604
rect 17037 2601 17049 2604
rect 17083 2601 17095 2635
rect 17037 2595 17095 2601
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 20496 2604 22017 2632
rect 20496 2592 20502 2604
rect 22005 2601 22017 2604
rect 22051 2601 22063 2635
rect 22005 2595 22063 2601
rect 23382 2592 23388 2644
rect 23440 2632 23446 2644
rect 24581 2635 24639 2641
rect 24581 2632 24593 2635
rect 23440 2604 24593 2632
rect 23440 2592 23446 2604
rect 24581 2601 24593 2604
rect 24627 2601 24639 2635
rect 24581 2595 24639 2601
rect 25406 2592 25412 2644
rect 25464 2632 25470 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 25464 2604 27169 2632
rect 25464 2592 25470 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 29730 2632 29736 2644
rect 29691 2604 29736 2632
rect 27157 2595 27215 2601
rect 29730 2592 29736 2604
rect 29788 2592 29794 2644
rect 30282 2592 30288 2644
rect 30340 2632 30346 2644
rect 32309 2635 32367 2641
rect 32309 2632 32321 2635
rect 30340 2604 32321 2632
rect 30340 2592 30346 2604
rect 32309 2601 32321 2604
rect 32355 2601 32367 2635
rect 32309 2595 32367 2601
rect 34330 2592 34336 2644
rect 34388 2632 34394 2644
rect 36725 2635 36783 2641
rect 36725 2632 36737 2635
rect 34388 2604 36737 2632
rect 34388 2592 34394 2604
rect 36725 2601 36737 2604
rect 36771 2601 36783 2635
rect 36725 2595 36783 2601
rect 4614 2524 4620 2576
rect 4672 2524 4678 2576
rect 30558 2524 30564 2576
rect 30616 2564 30622 2576
rect 34885 2567 34943 2573
rect 34885 2564 34897 2567
rect 30616 2536 34897 2564
rect 30616 2524 30622 2536
rect 34885 2533 34897 2536
rect 34931 2533 34943 2567
rect 34885 2527 34943 2533
rect 4632 2496 4660 2524
rect 12618 2496 12624 2508
rect 1872 2468 4660 2496
rect 12579 2468 12624 2496
rect 1872 2437 1900 2468
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 34422 2456 34428 2508
rect 34480 2496 34486 2508
rect 34480 2468 37504 2496
rect 34480 2456 34486 2468
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 2685 2431 2743 2437
rect 2685 2428 2697 2431
rect 2648 2400 2697 2428
rect 2648 2388 2654 2400
rect 2685 2397 2697 2400
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5868 2400 6561 2428
rect 5868 2388 5874 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7800 2400 7849 2428
rect 7800 2388 7806 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 9398 2428 9404 2440
rect 9359 2400 9404 2428
rect 7837 2391 7895 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12308 2400 12357 2428
rect 12308 2388 12314 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13596 2400 14289 2428
rect 13596 2388 13602 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15528 2400 15761 2428
rect 15528 2388 15534 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 18598 2428 18604 2440
rect 18559 2400 18604 2428
rect 16853 2391 16911 2397
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21324 2400 22201 2428
rect 21324 2388 21330 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 23290 2428 23296 2440
rect 23251 2400 23296 2428
rect 22189 2391 22247 2397
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24544 2400 24777 2428
rect 24544 2388 24550 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 26476 2400 27353 2428
rect 26476 2388 26482 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27798 2428 27804 2440
rect 27759 2400 27804 2428
rect 27341 2391 27399 2397
rect 27798 2388 27804 2400
rect 27856 2388 27862 2440
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 30006 2388 30012 2440
rect 30064 2428 30070 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30064 2400 31033 2428
rect 30064 2388 30070 2400
rect 31021 2397 31033 2400
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 32272 2400 32505 2428
rect 32272 2388 32278 2400
rect 32493 2397 32505 2400
rect 32539 2397 32551 2431
rect 32493 2391 32551 2397
rect 34146 2388 34152 2440
rect 34204 2428 34210 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34204 2400 35081 2428
rect 34204 2388 34210 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35069 2391 35127 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 37476 2437 37504 2468
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 36909 2431 36967 2437
rect 36909 2397 36921 2431
rect 36955 2397 36967 2431
rect 36909 2391 36967 2397
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 36924 2360 36952 2391
rect 38654 2360 38660 2372
rect 36924 2332 38660 2360
rect 38654 2320 38660 2332
rect 38712 2320 38718 2372
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 72 2264 1685 2292
rect 72 2252 78 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 9088 2264 9229 2292
rect 9088 2252 9094 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18748 2264 18797 2292
rect 18748 2252 18754 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 18785 2255 18843 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 20036 2264 20269 2292
rect 20036 2252 20042 2264
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23256 2264 23489 2292
rect 23256 2252 23262 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 27985 2295 28043 2301
rect 27985 2292 27997 2295
rect 27764 2264 27997 2292
rect 27764 2252 27770 2264
rect 27985 2261 27997 2264
rect 28031 2261 28043 2295
rect 27985 2255 28043 2261
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 30984 2264 31217 2292
rect 30984 2252 30990 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 33042 2252 33048 2304
rect 33100 2292 33106 2304
rect 35529 2295 35587 2301
rect 35529 2292 35541 2295
rect 33100 2264 35541 2292
rect 33100 2252 33106 2264
rect 35529 2261 35541 2264
rect 35575 2261 35587 2295
rect 35529 2255 35587 2261
rect 37366 2252 37372 2304
rect 37424 2292 37430 2304
rect 37645 2295 37703 2301
rect 37645 2292 37657 2295
rect 37424 2264 37657 2292
rect 37424 2252 37430 2264
rect 37645 2261 37657 2264
rect 37691 2261 37703 2295
rect 37645 2255 37703 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1860 37247 1912 37256
rect 1860 37213 1869 37247
rect 1869 37213 1903 37247
rect 1903 37213 1912 37247
rect 1860 37204 1912 37213
rect 1952 37204 2004 37256
rect 2964 37247 3016 37256
rect 2964 37213 2973 37247
rect 2973 37213 3007 37247
rect 3007 37213 3016 37247
rect 2964 37204 3016 37213
rect 4252 37247 4304 37256
rect 4252 37213 4261 37247
rect 4261 37213 4295 37247
rect 4295 37213 4304 37247
rect 4252 37204 4304 37213
rect 5540 37247 5592 37256
rect 5540 37213 5549 37247
rect 5549 37213 5583 37247
rect 5583 37213 5592 37247
rect 5540 37204 5592 37213
rect 7104 37204 7156 37256
rect 8392 37204 8444 37256
rect 10324 37204 10376 37256
rect 11612 37204 11664 37256
rect 12900 37204 12952 37256
rect 15200 37247 15252 37256
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 18144 37247 18196 37256
rect 18144 37213 18153 37247
rect 18153 37213 18187 37247
rect 18187 37213 18196 37247
rect 18144 37204 18196 37213
rect 18236 37204 18288 37256
rect 20720 37204 20772 37256
rect 22560 37204 22612 37256
rect 22928 37204 22980 37256
rect 24768 37204 24820 37256
rect 27068 37204 27120 37256
rect 27436 37204 27488 37256
rect 30380 37204 30432 37256
rect 31760 37204 31812 37256
rect 33508 37204 33560 37256
rect 34796 37204 34848 37256
rect 36728 37204 36780 37256
rect 2780 37136 2832 37188
rect 6552 37136 6604 37188
rect 19984 37136 20036 37188
rect 3148 37111 3200 37120
rect 3148 37077 3157 37111
rect 3157 37077 3191 37111
rect 3191 37077 3200 37111
rect 3148 37068 3200 37077
rect 3884 37068 3936 37120
rect 5172 37068 5224 37120
rect 7196 37111 7248 37120
rect 7196 37077 7205 37111
rect 7205 37077 7239 37111
rect 7239 37077 7248 37111
rect 7196 37068 7248 37077
rect 8300 37068 8352 37120
rect 10324 37068 10376 37120
rect 10876 37068 10928 37120
rect 14740 37068 14792 37120
rect 14832 37068 14884 37120
rect 16580 37068 16632 37120
rect 18052 37068 18104 37120
rect 19340 37068 19392 37120
rect 20720 37111 20772 37120
rect 20720 37077 20729 37111
rect 20729 37077 20763 37111
rect 20763 37077 20772 37111
rect 20720 37068 20772 37077
rect 29368 37136 29420 37188
rect 23848 37068 23900 37120
rect 25780 37068 25832 37120
rect 27160 37111 27212 37120
rect 27160 37077 27169 37111
rect 27169 37077 27203 37111
rect 27203 37077 27212 37111
rect 27160 37068 27212 37077
rect 29000 37068 29052 37120
rect 30472 37111 30524 37120
rect 30472 37077 30481 37111
rect 30481 37077 30515 37111
rect 30515 37077 30524 37111
rect 30472 37068 30524 37077
rect 32312 37111 32364 37120
rect 32312 37077 32321 37111
rect 32321 37077 32355 37111
rect 32355 37077 32364 37111
rect 32312 37068 32364 37077
rect 33968 37136 34020 37188
rect 34888 37111 34940 37120
rect 34888 37077 34897 37111
rect 34897 37077 34931 37111
rect 34931 37077 34940 37111
rect 34888 37068 34940 37077
rect 35900 37068 35952 37120
rect 38200 37111 38252 37120
rect 38200 37077 38209 37111
rect 38209 37077 38243 37111
rect 38243 37077 38252 37111
rect 38200 37068 38252 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 664 36864 716 36916
rect 1860 36864 1912 36916
rect 3976 36864 4028 36916
rect 30288 36864 30340 36916
rect 34888 36864 34940 36916
rect 4068 36728 4120 36780
rect 39304 36796 39356 36848
rect 37556 36771 37608 36780
rect 37556 36737 37565 36771
rect 37565 36737 37599 36771
rect 37599 36737 37608 36771
rect 37556 36728 37608 36737
rect 36728 36567 36780 36576
rect 36728 36533 36737 36567
rect 36737 36533 36771 36567
rect 36771 36533 36780 36567
rect 36728 36524 36780 36533
rect 37372 36524 37424 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 37188 36320 37240 36372
rect 1584 36159 1636 36168
rect 1584 36125 1593 36159
rect 1593 36125 1627 36159
rect 1627 36125 1636 36159
rect 1584 36116 1636 36125
rect 37372 36159 37424 36168
rect 37372 36125 37381 36159
rect 37381 36125 37415 36159
rect 37415 36125 37424 36159
rect 37372 36116 37424 36125
rect 6644 35980 6696 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 5540 35776 5592 35828
rect 16856 35819 16908 35828
rect 16856 35785 16865 35819
rect 16865 35785 16899 35819
rect 16899 35785 16908 35819
rect 16856 35776 16908 35785
rect 5908 35683 5960 35692
rect 5908 35649 5917 35683
rect 5917 35649 5951 35683
rect 5951 35649 5960 35683
rect 5908 35640 5960 35649
rect 17040 35683 17092 35692
rect 17040 35649 17049 35683
rect 17049 35649 17083 35683
rect 17083 35649 17092 35683
rect 17040 35640 17092 35649
rect 38016 35640 38068 35692
rect 33232 35436 33284 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3976 35232 4028 35284
rect 18144 35232 18196 35284
rect 18236 35164 18288 35216
rect 6736 35028 6788 35080
rect 16488 35028 16540 35080
rect 17500 35071 17552 35080
rect 17500 35037 17509 35071
rect 17509 35037 17543 35071
rect 17543 35037 17552 35071
rect 17500 35028 17552 35037
rect 35348 35028 35400 35080
rect 38200 34935 38252 34944
rect 38200 34901 38209 34935
rect 38209 34901 38243 34935
rect 38243 34901 38252 34935
rect 38200 34892 38252 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4068 34688 4120 34740
rect 15200 34688 15252 34740
rect 20076 34620 20128 34672
rect 24768 34688 24820 34740
rect 27436 34688 27488 34740
rect 3976 34552 4028 34604
rect 12072 34552 12124 34604
rect 14740 34552 14792 34604
rect 15660 34595 15712 34604
rect 15660 34561 15669 34595
rect 15669 34561 15703 34595
rect 15703 34561 15712 34595
rect 15660 34552 15712 34561
rect 20720 34595 20772 34604
rect 20720 34561 20729 34595
rect 20729 34561 20763 34595
rect 20763 34561 20772 34595
rect 20720 34552 20772 34561
rect 22928 34620 22980 34672
rect 21272 34552 21324 34604
rect 24676 34552 24728 34604
rect 33232 34595 33284 34604
rect 33232 34561 33241 34595
rect 33241 34561 33275 34595
rect 33275 34561 33284 34595
rect 33232 34552 33284 34561
rect 16120 34484 16172 34536
rect 20352 34484 20404 34536
rect 33140 34527 33192 34536
rect 33140 34493 33149 34527
rect 33149 34493 33183 34527
rect 33183 34493 33192 34527
rect 33140 34484 33192 34493
rect 1676 34391 1728 34400
rect 1676 34357 1685 34391
rect 1685 34357 1719 34391
rect 1719 34357 1728 34391
rect 1676 34348 1728 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 10876 34008 10928 34060
rect 10324 33983 10376 33992
rect 10324 33949 10333 33983
rect 10333 33949 10367 33983
rect 10367 33949 10376 33983
rect 10324 33940 10376 33949
rect 30288 33983 30340 33992
rect 30288 33949 30297 33983
rect 30297 33949 30331 33983
rect 30331 33949 30340 33983
rect 30288 33940 30340 33949
rect 8392 33804 8444 33856
rect 10232 33804 10284 33856
rect 18788 33804 18840 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 15660 33600 15712 33652
rect 13544 33464 13596 33516
rect 19984 33507 20036 33516
rect 19984 33473 19993 33507
rect 19993 33473 20027 33507
rect 20027 33473 20036 33507
rect 19984 33464 20036 33473
rect 29368 33507 29420 33516
rect 29368 33473 29377 33507
rect 29377 33473 29411 33507
rect 29411 33473 29420 33507
rect 29368 33464 29420 33473
rect 33508 33464 33560 33516
rect 12164 33328 12216 33380
rect 38200 33371 38252 33380
rect 38200 33337 38209 33371
rect 38209 33337 38243 33371
rect 38243 33337 38252 33371
rect 38200 33328 38252 33337
rect 17592 33260 17644 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1584 32895 1636 32904
rect 1584 32861 1593 32895
rect 1593 32861 1627 32895
rect 1627 32861 1636 32895
rect 1584 32852 1636 32861
rect 4620 32716 4672 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 33968 32555 34020 32564
rect 33968 32521 33977 32555
rect 33977 32521 34011 32555
rect 34011 32521 34020 32555
rect 33968 32512 34020 32521
rect 3148 32376 3200 32428
rect 33232 32376 33284 32428
rect 6184 32172 6236 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 33784 31900 33836 31952
rect 18972 31764 19024 31816
rect 27160 31764 27212 31816
rect 38292 31807 38344 31816
rect 38292 31773 38301 31807
rect 38301 31773 38335 31807
rect 38335 31773 38344 31807
rect 38292 31764 38344 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 17040 31424 17092 31476
rect 16672 31288 16724 31340
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3976 30923 4028 30932
rect 3976 30889 3985 30923
rect 3985 30889 4019 30923
rect 4019 30889 4028 30923
rect 3976 30880 4028 30889
rect 5908 30880 5960 30932
rect 35348 30880 35400 30932
rect 9128 30812 9180 30864
rect 1584 30719 1636 30728
rect 1584 30685 1593 30719
rect 1593 30685 1627 30719
rect 1627 30685 1636 30719
rect 1584 30676 1636 30685
rect 4068 30676 4120 30728
rect 6276 30719 6328 30728
rect 6276 30685 6285 30719
rect 6285 30685 6319 30719
rect 6319 30685 6328 30719
rect 6276 30676 6328 30685
rect 8300 30719 8352 30728
rect 8300 30685 8309 30719
rect 8309 30685 8343 30719
rect 8343 30685 8352 30719
rect 8300 30676 8352 30685
rect 33876 30676 33928 30728
rect 8208 30583 8260 30592
rect 8208 30549 8217 30583
rect 8217 30549 8251 30583
rect 8251 30549 8260 30583
rect 8208 30540 8260 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 6736 30268 6788 30320
rect 21272 30268 21324 30320
rect 2964 30200 3016 30252
rect 6552 30243 6604 30252
rect 6552 30209 6561 30243
rect 6561 30209 6595 30243
rect 6595 30209 6604 30243
rect 6552 30200 6604 30209
rect 12992 30200 13044 30252
rect 17132 30200 17184 30252
rect 35900 30268 35952 30320
rect 33324 30243 33376 30252
rect 2228 30132 2280 30184
rect 33324 30209 33333 30243
rect 33333 30209 33367 30243
rect 33367 30209 33376 30243
rect 33324 30200 33376 30209
rect 38292 30243 38344 30252
rect 38292 30209 38301 30243
rect 38301 30209 38335 30243
rect 38335 30209 38344 30243
rect 38292 30200 38344 30209
rect 32312 30132 32364 30184
rect 33508 30107 33560 30116
rect 33508 30073 33517 30107
rect 33517 30073 33551 30107
rect 33551 30073 33560 30107
rect 33508 30064 33560 30073
rect 7748 29996 7800 30048
rect 27252 30039 27304 30048
rect 27252 30005 27261 30039
rect 27261 30005 27295 30039
rect 27295 30005 27304 30039
rect 27252 29996 27304 30005
rect 29184 30039 29236 30048
rect 29184 30005 29193 30039
rect 29193 30005 29227 30039
rect 29227 30005 29236 30039
rect 29184 29996 29236 30005
rect 35440 29996 35492 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 12072 29835 12124 29844
rect 12072 29801 12081 29835
rect 12081 29801 12115 29835
rect 12115 29801 12124 29835
rect 12072 29792 12124 29801
rect 16488 29835 16540 29844
rect 16488 29801 16497 29835
rect 16497 29801 16531 29835
rect 16531 29801 16540 29835
rect 16488 29792 16540 29801
rect 17500 29792 17552 29844
rect 24676 29835 24728 29844
rect 24676 29801 24685 29835
rect 24685 29801 24719 29835
rect 24719 29801 24728 29835
rect 24676 29792 24728 29801
rect 2596 29699 2648 29708
rect 2596 29665 2605 29699
rect 2605 29665 2639 29699
rect 2639 29665 2648 29699
rect 2596 29656 2648 29665
rect 9864 29656 9916 29708
rect 2964 29588 3016 29640
rect 4988 29588 5040 29640
rect 3608 29520 3660 29572
rect 7472 29520 7524 29572
rect 14648 29588 14700 29640
rect 17040 29631 17092 29640
rect 17040 29597 17049 29631
rect 17049 29597 17083 29631
rect 17083 29597 17092 29631
rect 17040 29588 17092 29597
rect 23388 29588 23440 29640
rect 30472 29588 30524 29640
rect 36728 29588 36780 29640
rect 15384 29520 15436 29572
rect 1676 29495 1728 29504
rect 1676 29461 1685 29495
rect 1685 29461 1719 29495
rect 1719 29461 1728 29495
rect 1676 29452 1728 29461
rect 8024 29452 8076 29504
rect 25412 29495 25464 29504
rect 25412 29461 25421 29495
rect 25421 29461 25455 29495
rect 25455 29461 25464 29495
rect 25412 29452 25464 29461
rect 30472 29495 30524 29504
rect 30472 29461 30481 29495
rect 30481 29461 30515 29495
rect 30515 29461 30524 29495
rect 30472 29452 30524 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1584 29155 1636 29164
rect 1584 29121 1593 29155
rect 1593 29121 1627 29155
rect 1627 29121 1636 29155
rect 1584 29112 1636 29121
rect 4620 29112 4672 29164
rect 4988 29155 5040 29164
rect 2320 29044 2372 29096
rect 2964 29044 3016 29096
rect 4988 29121 4997 29155
rect 4997 29121 5031 29155
rect 5031 29121 5040 29155
rect 4988 29112 5040 29121
rect 38016 29155 38068 29164
rect 38016 29121 38025 29155
rect 38025 29121 38059 29155
rect 38059 29121 38068 29155
rect 38016 29112 38068 29121
rect 5080 29087 5132 29096
rect 5080 29053 5089 29087
rect 5089 29053 5123 29087
rect 5123 29053 5132 29087
rect 5080 29044 5132 29053
rect 3884 28976 3936 29028
rect 5356 28976 5408 29028
rect 38200 29019 38252 29028
rect 38200 28985 38209 29019
rect 38209 28985 38243 29019
rect 38243 28985 38252 29019
rect 38200 28976 38252 28985
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4068 28747 4120 28756
rect 4068 28713 4077 28747
rect 4077 28713 4111 28747
rect 4111 28713 4120 28747
rect 4068 28704 4120 28713
rect 20076 28704 20128 28756
rect 33324 28704 33376 28756
rect 2964 28500 3016 28552
rect 4896 28500 4948 28552
rect 15660 28500 15712 28552
rect 16304 28543 16356 28552
rect 16304 28509 16313 28543
rect 16313 28509 16347 28543
rect 16347 28509 16356 28543
rect 16304 28500 16356 28509
rect 19064 28500 19116 28552
rect 33324 28543 33376 28552
rect 33324 28509 33333 28543
rect 33333 28509 33367 28543
rect 33367 28509 33376 28543
rect 33324 28500 33376 28509
rect 35440 28500 35492 28552
rect 2504 28432 2556 28484
rect 17684 28364 17736 28416
rect 34060 28407 34112 28416
rect 34060 28373 34069 28407
rect 34069 28373 34103 28407
rect 34103 28373 34112 28407
rect 34060 28364 34112 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 18696 28160 18748 28212
rect 34060 28160 34112 28212
rect 2228 28024 2280 28076
rect 4068 28024 4120 28076
rect 6644 28024 6696 28076
rect 15844 28067 15896 28076
rect 15844 28033 15853 28067
rect 15853 28033 15887 28067
rect 15887 28033 15896 28067
rect 15844 28024 15896 28033
rect 16304 28024 16356 28076
rect 33784 28067 33836 28076
rect 33784 28033 33793 28067
rect 33793 28033 33827 28067
rect 33827 28033 33836 28067
rect 33784 28024 33836 28033
rect 2044 27863 2096 27872
rect 2044 27829 2053 27863
rect 2053 27829 2087 27863
rect 2087 27829 2096 27863
rect 2044 27820 2096 27829
rect 2688 27863 2740 27872
rect 2688 27829 2697 27863
rect 2697 27829 2731 27863
rect 2731 27829 2740 27863
rect 2688 27820 2740 27829
rect 3976 27820 4028 27872
rect 4988 27820 5040 27872
rect 7932 27820 7984 27872
rect 15936 27820 15988 27872
rect 16948 27863 17000 27872
rect 16948 27829 16957 27863
rect 16957 27829 16991 27863
rect 16991 27829 17000 27863
rect 16948 27820 17000 27829
rect 20720 27820 20772 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 16672 27591 16724 27600
rect 16672 27557 16681 27591
rect 16681 27557 16715 27591
rect 16715 27557 16724 27591
rect 16672 27548 16724 27557
rect 7104 27480 7156 27532
rect 2228 27412 2280 27464
rect 2320 27344 2372 27396
rect 4068 27412 4120 27464
rect 6828 27344 6880 27396
rect 1768 27276 1820 27328
rect 2872 27319 2924 27328
rect 2872 27285 2881 27319
rect 2881 27285 2915 27319
rect 2915 27285 2924 27319
rect 2872 27276 2924 27285
rect 3516 27276 3568 27328
rect 5632 27276 5684 27328
rect 5908 27319 5960 27328
rect 5908 27285 5917 27319
rect 5917 27285 5951 27319
rect 5951 27285 5960 27319
rect 5908 27276 5960 27285
rect 6092 27276 6144 27328
rect 7288 27412 7340 27464
rect 9128 27455 9180 27464
rect 9128 27421 9137 27455
rect 9137 27421 9171 27455
rect 9171 27421 9180 27455
rect 9128 27412 9180 27421
rect 12624 27412 12676 27464
rect 15936 27455 15988 27464
rect 15936 27421 15945 27455
rect 15945 27421 15979 27455
rect 15979 27421 15988 27455
rect 15936 27412 15988 27421
rect 17684 27455 17736 27464
rect 17684 27421 17693 27455
rect 17693 27421 17727 27455
rect 17727 27421 17736 27455
rect 17684 27412 17736 27421
rect 9220 27319 9272 27328
rect 9220 27285 9229 27319
rect 9229 27285 9263 27319
rect 9263 27285 9272 27319
rect 9220 27276 9272 27285
rect 12256 27276 12308 27328
rect 15752 27319 15804 27328
rect 15752 27285 15761 27319
rect 15761 27285 15795 27319
rect 15795 27285 15804 27319
rect 15752 27276 15804 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 3608 27115 3660 27124
rect 3608 27081 3617 27115
rect 3617 27081 3651 27115
rect 3651 27081 3660 27115
rect 3608 27072 3660 27081
rect 6276 27072 6328 27124
rect 16672 27072 16724 27124
rect 33232 27072 33284 27124
rect 4068 27004 4120 27056
rect 20 26936 72 26988
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 3792 26979 3844 26988
rect 3792 26945 3801 26979
rect 3801 26945 3835 26979
rect 3835 26945 3844 26979
rect 3792 26936 3844 26945
rect 4804 26936 4856 26988
rect 7288 26936 7340 26988
rect 9036 26936 9088 26988
rect 12624 26979 12676 26988
rect 5448 26868 5500 26920
rect 7656 26868 7708 26920
rect 8576 26868 8628 26920
rect 12624 26945 12633 26979
rect 12633 26945 12667 26979
rect 12667 26945 12676 26979
rect 12624 26936 12676 26945
rect 12440 26800 12492 26852
rect 15476 26911 15528 26920
rect 15476 26877 15485 26911
rect 15485 26877 15519 26911
rect 15519 26877 15528 26911
rect 15476 26868 15528 26877
rect 16948 26936 17000 26988
rect 17224 26868 17276 26920
rect 18144 26868 18196 26920
rect 20076 26936 20128 26988
rect 29736 26979 29788 26988
rect 29736 26945 29745 26979
rect 29745 26945 29779 26979
rect 29779 26945 29788 26979
rect 29736 26936 29788 26945
rect 35348 26936 35400 26988
rect 19432 26868 19484 26920
rect 1860 26732 1912 26784
rect 2504 26732 2556 26784
rect 3148 26732 3200 26784
rect 4712 26732 4764 26784
rect 5080 26732 5132 26784
rect 9956 26732 10008 26784
rect 13360 26732 13412 26784
rect 13636 26732 13688 26784
rect 14832 26732 14884 26784
rect 15200 26732 15252 26784
rect 15568 26732 15620 26784
rect 17684 26732 17736 26784
rect 18880 26775 18932 26784
rect 18880 26741 18889 26775
rect 18889 26741 18923 26775
rect 18923 26741 18932 26775
rect 18880 26732 18932 26741
rect 38200 26775 38252 26784
rect 38200 26741 38209 26775
rect 38209 26741 38243 26775
rect 38243 26741 38252 26775
rect 38200 26732 38252 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 4804 26528 4856 26580
rect 6276 26571 6328 26580
rect 6276 26537 6285 26571
rect 6285 26537 6319 26571
rect 6319 26537 6328 26571
rect 6276 26528 6328 26537
rect 18144 26571 18196 26580
rect 8208 26460 8260 26512
rect 5908 26435 5960 26444
rect 5908 26401 5917 26435
rect 5917 26401 5951 26435
rect 5951 26401 5960 26435
rect 5908 26392 5960 26401
rect 6092 26435 6144 26444
rect 6092 26401 6101 26435
rect 6101 26401 6135 26435
rect 6135 26401 6144 26435
rect 6092 26392 6144 26401
rect 13544 26460 13596 26512
rect 17592 26460 17644 26512
rect 18144 26537 18153 26571
rect 18153 26537 18187 26571
rect 18187 26537 18196 26571
rect 18144 26528 18196 26537
rect 20444 26528 20496 26580
rect 38016 26528 38068 26580
rect 14280 26392 14332 26444
rect 14464 26392 14516 26444
rect 2320 26367 2372 26376
rect 2320 26333 2329 26367
rect 2329 26333 2363 26367
rect 2363 26333 2372 26367
rect 2320 26324 2372 26333
rect 2964 26324 3016 26376
rect 1952 26256 2004 26308
rect 4068 26256 4120 26308
rect 4804 26324 4856 26376
rect 8208 26367 8260 26376
rect 8208 26333 8217 26367
rect 8217 26333 8251 26367
rect 8251 26333 8260 26367
rect 8208 26324 8260 26333
rect 9036 26324 9088 26376
rect 9956 26367 10008 26376
rect 9956 26333 9965 26367
rect 9965 26333 9999 26367
rect 9999 26333 10008 26367
rect 9956 26324 10008 26333
rect 10968 26367 11020 26376
rect 10968 26333 10977 26367
rect 10977 26333 11011 26367
rect 11011 26333 11020 26367
rect 10968 26324 11020 26333
rect 12072 26324 12124 26376
rect 12256 26367 12308 26376
rect 12256 26333 12265 26367
rect 12265 26333 12299 26367
rect 12299 26333 12308 26367
rect 12256 26324 12308 26333
rect 12532 26324 12584 26376
rect 15568 26367 15620 26376
rect 11060 26299 11112 26308
rect 11060 26265 11069 26299
rect 11069 26265 11103 26299
rect 11103 26265 11112 26299
rect 11060 26256 11112 26265
rect 11888 26256 11940 26308
rect 12900 26256 12952 26308
rect 15568 26333 15577 26367
rect 15577 26333 15611 26367
rect 15611 26333 15620 26367
rect 15568 26324 15620 26333
rect 17224 26392 17276 26444
rect 17684 26367 17736 26376
rect 17684 26333 17693 26367
rect 17693 26333 17727 26367
rect 17727 26333 17736 26367
rect 17684 26324 17736 26333
rect 18788 26435 18840 26444
rect 18788 26401 18797 26435
rect 18797 26401 18831 26435
rect 18831 26401 18840 26435
rect 18788 26392 18840 26401
rect 36084 26367 36136 26376
rect 15108 26256 15160 26308
rect 36084 26333 36093 26367
rect 36093 26333 36127 26367
rect 36127 26333 36136 26367
rect 36084 26324 36136 26333
rect 20628 26256 20680 26308
rect 4344 26231 4396 26240
rect 4344 26197 4353 26231
rect 4353 26197 4387 26231
rect 4387 26197 4396 26231
rect 4344 26188 4396 26197
rect 5172 26188 5224 26240
rect 7656 26188 7708 26240
rect 9772 26231 9824 26240
rect 9772 26197 9781 26231
rect 9781 26197 9815 26231
rect 9815 26197 9824 26231
rect 9772 26188 9824 26197
rect 12716 26188 12768 26240
rect 13728 26231 13780 26240
rect 13728 26197 13737 26231
rect 13737 26197 13771 26231
rect 13771 26197 13780 26231
rect 13728 26188 13780 26197
rect 16028 26188 16080 26240
rect 16212 26231 16264 26240
rect 16212 26197 16221 26231
rect 16221 26197 16255 26231
rect 16255 26197 16264 26231
rect 16212 26188 16264 26197
rect 19340 26188 19392 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 3792 26027 3844 26036
rect 3792 25993 3801 26027
rect 3801 25993 3835 26027
rect 3835 25993 3844 26027
rect 3792 25984 3844 25993
rect 7656 26027 7708 26036
rect 7656 25993 7665 26027
rect 7665 25993 7699 26027
rect 7699 25993 7708 26027
rect 7656 25984 7708 25993
rect 12348 25984 12400 26036
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 2228 25848 2280 25900
rect 4344 25916 4396 25968
rect 4804 25848 4856 25900
rect 1308 25712 1360 25764
rect 6828 25916 6880 25968
rect 7012 25848 7064 25900
rect 7380 25848 7432 25900
rect 8392 25848 8444 25900
rect 12440 25916 12492 25968
rect 10232 25891 10284 25900
rect 10232 25857 10241 25891
rect 10241 25857 10275 25891
rect 10275 25857 10284 25891
rect 10232 25848 10284 25857
rect 10324 25848 10376 25900
rect 10968 25848 11020 25900
rect 6828 25780 6880 25832
rect 9772 25780 9824 25832
rect 10048 25823 10100 25832
rect 10048 25789 10057 25823
rect 10057 25789 10091 25823
rect 10091 25789 10100 25823
rect 10048 25780 10100 25789
rect 11612 25848 11664 25900
rect 12624 25848 12676 25900
rect 13728 25916 13780 25968
rect 13176 25891 13228 25900
rect 13176 25857 13185 25891
rect 13185 25857 13219 25891
rect 13219 25857 13228 25891
rect 13176 25848 13228 25857
rect 15844 25984 15896 26036
rect 19432 25984 19484 26036
rect 20076 26027 20128 26036
rect 20076 25993 20085 26027
rect 20085 25993 20119 26027
rect 20119 25993 20128 26027
rect 20076 25984 20128 25993
rect 20628 25984 20680 26036
rect 33876 25984 33928 26036
rect 12808 25780 12860 25832
rect 15936 25848 15988 25900
rect 17500 25891 17552 25900
rect 17500 25857 17509 25891
rect 17509 25857 17543 25891
rect 17543 25857 17552 25891
rect 17500 25848 17552 25857
rect 19340 25848 19392 25900
rect 18696 25823 18748 25832
rect 18696 25789 18705 25823
rect 18705 25789 18739 25823
rect 18739 25789 18748 25823
rect 18696 25780 18748 25789
rect 19524 25780 19576 25832
rect 5908 25712 5960 25764
rect 1860 25644 1912 25696
rect 3240 25644 3292 25696
rect 4620 25644 4672 25696
rect 5540 25644 5592 25696
rect 6460 25644 6512 25696
rect 8668 25644 8720 25696
rect 9680 25644 9732 25696
rect 11704 25712 11756 25764
rect 11980 25644 12032 25696
rect 12348 25687 12400 25696
rect 12348 25653 12357 25687
rect 12357 25653 12391 25687
rect 12391 25653 12400 25687
rect 12348 25644 12400 25653
rect 12440 25644 12492 25696
rect 16396 25712 16448 25764
rect 16488 25712 16540 25764
rect 24032 25848 24084 25900
rect 13820 25644 13872 25696
rect 14740 25687 14792 25696
rect 14740 25653 14749 25687
rect 14749 25653 14783 25687
rect 14783 25653 14792 25687
rect 14740 25644 14792 25653
rect 16764 25644 16816 25696
rect 16856 25687 16908 25696
rect 16856 25653 16865 25687
rect 16865 25653 16899 25687
rect 16899 25653 16908 25687
rect 16856 25644 16908 25653
rect 18512 25644 18564 25696
rect 20536 25644 20588 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 4068 25440 4120 25492
rect 8116 25372 8168 25424
rect 10048 25440 10100 25492
rect 10416 25440 10468 25492
rect 13176 25440 13228 25492
rect 9772 25372 9824 25424
rect 14556 25440 14608 25492
rect 18144 25483 18196 25492
rect 18144 25449 18153 25483
rect 18153 25449 18187 25483
rect 18187 25449 18196 25483
rect 18144 25440 18196 25449
rect 36084 25440 36136 25492
rect 3700 25304 3752 25356
rect 1860 25279 1912 25288
rect 1860 25245 1869 25279
rect 1869 25245 1903 25279
rect 1903 25245 1912 25279
rect 1860 25236 1912 25245
rect 2412 25236 2464 25288
rect 5172 25279 5224 25288
rect 3056 25168 3108 25220
rect 2136 25100 2188 25152
rect 5172 25245 5181 25279
rect 5181 25245 5215 25279
rect 5215 25245 5224 25279
rect 5172 25236 5224 25245
rect 5816 25279 5868 25288
rect 5816 25245 5825 25279
rect 5825 25245 5859 25279
rect 5859 25245 5868 25279
rect 5816 25236 5868 25245
rect 6460 25279 6512 25288
rect 6460 25245 6469 25279
rect 6469 25245 6503 25279
rect 6503 25245 6512 25279
rect 6460 25236 6512 25245
rect 7380 25236 7432 25288
rect 6276 25168 6328 25220
rect 6828 25168 6880 25220
rect 8576 25279 8628 25288
rect 8576 25245 8585 25279
rect 8585 25245 8619 25279
rect 8619 25245 8628 25279
rect 8576 25236 8628 25245
rect 8760 25236 8812 25288
rect 12992 25347 13044 25356
rect 12992 25313 13001 25347
rect 13001 25313 13035 25347
rect 13035 25313 13044 25347
rect 12992 25304 13044 25313
rect 15200 25347 15252 25356
rect 15200 25313 15209 25347
rect 15209 25313 15243 25347
rect 15243 25313 15252 25347
rect 15200 25304 15252 25313
rect 16212 25304 16264 25356
rect 18880 25304 18932 25356
rect 9496 25168 9548 25220
rect 12716 25236 12768 25288
rect 15016 25279 15068 25288
rect 15016 25245 15025 25279
rect 15025 25245 15059 25279
rect 15059 25245 15068 25279
rect 15016 25236 15068 25245
rect 16028 25236 16080 25288
rect 16672 25236 16724 25288
rect 18236 25236 18288 25288
rect 18972 25236 19024 25288
rect 19524 25236 19576 25288
rect 13544 25211 13596 25220
rect 13544 25177 13553 25211
rect 13553 25177 13587 25211
rect 13587 25177 13596 25211
rect 13544 25168 13596 25177
rect 3608 25100 3660 25152
rect 5264 25143 5316 25152
rect 5264 25109 5273 25143
rect 5273 25109 5307 25143
rect 5307 25109 5316 25143
rect 5264 25100 5316 25109
rect 6552 25100 6604 25152
rect 6736 25100 6788 25152
rect 7656 25100 7708 25152
rect 7840 25143 7892 25152
rect 7840 25109 7849 25143
rect 7849 25109 7883 25143
rect 7883 25109 7892 25143
rect 7840 25100 7892 25109
rect 9312 25143 9364 25152
rect 9312 25109 9321 25143
rect 9321 25109 9355 25143
rect 9355 25109 9364 25143
rect 9312 25100 9364 25109
rect 9772 25100 9824 25152
rect 10324 25100 10376 25152
rect 10600 25143 10652 25152
rect 10600 25109 10609 25143
rect 10609 25109 10643 25143
rect 10643 25109 10652 25143
rect 10600 25100 10652 25109
rect 11152 25100 11204 25152
rect 13084 25100 13136 25152
rect 14372 25100 14424 25152
rect 17960 25100 18012 25152
rect 35624 25279 35676 25288
rect 35624 25245 35633 25279
rect 35633 25245 35667 25279
rect 35667 25245 35676 25279
rect 35624 25236 35676 25245
rect 38292 25279 38344 25288
rect 38292 25245 38301 25279
rect 38301 25245 38335 25279
rect 38335 25245 38344 25279
rect 38292 25236 38344 25245
rect 20904 25100 20956 25152
rect 34796 25100 34848 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 5816 24896 5868 24948
rect 6092 24896 6144 24948
rect 8760 24896 8812 24948
rect 9312 24896 9364 24948
rect 11796 24896 11848 24948
rect 11980 24896 12032 24948
rect 15936 24896 15988 24948
rect 5448 24828 5500 24880
rect 2412 24803 2464 24812
rect 2412 24769 2421 24803
rect 2421 24769 2455 24803
rect 2455 24769 2464 24803
rect 2412 24760 2464 24769
rect 3056 24803 3108 24812
rect 3056 24769 3065 24803
rect 3065 24769 3099 24803
rect 3099 24769 3108 24803
rect 3056 24760 3108 24769
rect 3240 24803 3292 24812
rect 3240 24769 3249 24803
rect 3249 24769 3283 24803
rect 3283 24769 3292 24803
rect 3240 24760 3292 24769
rect 4620 24760 4672 24812
rect 4896 24803 4948 24812
rect 4896 24769 4905 24803
rect 4905 24769 4939 24803
rect 4939 24769 4948 24803
rect 4896 24760 4948 24769
rect 5172 24760 5224 24812
rect 5816 24803 5868 24812
rect 5816 24769 5825 24803
rect 5825 24769 5859 24803
rect 5859 24769 5868 24803
rect 5816 24760 5868 24769
rect 3608 24692 3660 24744
rect 5448 24692 5500 24744
rect 1860 24624 1912 24676
rect 7840 24760 7892 24812
rect 7932 24735 7984 24744
rect 7932 24701 7941 24735
rect 7941 24701 7975 24735
rect 7975 24701 7984 24735
rect 8392 24760 8444 24812
rect 9680 24803 9732 24812
rect 9680 24769 9689 24803
rect 9689 24769 9723 24803
rect 9723 24769 9732 24803
rect 9680 24760 9732 24769
rect 12992 24828 13044 24880
rect 13360 24871 13412 24880
rect 13360 24837 13369 24871
rect 13369 24837 13403 24871
rect 13403 24837 13412 24871
rect 13360 24828 13412 24837
rect 18696 24871 18748 24880
rect 18696 24837 18705 24871
rect 18705 24837 18739 24871
rect 18739 24837 18748 24871
rect 18696 24828 18748 24837
rect 9956 24760 10008 24812
rect 10324 24803 10376 24812
rect 10324 24769 10333 24803
rect 10333 24769 10367 24803
rect 10367 24769 10376 24803
rect 10324 24760 10376 24769
rect 7932 24692 7984 24701
rect 8668 24692 8720 24744
rect 11152 24735 11204 24744
rect 11152 24701 11161 24735
rect 11161 24701 11195 24735
rect 11195 24701 11204 24735
rect 11152 24692 11204 24701
rect 11980 24760 12032 24812
rect 13636 24760 13688 24812
rect 15476 24760 15528 24812
rect 15752 24803 15804 24812
rect 15752 24769 15761 24803
rect 15761 24769 15795 24803
rect 15795 24769 15804 24803
rect 15752 24760 15804 24769
rect 16764 24760 16816 24812
rect 17684 24760 17736 24812
rect 18420 24760 18472 24812
rect 20536 24803 20588 24812
rect 20536 24769 20545 24803
rect 20545 24769 20579 24803
rect 20579 24769 20588 24803
rect 20536 24760 20588 24769
rect 20720 24803 20772 24812
rect 20720 24769 20729 24803
rect 20729 24769 20763 24803
rect 20763 24769 20772 24803
rect 20720 24760 20772 24769
rect 1676 24599 1728 24608
rect 1676 24565 1685 24599
rect 1685 24565 1719 24599
rect 1719 24565 1728 24599
rect 1676 24556 1728 24565
rect 6000 24556 6052 24608
rect 7840 24556 7892 24608
rect 8944 24556 8996 24608
rect 9128 24599 9180 24608
rect 9128 24565 9137 24599
rect 9137 24565 9171 24599
rect 9171 24565 9180 24599
rect 9128 24556 9180 24565
rect 9864 24599 9916 24608
rect 9864 24565 9873 24599
rect 9873 24565 9907 24599
rect 9907 24565 9916 24599
rect 9864 24556 9916 24565
rect 10416 24599 10468 24608
rect 10416 24565 10425 24599
rect 10425 24565 10459 24599
rect 10459 24565 10468 24599
rect 10416 24556 10468 24565
rect 11244 24556 11296 24608
rect 16580 24692 16632 24744
rect 16856 24692 16908 24744
rect 17868 24692 17920 24744
rect 18788 24692 18840 24744
rect 19984 24692 20036 24744
rect 37556 24760 37608 24812
rect 21088 24692 21140 24744
rect 15016 24624 15068 24676
rect 20812 24624 20864 24676
rect 17684 24556 17736 24608
rect 17776 24556 17828 24608
rect 20076 24599 20128 24608
rect 20076 24565 20085 24599
rect 20085 24565 20119 24599
rect 20119 24565 20128 24599
rect 20076 24556 20128 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2412 24352 2464 24404
rect 4252 24352 4304 24404
rect 4896 24352 4948 24404
rect 2964 24284 3016 24336
rect 7564 24352 7616 24404
rect 7748 24352 7800 24404
rect 9772 24352 9824 24404
rect 9864 24352 9916 24404
rect 11888 24352 11940 24404
rect 12716 24352 12768 24404
rect 16488 24352 16540 24404
rect 18696 24352 18748 24404
rect 35348 24395 35400 24404
rect 35348 24361 35357 24395
rect 35357 24361 35391 24395
rect 35391 24361 35400 24395
rect 35348 24352 35400 24361
rect 8944 24284 8996 24336
rect 4712 24216 4764 24268
rect 5172 24216 5224 24268
rect 5356 24259 5408 24268
rect 5356 24225 5365 24259
rect 5365 24225 5399 24259
rect 5399 24225 5408 24259
rect 5356 24216 5408 24225
rect 5540 24259 5592 24268
rect 5540 24225 5549 24259
rect 5549 24225 5583 24259
rect 5583 24225 5592 24259
rect 5540 24216 5592 24225
rect 6184 24216 6236 24268
rect 10048 24216 10100 24268
rect 1492 24148 1544 24200
rect 2136 24148 2188 24200
rect 2228 24148 2280 24200
rect 4988 24148 5040 24200
rect 5816 24148 5868 24200
rect 6276 24148 6328 24200
rect 9312 24191 9364 24200
rect 5172 24080 5224 24132
rect 6644 24123 6696 24132
rect 6644 24089 6653 24123
rect 6653 24089 6687 24123
rect 6687 24089 6696 24123
rect 7748 24123 7800 24132
rect 6644 24080 6696 24089
rect 7748 24089 7757 24123
rect 7757 24089 7791 24123
rect 7791 24089 7800 24123
rect 7748 24080 7800 24089
rect 7840 24123 7892 24132
rect 7840 24089 7849 24123
rect 7849 24089 7883 24123
rect 7883 24089 7892 24123
rect 7840 24080 7892 24089
rect 8208 24080 8260 24132
rect 9312 24157 9321 24191
rect 9321 24157 9355 24191
rect 9355 24157 9364 24191
rect 9312 24148 9364 24157
rect 12348 24284 12400 24336
rect 14648 24327 14700 24336
rect 14648 24293 14657 24327
rect 14657 24293 14691 24327
rect 14691 24293 14700 24327
rect 14648 24284 14700 24293
rect 11060 24216 11112 24268
rect 11520 24216 11572 24268
rect 25412 24284 25464 24336
rect 17592 24216 17644 24268
rect 17868 24216 17920 24268
rect 20904 24259 20956 24268
rect 8576 24080 8628 24132
rect 11336 24148 11388 24200
rect 14464 24148 14516 24200
rect 16304 24148 16356 24200
rect 16672 24148 16724 24200
rect 17960 24148 18012 24200
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 21088 24259 21140 24268
rect 21088 24225 21097 24259
rect 21097 24225 21131 24259
rect 21131 24225 21140 24259
rect 21088 24216 21140 24225
rect 27252 24148 27304 24200
rect 33140 24148 33192 24200
rect 3332 24055 3384 24064
rect 3332 24021 3341 24055
rect 3341 24021 3375 24055
rect 3375 24021 3384 24055
rect 3332 24012 3384 24021
rect 7380 24012 7432 24064
rect 8852 24012 8904 24064
rect 9404 24055 9456 24064
rect 9404 24021 9413 24055
rect 9413 24021 9447 24055
rect 9447 24021 9456 24055
rect 9404 24012 9456 24021
rect 10140 24055 10192 24064
rect 10140 24021 10149 24055
rect 10149 24021 10183 24055
rect 10183 24021 10192 24055
rect 10140 24012 10192 24021
rect 14188 24080 14240 24132
rect 14832 24080 14884 24132
rect 16580 24080 16632 24132
rect 17408 24080 17460 24132
rect 20076 24080 20128 24132
rect 11980 24012 12032 24064
rect 13452 24012 13504 24064
rect 13636 24055 13688 24064
rect 13636 24021 13645 24055
rect 13645 24021 13679 24055
rect 13679 24021 13688 24055
rect 13636 24012 13688 24021
rect 13912 24012 13964 24064
rect 17776 24012 17828 24064
rect 18972 24012 19024 24064
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1860 23808 1912 23860
rect 3884 23808 3936 23860
rect 4344 23783 4396 23792
rect 4344 23749 4353 23783
rect 4353 23749 4387 23783
rect 4387 23749 4396 23783
rect 4344 23740 4396 23749
rect 5264 23808 5316 23860
rect 2596 23672 2648 23724
rect 2780 23604 2832 23656
rect 2964 23715 3016 23724
rect 2964 23681 2973 23715
rect 2973 23681 3007 23715
rect 3007 23681 3016 23715
rect 2964 23672 3016 23681
rect 3884 23672 3936 23724
rect 4252 23715 4304 23724
rect 4252 23681 4261 23715
rect 4261 23681 4295 23715
rect 4295 23681 4304 23715
rect 4252 23672 4304 23681
rect 4712 23672 4764 23724
rect 4988 23672 5040 23724
rect 7012 23740 7064 23792
rect 7656 23783 7708 23792
rect 7656 23749 7665 23783
rect 7665 23749 7699 23783
rect 7699 23749 7708 23783
rect 7656 23740 7708 23749
rect 8668 23740 8720 23792
rect 4620 23604 4672 23656
rect 8576 23672 8628 23724
rect 9312 23808 9364 23860
rect 11612 23808 11664 23860
rect 13452 23808 13504 23860
rect 9404 23740 9456 23792
rect 13636 23740 13688 23792
rect 9128 23672 9180 23724
rect 11704 23672 11756 23724
rect 13912 23715 13964 23724
rect 5264 23604 5316 23656
rect 6368 23604 6420 23656
rect 8208 23604 8260 23656
rect 3056 23579 3108 23588
rect 3056 23545 3065 23579
rect 3065 23545 3099 23579
rect 3099 23545 3108 23579
rect 3056 23536 3108 23545
rect 5356 23536 5408 23588
rect 5448 23536 5500 23588
rect 11520 23604 11572 23656
rect 11980 23647 12032 23656
rect 11980 23613 11989 23647
rect 11989 23613 12023 23647
rect 12023 23613 12032 23647
rect 11980 23604 12032 23613
rect 13912 23681 13921 23715
rect 13921 23681 13955 23715
rect 13955 23681 13964 23715
rect 13912 23672 13964 23681
rect 14556 23715 14608 23724
rect 14556 23681 14565 23715
rect 14565 23681 14599 23715
rect 14599 23681 14608 23715
rect 14556 23672 14608 23681
rect 14740 23672 14792 23724
rect 13820 23604 13872 23656
rect 14004 23604 14056 23656
rect 14924 23604 14976 23656
rect 17408 23672 17460 23724
rect 20536 23808 20588 23860
rect 18972 23783 19024 23792
rect 18972 23749 18981 23783
rect 18981 23749 19015 23783
rect 19015 23749 19024 23783
rect 18972 23740 19024 23749
rect 19984 23740 20036 23792
rect 20444 23672 20496 23724
rect 34796 23672 34848 23724
rect 38292 23715 38344 23724
rect 38292 23681 38301 23715
rect 38301 23681 38335 23715
rect 38335 23681 38344 23715
rect 38292 23672 38344 23681
rect 9956 23536 10008 23588
rect 10968 23536 11020 23588
rect 14648 23536 14700 23588
rect 2596 23468 2648 23520
rect 4988 23511 5040 23520
rect 4988 23477 4997 23511
rect 4997 23477 5031 23511
rect 5031 23477 5040 23511
rect 4988 23468 5040 23477
rect 8484 23468 8536 23520
rect 8576 23468 8628 23520
rect 8944 23468 8996 23520
rect 9404 23468 9456 23520
rect 11060 23468 11112 23520
rect 13176 23468 13228 23520
rect 13912 23468 13964 23520
rect 14096 23511 14148 23520
rect 14096 23477 14105 23511
rect 14105 23477 14139 23511
rect 14139 23477 14148 23511
rect 14096 23468 14148 23477
rect 15476 23468 15528 23520
rect 19432 23604 19484 23656
rect 18144 23468 18196 23520
rect 18328 23511 18380 23520
rect 18328 23477 18337 23511
rect 18337 23477 18371 23511
rect 18371 23477 18380 23511
rect 18328 23468 18380 23477
rect 21916 23468 21968 23520
rect 34520 23468 34572 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1860 23264 1912 23316
rect 6092 23264 6144 23316
rect 10324 23264 10376 23316
rect 12532 23307 12584 23316
rect 12532 23273 12541 23307
rect 12541 23273 12575 23307
rect 12575 23273 12584 23307
rect 12532 23264 12584 23273
rect 14556 23264 14608 23316
rect 20536 23307 20588 23316
rect 20536 23273 20545 23307
rect 20545 23273 20579 23307
rect 20579 23273 20588 23307
rect 20536 23264 20588 23273
rect 5540 23196 5592 23248
rect 8300 23196 8352 23248
rect 2228 23128 2280 23180
rect 5264 23128 5316 23180
rect 3884 23060 3936 23112
rect 4712 23060 4764 23112
rect 5448 23060 5500 23112
rect 8208 23060 8260 23112
rect 8484 23128 8536 23180
rect 10600 23128 10652 23180
rect 11152 23128 11204 23180
rect 13084 23171 13136 23180
rect 13084 23137 13093 23171
rect 13093 23137 13127 23171
rect 13127 23137 13136 23171
rect 13084 23128 13136 23137
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 14004 23128 14056 23180
rect 14096 23128 14148 23180
rect 2136 22992 2188 23044
rect 4988 22992 5040 23044
rect 5172 22992 5224 23044
rect 3332 22967 3384 22976
rect 3332 22933 3341 22967
rect 3341 22933 3375 22967
rect 3375 22933 3384 22967
rect 3332 22924 3384 22933
rect 4712 22967 4764 22976
rect 4712 22933 4721 22967
rect 4721 22933 4755 22967
rect 4755 22933 4764 22967
rect 4712 22924 4764 22933
rect 6184 22924 6236 22976
rect 8944 22924 8996 22976
rect 13728 23060 13780 23112
rect 15108 23103 15160 23112
rect 9220 23035 9272 23044
rect 9220 23001 9230 23035
rect 9230 23001 9264 23035
rect 9264 23001 9272 23035
rect 9220 22992 9272 23001
rect 9864 23035 9916 23044
rect 9864 23001 9873 23035
rect 9873 23001 9907 23035
rect 9907 23001 9916 23035
rect 9864 22992 9916 23001
rect 13176 23035 13228 23044
rect 13176 23001 13185 23035
rect 13185 23001 13219 23035
rect 13219 23001 13228 23035
rect 13176 22992 13228 23001
rect 14832 22992 14884 23044
rect 14096 22924 14148 22976
rect 14280 22924 14332 22976
rect 15108 23069 15117 23103
rect 15117 23069 15151 23103
rect 15151 23069 15160 23103
rect 15108 23060 15160 23069
rect 17776 23196 17828 23248
rect 15936 23128 15988 23180
rect 18236 23171 18288 23180
rect 18236 23137 18245 23171
rect 18245 23137 18279 23171
rect 18279 23137 18288 23171
rect 18236 23128 18288 23137
rect 18328 23128 18380 23180
rect 33232 23128 33284 23180
rect 17316 23103 17368 23112
rect 17316 23069 17325 23103
rect 17325 23069 17359 23103
rect 17359 23069 17368 23103
rect 17316 23060 17368 23069
rect 19248 23060 19300 23112
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 15660 22924 15712 22976
rect 16764 23035 16816 23044
rect 16764 23001 16773 23035
rect 16773 23001 16807 23035
rect 16807 23001 16816 23035
rect 16764 22992 16816 23001
rect 17408 22967 17460 22976
rect 17408 22933 17417 22967
rect 17417 22933 17451 22967
rect 17451 22933 17460 22967
rect 17408 22924 17460 22933
rect 18880 22967 18932 22976
rect 18880 22933 18889 22967
rect 18889 22933 18923 22967
rect 18923 22933 18932 22967
rect 18880 22924 18932 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1860 22720 1912 22772
rect 2136 22720 2188 22772
rect 3424 22720 3476 22772
rect 3792 22652 3844 22704
rect 5264 22695 5316 22704
rect 5264 22661 5273 22695
rect 5273 22661 5307 22695
rect 5307 22661 5316 22695
rect 5264 22652 5316 22661
rect 1584 22627 1636 22636
rect 1584 22593 1593 22627
rect 1593 22593 1627 22627
rect 1627 22593 1636 22627
rect 1584 22584 1636 22593
rect 2228 22627 2280 22636
rect 2228 22593 2237 22627
rect 2237 22593 2271 22627
rect 2271 22593 2280 22627
rect 2228 22584 2280 22593
rect 4620 22627 4672 22636
rect 4620 22593 4629 22627
rect 4629 22593 4663 22627
rect 4663 22593 4672 22627
rect 4620 22584 4672 22593
rect 4988 22584 5040 22636
rect 7932 22720 7984 22772
rect 8208 22720 8260 22772
rect 9128 22720 9180 22772
rect 6184 22652 6236 22704
rect 6736 22695 6788 22704
rect 6736 22661 6745 22695
rect 6745 22661 6779 22695
rect 6779 22661 6788 22695
rect 6736 22652 6788 22661
rect 6920 22652 6972 22704
rect 8944 22652 8996 22704
rect 9588 22720 9640 22772
rect 12992 22720 13044 22772
rect 2320 22380 2372 22432
rect 2596 22380 2648 22432
rect 5172 22516 5224 22568
rect 3608 22448 3660 22500
rect 8116 22584 8168 22636
rect 9588 22584 9640 22636
rect 9956 22584 10008 22636
rect 10140 22584 10192 22636
rect 11060 22652 11112 22704
rect 11428 22652 11480 22704
rect 13820 22695 13872 22704
rect 13820 22661 13829 22695
rect 13829 22661 13863 22695
rect 13863 22661 13872 22695
rect 13820 22652 13872 22661
rect 14924 22720 14976 22772
rect 19248 22763 19300 22772
rect 15292 22652 15344 22704
rect 15476 22695 15528 22704
rect 15476 22661 15485 22695
rect 15485 22661 15519 22695
rect 15519 22661 15528 22695
rect 15476 22652 15528 22661
rect 19248 22729 19257 22763
rect 19257 22729 19291 22763
rect 19291 22729 19300 22763
rect 19248 22720 19300 22729
rect 17408 22695 17460 22704
rect 17408 22661 17417 22695
rect 17417 22661 17451 22695
rect 17451 22661 17460 22695
rect 17408 22652 17460 22661
rect 17868 22652 17920 22704
rect 12716 22584 12768 22636
rect 13084 22584 13136 22636
rect 17960 22584 18012 22636
rect 18420 22584 18472 22636
rect 20720 22652 20772 22704
rect 19248 22584 19300 22636
rect 21180 22584 21232 22636
rect 21456 22627 21508 22636
rect 21456 22593 21465 22627
rect 21465 22593 21499 22627
rect 21499 22593 21508 22627
rect 21456 22584 21508 22593
rect 7104 22448 7156 22500
rect 5816 22380 5868 22432
rect 7656 22380 7708 22432
rect 9772 22516 9824 22568
rect 10968 22516 11020 22568
rect 11888 22559 11940 22568
rect 11888 22525 11897 22559
rect 11897 22525 11931 22559
rect 11931 22525 11940 22559
rect 11888 22516 11940 22525
rect 13728 22559 13780 22568
rect 13728 22525 13737 22559
rect 13737 22525 13771 22559
rect 13771 22525 13780 22559
rect 13728 22516 13780 22525
rect 16764 22516 16816 22568
rect 10784 22448 10836 22500
rect 11980 22448 12032 22500
rect 17040 22448 17092 22500
rect 17408 22516 17460 22568
rect 18052 22559 18104 22568
rect 18052 22525 18061 22559
rect 18061 22525 18095 22559
rect 18095 22525 18104 22559
rect 18052 22516 18104 22525
rect 18604 22516 18656 22568
rect 20812 22559 20864 22568
rect 20812 22525 20821 22559
rect 20821 22525 20855 22559
rect 20855 22525 20864 22559
rect 20812 22516 20864 22525
rect 30472 22516 30524 22568
rect 9772 22380 9824 22432
rect 9864 22380 9916 22432
rect 12992 22380 13044 22432
rect 15200 22380 15252 22432
rect 15292 22380 15344 22432
rect 18788 22380 18840 22432
rect 20444 22423 20496 22432
rect 20444 22389 20453 22423
rect 20453 22389 20487 22423
rect 20487 22389 20496 22423
rect 20444 22380 20496 22389
rect 33324 22380 33376 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2964 22176 3016 22228
rect 4068 22176 4120 22228
rect 5264 22176 5316 22228
rect 5448 22176 5500 22228
rect 9036 22176 9088 22228
rect 9220 22176 9272 22228
rect 12532 22176 12584 22228
rect 13452 22176 13504 22228
rect 18880 22176 18932 22228
rect 7288 22108 7340 22160
rect 9312 22108 9364 22160
rect 13544 22108 13596 22160
rect 2136 22040 2188 22092
rect 4528 22040 4580 22092
rect 5540 22040 5592 22092
rect 3884 21972 3936 22024
rect 8944 22040 8996 22092
rect 9588 22040 9640 22092
rect 11244 22040 11296 22092
rect 11704 22040 11756 22092
rect 11888 22040 11940 22092
rect 13636 22040 13688 22092
rect 14372 22083 14424 22092
rect 14372 22049 14381 22083
rect 14381 22049 14415 22083
rect 14415 22049 14424 22083
rect 14372 22040 14424 22049
rect 14648 22083 14700 22092
rect 14648 22049 14657 22083
rect 14657 22049 14691 22083
rect 14691 22049 14700 22083
rect 14648 22040 14700 22049
rect 16120 22083 16172 22092
rect 16120 22049 16129 22083
rect 16129 22049 16163 22083
rect 16163 22049 16172 22083
rect 16120 22040 16172 22049
rect 18420 22040 18472 22092
rect 18696 22040 18748 22092
rect 18880 22083 18932 22092
rect 18880 22049 18889 22083
rect 18889 22049 18923 22083
rect 18923 22049 18932 22083
rect 18880 22040 18932 22049
rect 21916 22083 21968 22092
rect 21916 22049 21925 22083
rect 21925 22049 21959 22083
rect 21959 22049 21968 22083
rect 21916 22040 21968 22049
rect 2596 21904 2648 21956
rect 1400 21836 1452 21888
rect 1860 21836 1912 21888
rect 10416 21972 10468 22024
rect 4252 21904 4304 21956
rect 4804 21904 4856 21956
rect 5356 21904 5408 21956
rect 9128 21947 9180 21956
rect 9128 21913 9137 21947
rect 9137 21913 9171 21947
rect 9171 21913 9180 21947
rect 9128 21904 9180 21913
rect 5816 21836 5868 21888
rect 6276 21836 6328 21888
rect 6644 21836 6696 21888
rect 6828 21836 6880 21888
rect 12348 21972 12400 22024
rect 15108 21972 15160 22024
rect 17500 22015 17552 22024
rect 12072 21947 12124 21956
rect 12072 21913 12081 21947
rect 12081 21913 12115 21947
rect 12115 21913 12124 21947
rect 12072 21904 12124 21913
rect 12256 21904 12308 21956
rect 13820 21904 13872 21956
rect 14188 21904 14240 21956
rect 14556 21904 14608 21956
rect 17500 21981 17509 22015
rect 17509 21981 17543 22015
rect 17543 21981 17552 22015
rect 17500 21972 17552 21981
rect 19340 21972 19392 22024
rect 20168 21972 20220 22024
rect 38292 22015 38344 22024
rect 38292 21981 38301 22015
rect 38301 21981 38335 22015
rect 38335 21981 38344 22015
rect 38292 21972 38344 21981
rect 18052 21904 18104 21956
rect 18328 21947 18380 21956
rect 18328 21913 18330 21947
rect 18330 21913 18364 21947
rect 18364 21913 18380 21947
rect 18328 21904 18380 21913
rect 18696 21904 18748 21956
rect 21272 21947 21324 21956
rect 21272 21913 21281 21947
rect 21281 21913 21315 21947
rect 21315 21913 21324 21947
rect 21272 21904 21324 21913
rect 21824 21947 21876 21956
rect 21824 21913 21833 21947
rect 21833 21913 21867 21947
rect 21867 21913 21876 21947
rect 21824 21904 21876 21913
rect 13544 21836 13596 21888
rect 17960 21836 18012 21888
rect 18972 21836 19024 21888
rect 19984 21836 20036 21888
rect 32220 21836 32272 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4252 21675 4304 21684
rect 4252 21641 4261 21675
rect 4261 21641 4295 21675
rect 4295 21641 4304 21675
rect 4252 21632 4304 21641
rect 2044 21564 2096 21616
rect 3240 21564 3292 21616
rect 6460 21564 6512 21616
rect 3700 21496 3752 21548
rect 6184 21496 6236 21548
rect 2136 21428 2188 21480
rect 8300 21632 8352 21684
rect 8484 21632 8536 21684
rect 7472 21564 7524 21616
rect 12256 21632 12308 21684
rect 16856 21632 16908 21684
rect 17500 21632 17552 21684
rect 20168 21675 20220 21684
rect 20168 21641 20177 21675
rect 20177 21641 20211 21675
rect 20211 21641 20220 21675
rect 20168 21632 20220 21641
rect 21824 21632 21876 21684
rect 33140 21632 33192 21684
rect 10140 21607 10192 21616
rect 10140 21573 10149 21607
rect 10149 21573 10183 21607
rect 10183 21573 10192 21607
rect 10140 21564 10192 21573
rect 14464 21564 14516 21616
rect 16948 21564 17000 21616
rect 8484 21428 8536 21480
rect 8852 21428 8904 21480
rect 9220 21471 9272 21480
rect 9220 21437 9229 21471
rect 9229 21437 9263 21471
rect 9263 21437 9272 21471
rect 9220 21428 9272 21437
rect 2228 21360 2280 21412
rect 4620 21360 4672 21412
rect 7104 21292 7156 21344
rect 8484 21292 8536 21344
rect 9128 21292 9180 21344
rect 10324 21496 10376 21548
rect 12808 21496 12860 21548
rect 13360 21539 13412 21548
rect 13360 21505 13369 21539
rect 13369 21505 13403 21539
rect 13403 21505 13412 21539
rect 13360 21496 13412 21505
rect 14004 21539 14056 21548
rect 14004 21505 14013 21539
rect 14013 21505 14047 21539
rect 14047 21505 14056 21539
rect 14004 21496 14056 21505
rect 15844 21539 15896 21548
rect 15844 21505 15853 21539
rect 15853 21505 15887 21539
rect 15887 21505 15896 21539
rect 15844 21496 15896 21505
rect 16856 21539 16908 21548
rect 16856 21505 16865 21539
rect 16865 21505 16899 21539
rect 16899 21505 16908 21539
rect 16856 21496 16908 21505
rect 17132 21564 17184 21616
rect 18972 21607 19024 21616
rect 18972 21573 18981 21607
rect 18981 21573 19015 21607
rect 19015 21573 19024 21607
rect 18972 21564 19024 21573
rect 18144 21496 18196 21548
rect 21180 21539 21232 21548
rect 9588 21360 9640 21412
rect 11888 21360 11940 21412
rect 13268 21428 13320 21480
rect 15660 21471 15712 21480
rect 14556 21360 14608 21412
rect 14924 21292 14976 21344
rect 15660 21437 15669 21471
rect 15669 21437 15703 21471
rect 15703 21437 15712 21471
rect 15660 21428 15712 21437
rect 18420 21428 18472 21480
rect 19340 21428 19392 21480
rect 21180 21505 21189 21539
rect 21189 21505 21223 21539
rect 21223 21505 21232 21539
rect 21180 21496 21232 21505
rect 21364 21496 21416 21548
rect 21548 21496 21600 21548
rect 25320 21496 25372 21548
rect 34520 21496 34572 21548
rect 21916 21428 21968 21480
rect 20076 21360 20128 21412
rect 35624 21360 35676 21412
rect 16856 21292 16908 21344
rect 23664 21292 23716 21344
rect 29000 21292 29052 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2044 21088 2096 21140
rect 2228 21088 2280 21140
rect 5356 21088 5408 21140
rect 1400 21020 1452 21072
rect 4160 21020 4212 21072
rect 4712 21020 4764 21072
rect 4896 21020 4948 21072
rect 11612 20952 11664 21004
rect 12164 20952 12216 21004
rect 17132 21088 17184 21140
rect 13912 21020 13964 21072
rect 16580 21020 16632 21072
rect 19064 21020 19116 21072
rect 20076 21063 20128 21072
rect 15660 20952 15712 21004
rect 16488 20952 16540 21004
rect 16856 20995 16908 21004
rect 16856 20961 16865 20995
rect 16865 20961 16899 20995
rect 16899 20961 16908 20995
rect 16856 20952 16908 20961
rect 19340 20952 19392 21004
rect 20076 21029 20085 21063
rect 20085 21029 20119 21063
rect 20119 21029 20128 21063
rect 20076 21020 20128 21029
rect 21272 21020 21324 21072
rect 23388 21020 23440 21072
rect 21916 20995 21968 21004
rect 21916 20961 21925 20995
rect 21925 20961 21959 20995
rect 21959 20961 21968 20995
rect 21916 20952 21968 20961
rect 22468 20952 22520 21004
rect 4896 20884 4948 20936
rect 5172 20884 5224 20936
rect 5356 20884 5408 20936
rect 7472 20884 7524 20936
rect 5908 20816 5960 20868
rect 8208 20816 8260 20868
rect 6828 20748 6880 20800
rect 7288 20748 7340 20800
rect 7748 20748 7800 20800
rect 8852 20884 8904 20936
rect 9128 20927 9180 20936
rect 9128 20893 9137 20927
rect 9137 20893 9171 20927
rect 9171 20893 9180 20927
rect 9128 20884 9180 20893
rect 11060 20884 11112 20936
rect 13544 20927 13596 20936
rect 13544 20893 13553 20927
rect 13553 20893 13587 20927
rect 13587 20893 13596 20927
rect 13544 20884 13596 20893
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 14372 20884 14424 20936
rect 8484 20816 8536 20868
rect 9864 20816 9916 20868
rect 8852 20748 8904 20800
rect 9496 20748 9548 20800
rect 9680 20748 9732 20800
rect 13912 20816 13964 20868
rect 14004 20816 14056 20868
rect 15108 20816 15160 20868
rect 15660 20816 15712 20868
rect 12348 20748 12400 20800
rect 15016 20748 15068 20800
rect 15476 20748 15528 20800
rect 15936 20748 15988 20800
rect 18788 20816 18840 20868
rect 21180 20884 21232 20936
rect 32220 20927 32272 20936
rect 32220 20893 32229 20927
rect 32229 20893 32263 20927
rect 32263 20893 32272 20927
rect 32220 20884 32272 20893
rect 19984 20816 20036 20868
rect 22836 20859 22888 20868
rect 20076 20748 20128 20800
rect 22836 20825 22845 20859
rect 22845 20825 22879 20859
rect 22879 20825 22888 20859
rect 22836 20816 22888 20825
rect 23572 20748 23624 20800
rect 32128 20791 32180 20800
rect 32128 20757 32137 20791
rect 32137 20757 32171 20791
rect 32171 20757 32180 20791
rect 32128 20748 32180 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 3976 20544 4028 20596
rect 6920 20544 6972 20596
rect 10232 20587 10284 20596
rect 3148 20476 3200 20528
rect 4160 20519 4212 20528
rect 4160 20485 4169 20519
rect 4169 20485 4203 20519
rect 4203 20485 4212 20519
rect 4160 20476 4212 20485
rect 2872 20408 2924 20460
rect 3424 20340 3476 20392
rect 4620 20340 4672 20392
rect 5540 20476 5592 20528
rect 7840 20476 7892 20528
rect 8760 20476 8812 20528
rect 5172 20451 5224 20460
rect 5172 20417 5181 20451
rect 5181 20417 5215 20451
rect 5215 20417 5224 20451
rect 5172 20408 5224 20417
rect 6276 20408 6328 20460
rect 7104 20408 7156 20460
rect 9036 20408 9088 20460
rect 9864 20408 9916 20460
rect 10232 20553 10241 20587
rect 10241 20553 10275 20587
rect 10275 20553 10284 20587
rect 10232 20544 10284 20553
rect 12348 20587 12400 20596
rect 12348 20553 12357 20587
rect 12357 20553 12391 20587
rect 12391 20553 12400 20587
rect 12348 20544 12400 20553
rect 14188 20544 14240 20596
rect 14832 20587 14884 20596
rect 14832 20553 14841 20587
rect 14841 20553 14875 20587
rect 14875 20553 14884 20587
rect 14832 20544 14884 20553
rect 16028 20544 16080 20596
rect 18512 20544 18564 20596
rect 19340 20544 19392 20596
rect 20076 20544 20128 20596
rect 21180 20544 21232 20596
rect 22836 20587 22888 20596
rect 22836 20553 22845 20587
rect 22845 20553 22879 20587
rect 22879 20553 22888 20587
rect 22836 20544 22888 20553
rect 23572 20544 23624 20596
rect 14280 20476 14332 20528
rect 11612 20408 11664 20460
rect 12716 20408 12768 20460
rect 14004 20451 14056 20460
rect 14004 20417 14013 20451
rect 14013 20417 14047 20451
rect 14047 20417 14056 20451
rect 14004 20408 14056 20417
rect 6368 20340 6420 20392
rect 7472 20383 7524 20392
rect 7472 20349 7481 20383
rect 7481 20349 7515 20383
rect 7515 20349 7524 20383
rect 7472 20340 7524 20349
rect 3424 20204 3476 20256
rect 7288 20272 7340 20324
rect 7840 20340 7892 20392
rect 9496 20383 9548 20392
rect 9496 20349 9505 20383
rect 9505 20349 9539 20383
rect 9539 20349 9548 20383
rect 9496 20340 9548 20349
rect 11060 20340 11112 20392
rect 11336 20340 11388 20392
rect 14924 20408 14976 20460
rect 15384 20408 15436 20460
rect 17316 20451 17368 20460
rect 17316 20417 17325 20451
rect 17325 20417 17359 20451
rect 17359 20417 17368 20451
rect 17316 20408 17368 20417
rect 17684 20408 17736 20460
rect 18144 20408 18196 20460
rect 18696 20408 18748 20460
rect 18052 20340 18104 20392
rect 21364 20408 21416 20460
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 23664 20451 23716 20460
rect 23664 20417 23673 20451
rect 23673 20417 23707 20451
rect 23707 20417 23716 20451
rect 23664 20408 23716 20417
rect 21088 20340 21140 20392
rect 24584 20340 24636 20392
rect 5540 20204 5592 20256
rect 7380 20204 7432 20256
rect 7472 20204 7524 20256
rect 9128 20204 9180 20256
rect 9588 20204 9640 20256
rect 13268 20204 13320 20256
rect 13544 20247 13596 20256
rect 13544 20213 13553 20247
rect 13553 20213 13587 20247
rect 13587 20213 13596 20247
rect 13544 20204 13596 20213
rect 13728 20204 13780 20256
rect 15476 20204 15528 20256
rect 22284 20204 22336 20256
rect 25504 20204 25556 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3424 20043 3476 20052
rect 3424 20009 3433 20043
rect 3433 20009 3467 20043
rect 3467 20009 3476 20043
rect 3424 20000 3476 20009
rect 5172 20000 5224 20052
rect 2044 19864 2096 19916
rect 4160 19796 4212 19848
rect 4896 19932 4948 19984
rect 6184 20000 6236 20052
rect 6276 20000 6328 20052
rect 6920 20000 6972 20052
rect 9036 20000 9088 20052
rect 9220 20000 9272 20052
rect 6276 19864 6328 19916
rect 6368 19864 6420 19916
rect 7380 19932 7432 19984
rect 12072 20000 12124 20052
rect 16028 20000 16080 20052
rect 16948 20000 17000 20052
rect 18236 20000 18288 20052
rect 14372 19932 14424 19984
rect 16488 19932 16540 19984
rect 7012 19864 7064 19916
rect 8852 19864 8904 19916
rect 9036 19864 9088 19916
rect 9128 19864 9180 19916
rect 11796 19864 11848 19916
rect 12992 19864 13044 19916
rect 29184 20000 29236 20052
rect 20168 19932 20220 19984
rect 2688 19728 2740 19780
rect 4620 19728 4672 19780
rect 8208 19796 8260 19848
rect 5724 19728 5776 19780
rect 8760 19728 8812 19780
rect 10324 19728 10376 19780
rect 10876 19728 10928 19780
rect 14280 19796 14332 19848
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 17684 19796 17736 19848
rect 21364 19864 21416 19916
rect 20168 19796 20220 19848
rect 20996 19839 21048 19848
rect 20996 19805 21005 19839
rect 21005 19805 21039 19839
rect 21039 19805 21048 19839
rect 20996 19796 21048 19805
rect 15752 19771 15804 19780
rect 3424 19660 3476 19712
rect 3976 19660 4028 19712
rect 4804 19660 4856 19712
rect 5908 19660 5960 19712
rect 7104 19660 7156 19712
rect 8392 19660 8444 19712
rect 15752 19737 15761 19771
rect 15761 19737 15795 19771
rect 15795 19737 15804 19771
rect 15752 19728 15804 19737
rect 15844 19771 15896 19780
rect 15844 19737 15853 19771
rect 15853 19737 15887 19771
rect 15887 19737 15896 19771
rect 16396 19771 16448 19780
rect 15844 19728 15896 19737
rect 16396 19737 16405 19771
rect 16405 19737 16439 19771
rect 16439 19737 16448 19771
rect 16396 19728 16448 19737
rect 17040 19771 17092 19780
rect 17040 19737 17049 19771
rect 17049 19737 17083 19771
rect 17083 19737 17092 19771
rect 17040 19728 17092 19737
rect 17224 19728 17276 19780
rect 29736 19932 29788 19984
rect 24032 19907 24084 19916
rect 24032 19873 24041 19907
rect 24041 19873 24075 19907
rect 24075 19873 24084 19907
rect 24032 19864 24084 19873
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 25412 19839 25464 19848
rect 25412 19805 25421 19839
rect 25421 19805 25455 19839
rect 25455 19805 25464 19839
rect 25412 19796 25464 19805
rect 38292 19839 38344 19848
rect 38292 19805 38301 19839
rect 38301 19805 38335 19839
rect 38335 19805 38344 19839
rect 38292 19796 38344 19805
rect 23112 19728 23164 19780
rect 20076 19660 20128 19712
rect 20260 19703 20312 19712
rect 20260 19669 20269 19703
rect 20269 19669 20303 19703
rect 20303 19669 20312 19703
rect 20260 19660 20312 19669
rect 20812 19703 20864 19712
rect 20812 19669 20821 19703
rect 20821 19669 20855 19703
rect 20855 19669 20864 19703
rect 20812 19660 20864 19669
rect 22100 19703 22152 19712
rect 22100 19669 22109 19703
rect 22109 19669 22143 19703
rect 22143 19669 22152 19703
rect 25228 19703 25280 19712
rect 22100 19660 22152 19669
rect 25228 19669 25237 19703
rect 25237 19669 25271 19703
rect 25271 19669 25280 19703
rect 25228 19660 25280 19669
rect 35532 19660 35584 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 2228 19456 2280 19508
rect 8116 19456 8168 19508
rect 8392 19456 8444 19508
rect 3884 19388 3936 19440
rect 4068 19388 4120 19440
rect 5908 19388 5960 19440
rect 9680 19388 9732 19440
rect 9956 19499 10008 19508
rect 9956 19465 9965 19499
rect 9965 19465 9999 19499
rect 9999 19465 10008 19499
rect 9956 19456 10008 19465
rect 13728 19456 13780 19508
rect 14280 19499 14332 19508
rect 14280 19465 14289 19499
rect 14289 19465 14323 19499
rect 14323 19465 14332 19499
rect 14280 19456 14332 19465
rect 14372 19456 14424 19508
rect 15844 19456 15896 19508
rect 2320 19363 2372 19372
rect 2320 19329 2329 19363
rect 2329 19329 2363 19363
rect 2363 19329 2372 19363
rect 2320 19320 2372 19329
rect 3332 19320 3384 19372
rect 3700 19320 3752 19372
rect 7288 19320 7340 19372
rect 3976 19252 4028 19304
rect 5724 19252 5776 19304
rect 9588 19320 9640 19372
rect 9680 19252 9732 19304
rect 9864 19363 9916 19372
rect 9864 19329 9873 19363
rect 9873 19329 9907 19363
rect 9907 19329 9916 19363
rect 9864 19320 9916 19329
rect 10324 19320 10376 19372
rect 10968 19320 11020 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 13544 19388 13596 19440
rect 18420 19456 18472 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 21180 19456 21232 19508
rect 16120 19431 16172 19440
rect 14372 19320 14424 19372
rect 14464 19363 14516 19372
rect 14464 19329 14473 19363
rect 14473 19329 14507 19363
rect 14507 19329 14516 19363
rect 14464 19320 14516 19329
rect 14648 19320 14700 19372
rect 12072 19295 12124 19304
rect 10600 19184 10652 19236
rect 7104 19159 7156 19168
rect 7104 19125 7113 19159
rect 7113 19125 7147 19159
rect 7147 19125 7156 19159
rect 7104 19116 7156 19125
rect 7196 19116 7248 19168
rect 7656 19159 7708 19168
rect 7656 19125 7665 19159
rect 7665 19125 7699 19159
rect 7699 19125 7708 19159
rect 7656 19116 7708 19125
rect 9588 19116 9640 19168
rect 12072 19261 12081 19295
rect 12081 19261 12115 19295
rect 12115 19261 12124 19295
rect 12072 19252 12124 19261
rect 13268 19252 13320 19304
rect 13636 19295 13688 19304
rect 13636 19261 13645 19295
rect 13645 19261 13679 19295
rect 13679 19261 13688 19295
rect 13636 19252 13688 19261
rect 16120 19397 16129 19431
rect 16129 19397 16163 19431
rect 16163 19397 16172 19431
rect 16120 19388 16172 19397
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 17776 19295 17828 19304
rect 17776 19261 17785 19295
rect 17785 19261 17819 19295
rect 17819 19261 17828 19295
rect 17776 19252 17828 19261
rect 19432 19320 19484 19372
rect 20260 19320 20312 19372
rect 20352 19363 20404 19372
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 20352 19320 20404 19329
rect 21180 19320 21232 19372
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 23112 19363 23164 19372
rect 23112 19329 23121 19363
rect 23121 19329 23155 19363
rect 23155 19329 23164 19363
rect 23112 19320 23164 19329
rect 32128 19388 32180 19440
rect 25504 19363 25556 19372
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 18788 19252 18840 19304
rect 15660 19184 15712 19236
rect 22100 19184 22152 19236
rect 24768 19252 24820 19304
rect 25504 19329 25513 19363
rect 25513 19329 25547 19363
rect 25547 19329 25556 19363
rect 25504 19320 25556 19329
rect 25044 19252 25096 19304
rect 25872 19252 25924 19304
rect 25228 19184 25280 19236
rect 11060 19159 11112 19168
rect 11060 19125 11069 19159
rect 11069 19125 11103 19159
rect 11103 19125 11112 19159
rect 11060 19116 11112 19125
rect 12440 19116 12492 19168
rect 21272 19116 21324 19168
rect 24676 19116 24728 19168
rect 24860 19116 24912 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 6092 18844 6144 18896
rect 6368 18844 6420 18896
rect 1952 18776 2004 18828
rect 4620 18776 4672 18828
rect 4804 18819 4856 18828
rect 4804 18785 4813 18819
rect 4813 18785 4847 18819
rect 4847 18785 4856 18819
rect 4804 18776 4856 18785
rect 5724 18776 5776 18828
rect 8116 18819 8168 18828
rect 8116 18785 8125 18819
rect 8125 18785 8159 18819
rect 8159 18785 8168 18819
rect 8116 18776 8168 18785
rect 12440 18912 12492 18964
rect 12992 18955 13044 18964
rect 12992 18921 13001 18955
rect 13001 18921 13035 18955
rect 13035 18921 13044 18955
rect 12992 18912 13044 18921
rect 13084 18912 13136 18964
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 20996 18912 21048 18964
rect 21456 18912 21508 18964
rect 25412 18912 25464 18964
rect 25872 18912 25924 18964
rect 8668 18844 8720 18896
rect 18328 18844 18380 18896
rect 21548 18844 21600 18896
rect 24768 18844 24820 18896
rect 9220 18776 9272 18828
rect 4436 18708 4488 18760
rect 6920 18708 6972 18760
rect 7840 18708 7892 18760
rect 11060 18776 11112 18828
rect 11152 18776 11204 18828
rect 9496 18708 9548 18760
rect 10876 18751 10928 18760
rect 10876 18717 10885 18751
rect 10885 18717 10919 18751
rect 10919 18717 10928 18751
rect 10876 18708 10928 18717
rect 11796 18751 11848 18760
rect 3056 18640 3108 18692
rect 5172 18640 5224 18692
rect 5632 18640 5684 18692
rect 10600 18683 10652 18692
rect 8944 18572 8996 18624
rect 10600 18649 10609 18683
rect 10609 18649 10643 18683
rect 10643 18649 10652 18683
rect 10600 18640 10652 18649
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 13268 18776 13320 18828
rect 15568 18819 15620 18828
rect 15568 18785 15577 18819
rect 15577 18785 15611 18819
rect 15611 18785 15620 18819
rect 15568 18776 15620 18785
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 19432 18776 19484 18828
rect 24032 18819 24084 18828
rect 24032 18785 24041 18819
rect 24041 18785 24075 18819
rect 24075 18785 24084 18819
rect 24032 18776 24084 18785
rect 24676 18819 24728 18828
rect 24676 18785 24685 18819
rect 24685 18785 24719 18819
rect 24719 18785 24728 18819
rect 24676 18776 24728 18785
rect 25320 18819 25372 18828
rect 25320 18785 25329 18819
rect 25329 18785 25363 18819
rect 25363 18785 25372 18819
rect 25320 18776 25372 18785
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 14832 18751 14884 18760
rect 14832 18717 14841 18751
rect 14841 18717 14875 18751
rect 14875 18717 14884 18751
rect 14832 18708 14884 18717
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 19984 18708 20036 18760
rect 20904 18708 20956 18760
rect 20996 18708 21048 18760
rect 26608 18751 26660 18760
rect 13820 18640 13872 18692
rect 16580 18683 16632 18692
rect 10692 18572 10744 18624
rect 10784 18572 10836 18624
rect 12348 18572 12400 18624
rect 16580 18649 16589 18683
rect 16589 18649 16623 18683
rect 16623 18649 16632 18683
rect 16580 18640 16632 18649
rect 16672 18683 16724 18692
rect 16672 18649 16681 18683
rect 16681 18649 16715 18683
rect 16715 18649 16724 18683
rect 23388 18683 23440 18692
rect 16672 18640 16724 18649
rect 23388 18649 23397 18683
rect 23397 18649 23431 18683
rect 23431 18649 23440 18683
rect 23388 18640 23440 18649
rect 24768 18683 24820 18692
rect 20720 18572 20772 18624
rect 22652 18615 22704 18624
rect 22652 18581 22661 18615
rect 22661 18581 22695 18615
rect 22695 18581 22704 18615
rect 22652 18572 22704 18581
rect 24768 18649 24777 18683
rect 24777 18649 24811 18683
rect 24811 18649 24820 18683
rect 24768 18640 24820 18649
rect 25136 18640 25188 18692
rect 26608 18717 26617 18751
rect 26617 18717 26651 18751
rect 26651 18717 26660 18751
rect 26608 18708 26660 18717
rect 38292 18751 38344 18760
rect 24860 18572 24912 18624
rect 38292 18717 38301 18751
rect 38301 18717 38335 18751
rect 38335 18717 38344 18751
rect 38292 18708 38344 18717
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 3240 18368 3292 18420
rect 4436 18368 4488 18420
rect 7196 18368 7248 18420
rect 8300 18368 8352 18420
rect 8760 18368 8812 18420
rect 10232 18368 10284 18420
rect 3516 18300 3568 18352
rect 4712 18300 4764 18352
rect 5356 18300 5408 18352
rect 8208 18300 8260 18352
rect 5724 18275 5776 18284
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 8944 18300 8996 18352
rect 10048 18300 10100 18352
rect 10692 18300 10744 18352
rect 5724 18232 5776 18241
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 2044 18164 2096 18216
rect 3424 18071 3476 18080
rect 3424 18037 3433 18071
rect 3433 18037 3467 18071
rect 3467 18037 3476 18071
rect 3424 18028 3476 18037
rect 3792 18028 3844 18080
rect 4160 18028 4212 18080
rect 6092 18164 6144 18216
rect 6644 18207 6696 18216
rect 6644 18173 6653 18207
rect 6653 18173 6687 18207
rect 6687 18173 6696 18207
rect 6644 18164 6696 18173
rect 7472 18164 7524 18216
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 10876 18232 10928 18284
rect 12624 18300 12676 18352
rect 13452 18343 13504 18352
rect 13452 18309 13461 18343
rect 13461 18309 13495 18343
rect 13495 18309 13504 18343
rect 15752 18368 15804 18420
rect 16580 18368 16632 18420
rect 19340 18368 19392 18420
rect 19984 18368 20036 18420
rect 13452 18300 13504 18309
rect 17316 18300 17368 18352
rect 17592 18300 17644 18352
rect 22376 18368 22428 18420
rect 23388 18368 23440 18420
rect 24676 18368 24728 18420
rect 24768 18368 24820 18420
rect 9680 18164 9732 18216
rect 9956 18164 10008 18216
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 11060 18164 11112 18216
rect 12808 18096 12860 18148
rect 16764 18232 16816 18284
rect 17868 18232 17920 18284
rect 20812 18232 20864 18284
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 22652 18232 22704 18284
rect 29000 18300 29052 18352
rect 24952 18275 25004 18284
rect 24952 18241 24961 18275
rect 24961 18241 24995 18275
rect 24995 18241 25004 18275
rect 24952 18232 25004 18241
rect 25596 18275 25648 18284
rect 25596 18241 25605 18275
rect 25605 18241 25639 18275
rect 25639 18241 25648 18275
rect 25596 18232 25648 18241
rect 26240 18275 26292 18284
rect 26240 18241 26249 18275
rect 26249 18241 26283 18275
rect 26283 18241 26292 18275
rect 26240 18232 26292 18241
rect 35532 18232 35584 18284
rect 15292 18164 15344 18216
rect 15752 18164 15804 18216
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 17040 18207 17092 18216
rect 17040 18173 17049 18207
rect 17049 18173 17083 18207
rect 17083 18173 17092 18207
rect 17040 18164 17092 18173
rect 18512 18207 18564 18216
rect 18512 18173 18521 18207
rect 18521 18173 18555 18207
rect 18555 18173 18564 18207
rect 18512 18164 18564 18173
rect 18880 18164 18932 18216
rect 18144 18096 18196 18148
rect 21364 18164 21416 18216
rect 22284 18164 22336 18216
rect 25044 18096 25096 18148
rect 16488 18028 16540 18080
rect 20720 18028 20772 18080
rect 24768 18071 24820 18080
rect 24768 18037 24777 18071
rect 24777 18037 24811 18071
rect 24811 18037 24820 18071
rect 24768 18028 24820 18037
rect 34244 18071 34296 18080
rect 34244 18037 34253 18071
rect 34253 18037 34287 18071
rect 34287 18037 34296 18071
rect 34244 18028 34296 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 8576 17867 8628 17876
rect 5356 17756 5408 17808
rect 4804 17688 4856 17740
rect 7380 17688 7432 17740
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 8668 17824 8720 17876
rect 7840 17756 7892 17808
rect 8760 17756 8812 17808
rect 11428 17731 11480 17740
rect 11428 17697 11437 17731
rect 11437 17697 11471 17731
rect 11471 17697 11480 17731
rect 11428 17688 11480 17697
rect 11704 17756 11756 17808
rect 12624 17688 12676 17740
rect 15016 17688 15068 17740
rect 17776 17824 17828 17876
rect 22376 17824 22428 17876
rect 23112 17867 23164 17876
rect 23112 17833 23121 17867
rect 23121 17833 23155 17867
rect 23155 17833 23164 17867
rect 23112 17824 23164 17833
rect 24952 17824 25004 17876
rect 26608 17824 26660 17876
rect 18512 17756 18564 17808
rect 3424 17620 3476 17672
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 1768 17552 1820 17604
rect 3700 17552 3752 17604
rect 3424 17484 3476 17536
rect 3792 17484 3844 17536
rect 4620 17595 4672 17604
rect 4620 17561 4629 17595
rect 4629 17561 4663 17595
rect 4663 17561 4672 17595
rect 4620 17552 4672 17561
rect 5080 17552 5132 17604
rect 6368 17595 6420 17604
rect 6368 17561 6377 17595
rect 6377 17561 6411 17595
rect 6411 17561 6420 17595
rect 6368 17552 6420 17561
rect 7472 17620 7524 17672
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 14096 17620 14148 17672
rect 14924 17663 14976 17672
rect 14924 17629 14933 17663
rect 14933 17629 14967 17663
rect 14967 17629 14976 17663
rect 14924 17620 14976 17629
rect 15292 17620 15344 17672
rect 8300 17552 8352 17604
rect 8484 17552 8536 17604
rect 8576 17552 8628 17604
rect 10508 17552 10560 17604
rect 11152 17552 11204 17604
rect 12164 17552 12216 17604
rect 12808 17552 12860 17604
rect 13544 17595 13596 17604
rect 13544 17561 13553 17595
rect 13553 17561 13587 17595
rect 13587 17561 13596 17595
rect 13544 17552 13596 17561
rect 15568 17595 15620 17604
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 7196 17484 7248 17536
rect 7840 17484 7892 17536
rect 10232 17484 10284 17536
rect 13176 17484 13228 17536
rect 13452 17484 13504 17536
rect 15568 17561 15577 17595
rect 15577 17561 15611 17595
rect 15611 17561 15620 17595
rect 15568 17552 15620 17561
rect 19984 17688 20036 17740
rect 16948 17620 17000 17672
rect 17316 17663 17368 17672
rect 17316 17629 17325 17663
rect 17325 17629 17359 17663
rect 17359 17629 17368 17663
rect 17316 17620 17368 17629
rect 20904 17688 20956 17740
rect 22376 17688 22428 17740
rect 24768 17688 24820 17740
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 23572 17663 23624 17672
rect 23572 17629 23581 17663
rect 23581 17629 23615 17663
rect 23615 17629 23624 17663
rect 23572 17620 23624 17629
rect 20536 17595 20588 17604
rect 20536 17561 20545 17595
rect 20545 17561 20579 17595
rect 20579 17561 20588 17595
rect 20536 17552 20588 17561
rect 21456 17552 21508 17604
rect 23848 17620 23900 17672
rect 25136 17620 25188 17672
rect 25596 17620 25648 17672
rect 26148 17620 26200 17672
rect 34796 17552 34848 17604
rect 17776 17484 17828 17536
rect 18144 17484 18196 17536
rect 21272 17484 21324 17536
rect 25504 17484 25556 17536
rect 33784 17484 33836 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 8668 17280 8720 17332
rect 8944 17280 8996 17332
rect 2136 17255 2188 17264
rect 2136 17221 2145 17255
rect 2145 17221 2179 17255
rect 2179 17221 2188 17255
rect 2136 17212 2188 17221
rect 3148 17212 3200 17264
rect 3792 17212 3844 17264
rect 7012 17212 7064 17264
rect 7656 17212 7708 17264
rect 9404 17212 9456 17264
rect 10232 17280 10284 17332
rect 11980 17255 12032 17264
rect 11980 17221 11989 17255
rect 11989 17221 12023 17255
rect 12023 17221 12032 17255
rect 11980 17212 12032 17221
rect 14832 17212 14884 17264
rect 4804 17144 4856 17196
rect 4896 17144 4948 17196
rect 3332 17076 3384 17128
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 6644 17144 6696 17196
rect 7196 17144 7248 17196
rect 9128 17144 9180 17196
rect 9496 17144 9548 17196
rect 10876 17144 10928 17196
rect 13084 17144 13136 17196
rect 7380 17119 7432 17128
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 6552 17008 6604 17060
rect 4068 16940 4120 16992
rect 5356 16983 5408 16992
rect 5356 16949 5365 16983
rect 5365 16949 5399 16983
rect 5399 16949 5408 16983
rect 5356 16940 5408 16949
rect 6644 16940 6696 16992
rect 10600 17076 10652 17128
rect 10692 17076 10744 17128
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 15476 17144 15528 17153
rect 16488 17212 16540 17264
rect 17224 17187 17276 17196
rect 17224 17153 17233 17187
rect 17233 17153 17267 17187
rect 17267 17153 17276 17187
rect 17224 17144 17276 17153
rect 17868 17187 17920 17196
rect 17868 17153 17877 17187
rect 17877 17153 17911 17187
rect 17911 17153 17920 17187
rect 17868 17144 17920 17153
rect 20720 17212 20772 17264
rect 20904 17212 20956 17264
rect 22192 17323 22244 17332
rect 22192 17289 22201 17323
rect 22201 17289 22235 17323
rect 22235 17289 22244 17323
rect 22652 17323 22704 17332
rect 22192 17280 22244 17289
rect 22652 17289 22661 17323
rect 22661 17289 22695 17323
rect 22695 17289 22704 17323
rect 22652 17280 22704 17289
rect 26240 17280 26292 17332
rect 25136 17255 25188 17264
rect 20076 17144 20128 17196
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 25136 17221 25145 17255
rect 25145 17221 25179 17255
rect 25179 17221 25188 17255
rect 25136 17212 25188 17221
rect 26148 17187 26200 17196
rect 26148 17153 26157 17187
rect 26157 17153 26191 17187
rect 26191 17153 26200 17187
rect 26148 17144 26200 17153
rect 33784 17187 33836 17196
rect 33784 17153 33793 17187
rect 33793 17153 33827 17187
rect 33827 17153 33836 17187
rect 33784 17144 33836 17153
rect 13452 17119 13504 17128
rect 13452 17085 13461 17119
rect 13461 17085 13495 17119
rect 13495 17085 13504 17119
rect 13452 17076 13504 17085
rect 14004 17076 14056 17128
rect 15384 17076 15436 17128
rect 11612 17008 11664 17060
rect 9128 16983 9180 16992
rect 9128 16949 9137 16983
rect 9137 16949 9171 16983
rect 9171 16949 9180 16983
rect 9128 16940 9180 16949
rect 9220 16940 9272 16992
rect 11980 16940 12032 16992
rect 12348 16940 12400 16992
rect 17316 17008 17368 17060
rect 17684 17008 17736 17060
rect 16672 16940 16724 16992
rect 17960 17076 18012 17128
rect 19156 17119 19208 17128
rect 19156 17085 19165 17119
rect 19165 17085 19199 17119
rect 19199 17085 19208 17119
rect 19156 17076 19208 17085
rect 21732 17076 21784 17128
rect 24492 17119 24544 17128
rect 17868 17008 17920 17060
rect 19432 17008 19484 17060
rect 20996 16940 21048 16992
rect 21824 16940 21876 16992
rect 24124 16983 24176 16992
rect 24124 16949 24133 16983
rect 24133 16949 24167 16983
rect 24167 16949 24176 16983
rect 24124 16940 24176 16949
rect 24492 17085 24501 17119
rect 24501 17085 24535 17119
rect 24535 17085 24544 17119
rect 24492 17076 24544 17085
rect 24584 17076 24636 17128
rect 25320 17119 25372 17128
rect 25320 17085 25329 17119
rect 25329 17085 25363 17119
rect 25363 17085 25372 17119
rect 25320 17076 25372 17085
rect 38200 17051 38252 17060
rect 38200 17017 38209 17051
rect 38209 17017 38243 17051
rect 38243 17017 38252 17051
rect 38200 17008 38252 17017
rect 27160 16983 27212 16992
rect 27160 16949 27169 16983
rect 27169 16949 27203 16983
rect 27203 16949 27212 16983
rect 27160 16940 27212 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1676 16736 1728 16788
rect 4068 16600 4120 16652
rect 4620 16736 4672 16788
rect 4896 16736 4948 16788
rect 9128 16736 9180 16788
rect 9496 16736 9548 16788
rect 11704 16736 11756 16788
rect 11980 16736 12032 16788
rect 15384 16736 15436 16788
rect 15476 16736 15528 16788
rect 17224 16736 17276 16788
rect 23572 16736 23624 16788
rect 24124 16736 24176 16788
rect 24584 16779 24636 16788
rect 24584 16745 24593 16779
rect 24593 16745 24627 16779
rect 24627 16745 24636 16779
rect 24584 16736 24636 16745
rect 25136 16736 25188 16788
rect 7012 16668 7064 16720
rect 8944 16668 8996 16720
rect 4804 16600 4856 16652
rect 9312 16600 9364 16652
rect 14004 16668 14056 16720
rect 14372 16668 14424 16720
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 11612 16600 11664 16652
rect 16396 16668 16448 16720
rect 21640 16668 21692 16720
rect 6828 16575 6880 16584
rect 6828 16541 6837 16575
rect 6837 16541 6871 16575
rect 6871 16541 6880 16575
rect 6828 16532 6880 16541
rect 8852 16532 8904 16584
rect 9220 16532 9272 16584
rect 9496 16532 9548 16584
rect 14188 16532 14240 16584
rect 18696 16600 18748 16652
rect 3608 16464 3660 16516
rect 3332 16396 3384 16448
rect 4528 16464 4580 16516
rect 5908 16464 5960 16516
rect 4068 16396 4120 16448
rect 8208 16396 8260 16448
rect 10508 16464 10560 16516
rect 11612 16507 11664 16516
rect 11612 16473 11621 16507
rect 11621 16473 11655 16507
rect 11655 16473 11664 16507
rect 11612 16464 11664 16473
rect 12624 16464 12676 16516
rect 15936 16532 15988 16584
rect 16488 16575 16540 16584
rect 16488 16541 16497 16575
rect 16497 16541 16531 16575
rect 16531 16541 16540 16575
rect 16488 16532 16540 16541
rect 15200 16507 15252 16516
rect 10876 16396 10928 16448
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 13820 16396 13872 16448
rect 15200 16473 15209 16507
rect 15209 16473 15243 16507
rect 15243 16473 15252 16507
rect 15200 16464 15252 16473
rect 15384 16464 15436 16516
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 18972 16600 19024 16652
rect 22652 16600 22704 16652
rect 34244 16668 34296 16720
rect 21456 16575 21508 16584
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 21456 16532 21508 16541
rect 21548 16575 21600 16584
rect 21548 16541 21557 16575
rect 21557 16541 21591 16575
rect 21591 16541 21600 16575
rect 23756 16600 23808 16652
rect 23848 16600 23900 16652
rect 25504 16600 25556 16652
rect 21548 16532 21600 16541
rect 25044 16575 25096 16584
rect 18236 16464 18288 16516
rect 18328 16464 18380 16516
rect 22008 16464 22060 16516
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 27160 16532 27212 16584
rect 34796 16532 34848 16584
rect 38108 16600 38160 16652
rect 16948 16396 17000 16448
rect 18880 16396 18932 16448
rect 20628 16439 20680 16448
rect 20628 16405 20637 16439
rect 20637 16405 20671 16439
rect 20671 16405 20680 16439
rect 20628 16396 20680 16405
rect 22652 16396 22704 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 1584 16192 1636 16244
rect 3884 16192 3936 16244
rect 5080 16124 5132 16176
rect 1952 16056 2004 16108
rect 4528 16056 4580 16108
rect 6828 16192 6880 16244
rect 13728 16192 13780 16244
rect 22652 16235 22704 16244
rect 2872 16031 2924 16040
rect 2872 15997 2881 16031
rect 2881 15997 2915 16031
rect 2915 15997 2924 16031
rect 2872 15988 2924 15997
rect 3240 15988 3292 16040
rect 4896 16031 4948 16040
rect 4896 15997 4905 16031
rect 4905 15997 4939 16031
rect 4939 15997 4948 16031
rect 4896 15988 4948 15997
rect 6552 15988 6604 16040
rect 7840 16124 7892 16176
rect 8760 16124 8812 16176
rect 9772 16124 9824 16176
rect 10232 16167 10284 16176
rect 10232 16133 10241 16167
rect 10241 16133 10275 16167
rect 10275 16133 10284 16167
rect 10232 16124 10284 16133
rect 2320 15852 2372 15904
rect 9128 16056 9180 16108
rect 11704 16099 11756 16108
rect 7380 15988 7432 16040
rect 7748 16031 7800 16040
rect 6920 15963 6972 15972
rect 6920 15929 6929 15963
rect 6929 15929 6963 15963
rect 6963 15929 6972 15963
rect 6920 15920 6972 15929
rect 7104 15852 7156 15904
rect 7748 15997 7757 16031
rect 7757 15997 7791 16031
rect 7791 15997 7800 16031
rect 7748 15988 7800 15997
rect 8116 15988 8168 16040
rect 9680 15988 9732 16040
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 13728 15988 13780 16040
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 13912 15988 13964 15997
rect 14004 15988 14056 16040
rect 15936 16124 15988 16176
rect 16396 16124 16448 16176
rect 16672 16056 16724 16108
rect 16028 15988 16080 16040
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 16580 15988 16632 16040
rect 17684 15988 17736 16040
rect 10324 15920 10376 15972
rect 10876 15920 10928 15972
rect 11980 15920 12032 15972
rect 8208 15852 8260 15904
rect 9128 15852 9180 15904
rect 9404 15852 9456 15904
rect 13544 15852 13596 15904
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 14556 15920 14608 15972
rect 18420 15988 18472 16040
rect 20628 16124 20680 16176
rect 20904 16167 20956 16176
rect 20904 16133 20913 16167
rect 20913 16133 20947 16167
rect 20947 16133 20956 16167
rect 22652 16201 22661 16235
rect 22661 16201 22695 16235
rect 22695 16201 22704 16235
rect 22652 16192 22704 16201
rect 22744 16192 22796 16244
rect 23756 16235 23808 16244
rect 23756 16201 23765 16235
rect 23765 16201 23799 16235
rect 23799 16201 23808 16235
rect 23756 16192 23808 16201
rect 25044 16235 25096 16244
rect 25044 16201 25053 16235
rect 25053 16201 25087 16235
rect 25087 16201 25096 16235
rect 25044 16192 25096 16201
rect 20904 16124 20956 16133
rect 21548 16056 21600 16108
rect 18144 15963 18196 15972
rect 18144 15929 18153 15963
rect 18153 15929 18187 15963
rect 18187 15929 18196 15963
rect 18144 15920 18196 15929
rect 21456 15920 21508 15972
rect 21916 15988 21968 16040
rect 22192 16031 22244 16040
rect 22192 15997 22201 16031
rect 22201 15997 22235 16031
rect 22235 15997 22244 16031
rect 22192 15988 22244 15997
rect 22468 15988 22520 16040
rect 24308 15988 24360 16040
rect 23756 15920 23808 15972
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 16488 15852 16540 15904
rect 22560 15852 22612 15904
rect 26148 16056 26200 16108
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3240 15648 3292 15700
rect 11612 15648 11664 15700
rect 14280 15648 14332 15700
rect 14556 15691 14608 15700
rect 14556 15657 14565 15691
rect 14565 15657 14599 15691
rect 14599 15657 14608 15691
rect 14556 15648 14608 15657
rect 14648 15648 14700 15700
rect 16580 15648 16632 15700
rect 18328 15648 18380 15700
rect 20076 15691 20128 15700
rect 20076 15657 20085 15691
rect 20085 15657 20119 15691
rect 20119 15657 20128 15691
rect 20076 15648 20128 15657
rect 20536 15648 20588 15700
rect 22192 15648 22244 15700
rect 38108 15691 38160 15700
rect 38108 15657 38117 15691
rect 38117 15657 38151 15691
rect 38151 15657 38160 15691
rect 38108 15648 38160 15657
rect 2872 15512 2924 15564
rect 3608 15512 3660 15564
rect 6736 15580 6788 15632
rect 8944 15580 8996 15632
rect 10508 15580 10560 15632
rect 22560 15580 22612 15632
rect 27436 15580 27488 15632
rect 12348 15555 12400 15564
rect 3884 15376 3936 15428
rect 4896 15444 4948 15496
rect 6920 15444 6972 15496
rect 5264 15376 5316 15428
rect 5540 15419 5592 15428
rect 5540 15385 5549 15419
rect 5549 15385 5583 15419
rect 5583 15385 5592 15419
rect 5540 15376 5592 15385
rect 6000 15376 6052 15428
rect 7288 15419 7340 15428
rect 7288 15385 7297 15419
rect 7297 15385 7331 15419
rect 7331 15385 7340 15419
rect 7288 15376 7340 15385
rect 7472 15444 7524 15496
rect 8852 15444 8904 15496
rect 8944 15376 8996 15428
rect 10140 15376 10192 15428
rect 4068 15308 4120 15360
rect 8392 15308 8444 15360
rect 8484 15308 8536 15360
rect 9680 15308 9732 15360
rect 10416 15308 10468 15360
rect 12348 15521 12357 15555
rect 12357 15521 12391 15555
rect 12391 15521 12400 15555
rect 12348 15512 12400 15521
rect 13820 15512 13872 15564
rect 14188 15512 14240 15564
rect 15476 15512 15528 15564
rect 16396 15512 16448 15564
rect 18972 15512 19024 15564
rect 21180 15555 21232 15564
rect 21180 15521 21189 15555
rect 21189 15521 21223 15555
rect 21223 15521 21232 15555
rect 21180 15512 21232 15521
rect 21456 15555 21508 15564
rect 21456 15521 21465 15555
rect 21465 15521 21499 15555
rect 21499 15521 21508 15555
rect 23112 15555 23164 15564
rect 21456 15512 21508 15521
rect 23112 15521 23121 15555
rect 23121 15521 23155 15555
rect 23155 15521 23164 15555
rect 23112 15512 23164 15521
rect 16764 15487 16816 15496
rect 11520 15376 11572 15428
rect 12072 15376 12124 15428
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 24032 15487 24084 15496
rect 15108 15419 15160 15428
rect 15108 15385 15117 15419
rect 15117 15385 15151 15419
rect 15151 15385 15160 15419
rect 15108 15376 15160 15385
rect 15292 15376 15344 15428
rect 17408 15419 17460 15428
rect 17408 15385 17417 15419
rect 17417 15385 17451 15419
rect 17451 15385 17460 15419
rect 17408 15376 17460 15385
rect 17776 15308 17828 15360
rect 20352 15376 20404 15428
rect 18144 15308 18196 15360
rect 24032 15453 24041 15487
rect 24041 15453 24075 15487
rect 24075 15453 24084 15487
rect 24032 15444 24084 15453
rect 24584 15487 24636 15496
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 24584 15444 24636 15453
rect 38292 15487 38344 15496
rect 38292 15453 38301 15487
rect 38301 15453 38335 15487
rect 38335 15453 38344 15487
rect 38292 15444 38344 15453
rect 21272 15419 21324 15428
rect 21272 15385 21281 15419
rect 21281 15385 21315 15419
rect 21315 15385 21324 15419
rect 22744 15419 22796 15428
rect 21272 15376 21324 15385
rect 22744 15385 22753 15419
rect 22753 15385 22787 15419
rect 22787 15385 22796 15419
rect 22744 15376 22796 15385
rect 22468 15308 22520 15360
rect 23664 15308 23716 15360
rect 23848 15351 23900 15360
rect 23848 15317 23857 15351
rect 23857 15317 23891 15351
rect 23891 15317 23900 15351
rect 23848 15308 23900 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2044 15104 2096 15156
rect 3700 15104 3752 15156
rect 11704 15104 11756 15156
rect 3792 15036 3844 15088
rect 4896 15036 4948 15088
rect 1768 14968 1820 15020
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 3608 15011 3660 15020
rect 2780 14764 2832 14816
rect 3608 14977 3617 15011
rect 3617 14977 3651 15011
rect 3651 14977 3660 15011
rect 3608 14968 3660 14977
rect 6920 15036 6972 15088
rect 9036 15036 9088 15088
rect 10968 15036 11020 15088
rect 12256 15079 12308 15088
rect 12256 15045 12265 15079
rect 12265 15045 12299 15079
rect 12299 15045 12308 15079
rect 12256 15036 12308 15045
rect 16764 15104 16816 15156
rect 17592 15104 17644 15156
rect 5264 14832 5316 14884
rect 7932 14968 7984 15020
rect 10508 14968 10560 15020
rect 6460 14900 6512 14952
rect 7840 14900 7892 14952
rect 8852 14943 8904 14952
rect 6276 14764 6328 14816
rect 7380 14764 7432 14816
rect 8852 14909 8861 14943
rect 8861 14909 8895 14943
rect 8895 14909 8904 14943
rect 8852 14900 8904 14909
rect 9220 14900 9272 14952
rect 11060 14900 11112 14952
rect 14188 15036 14240 15088
rect 14280 15036 14332 15088
rect 16948 15036 17000 15088
rect 12992 14968 13044 15020
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 13084 14943 13136 14952
rect 12900 14900 12952 14909
rect 13084 14909 13093 14943
rect 13093 14909 13127 14943
rect 13127 14909 13136 14943
rect 13084 14900 13136 14909
rect 13820 14900 13872 14952
rect 14556 14900 14608 14952
rect 14832 14900 14884 14952
rect 16672 14968 16724 15020
rect 18052 15036 18104 15088
rect 20076 15104 20128 15156
rect 20904 15104 20956 15156
rect 20168 15036 20220 15088
rect 21180 14968 21232 15020
rect 23848 15104 23900 15156
rect 24584 15036 24636 15088
rect 23572 14968 23624 15020
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 17868 14943 17920 14952
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 17868 14900 17920 14909
rect 18236 14900 18288 14952
rect 19064 14943 19116 14952
rect 19064 14909 19073 14943
rect 19073 14909 19107 14943
rect 19107 14909 19116 14943
rect 19064 14900 19116 14909
rect 20812 14943 20864 14952
rect 10232 14832 10284 14884
rect 11520 14832 11572 14884
rect 13360 14832 13412 14884
rect 9864 14764 9916 14816
rect 10508 14764 10560 14816
rect 11060 14764 11112 14816
rect 13728 14764 13780 14816
rect 15108 14807 15160 14816
rect 15108 14773 15117 14807
rect 15117 14773 15151 14807
rect 15151 14773 15160 14807
rect 15108 14764 15160 14773
rect 18788 14832 18840 14884
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 23112 14943 23164 14952
rect 23112 14909 23121 14943
rect 23121 14909 23155 14943
rect 23155 14909 23164 14943
rect 23112 14900 23164 14909
rect 23296 14900 23348 14952
rect 23664 14900 23716 14952
rect 19432 14764 19484 14816
rect 19984 14764 20036 14816
rect 21548 14764 21600 14816
rect 29276 14807 29328 14816
rect 29276 14773 29285 14807
rect 29285 14773 29319 14807
rect 29319 14773 29328 14807
rect 29276 14764 29328 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2780 14560 2832 14612
rect 4436 14560 4488 14612
rect 10048 14560 10100 14612
rect 10876 14603 10928 14612
rect 10876 14569 10885 14603
rect 10885 14569 10919 14603
rect 10919 14569 10928 14603
rect 10876 14560 10928 14569
rect 12348 14560 12400 14612
rect 14556 14560 14608 14612
rect 15108 14560 15160 14612
rect 17776 14560 17828 14612
rect 20260 14560 20312 14612
rect 20444 14560 20496 14612
rect 21272 14560 21324 14612
rect 21456 14560 21508 14612
rect 24584 14603 24636 14612
rect 3056 14492 3108 14544
rect 5264 14492 5316 14544
rect 7840 14492 7892 14544
rect 1676 14467 1728 14476
rect 1676 14433 1685 14467
rect 1685 14433 1719 14467
rect 1719 14433 1728 14467
rect 1676 14424 1728 14433
rect 7012 14424 7064 14476
rect 7380 14424 7432 14476
rect 9036 14424 9088 14476
rect 10600 14424 10652 14476
rect 10876 14424 10928 14476
rect 11612 14424 11664 14476
rect 12164 14467 12216 14476
rect 12164 14433 12173 14467
rect 12173 14433 12207 14467
rect 12207 14433 12216 14467
rect 12164 14424 12216 14433
rect 12624 14492 12676 14544
rect 12900 14492 12952 14544
rect 13360 14424 13412 14476
rect 13636 14492 13688 14544
rect 15200 14492 15252 14544
rect 15476 14535 15528 14544
rect 15476 14501 15485 14535
rect 15485 14501 15519 14535
rect 15519 14501 15528 14535
rect 15476 14492 15528 14501
rect 16028 14492 16080 14544
rect 17592 14492 17644 14544
rect 18788 14492 18840 14544
rect 24308 14492 24360 14544
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 25228 14603 25280 14612
rect 25228 14569 25237 14603
rect 25237 14569 25271 14603
rect 25271 14569 25280 14603
rect 25228 14560 25280 14569
rect 26148 14492 26200 14544
rect 14648 14424 14700 14476
rect 18420 14424 18472 14476
rect 2964 14356 3016 14408
rect 3240 14288 3292 14340
rect 4620 14356 4672 14408
rect 4804 14399 4856 14408
rect 4804 14365 4813 14399
rect 4813 14365 4847 14399
rect 4847 14365 4856 14399
rect 4804 14356 4856 14365
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 12900 14356 12952 14408
rect 14188 14356 14240 14408
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 16580 14399 16632 14408
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 17316 14356 17368 14408
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 20720 14399 20772 14408
rect 5724 14288 5776 14340
rect 7380 14331 7432 14340
rect 7380 14297 7389 14331
rect 7389 14297 7423 14331
rect 7423 14297 7432 14331
rect 7380 14288 7432 14297
rect 8116 14288 8168 14340
rect 9128 14288 9180 14340
rect 9404 14331 9456 14340
rect 9404 14297 9413 14331
rect 9413 14297 9447 14331
rect 9447 14297 9456 14331
rect 9404 14288 9456 14297
rect 9956 14288 10008 14340
rect 8576 14263 8628 14272
rect 8576 14229 8585 14263
rect 8585 14229 8619 14263
rect 8619 14229 8628 14263
rect 8576 14220 8628 14229
rect 9588 14220 9640 14272
rect 11520 14220 11572 14272
rect 12164 14288 12216 14340
rect 11980 14220 12032 14272
rect 13820 14220 13872 14272
rect 15200 14288 15252 14340
rect 17408 14288 17460 14340
rect 14556 14220 14608 14272
rect 16396 14220 16448 14272
rect 19984 14288 20036 14340
rect 20720 14365 20729 14399
rect 20729 14365 20763 14399
rect 20763 14365 20772 14399
rect 20720 14356 20772 14365
rect 21732 14424 21784 14476
rect 21548 14356 21600 14408
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 23296 14399 23348 14408
rect 23296 14365 23305 14399
rect 23305 14365 23339 14399
rect 23339 14365 23348 14399
rect 23296 14356 23348 14365
rect 23480 14356 23532 14408
rect 25228 14356 25280 14408
rect 36912 14356 36964 14408
rect 18512 14220 18564 14272
rect 18604 14220 18656 14272
rect 19248 14220 19300 14272
rect 21456 14220 21508 14272
rect 22376 14220 22428 14272
rect 24768 14220 24820 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1676 14016 1728 14068
rect 1308 13948 1360 14000
rect 3516 13948 3568 14000
rect 4712 14016 4764 14068
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 8576 14016 8628 14068
rect 13636 14059 13688 14068
rect 5356 13948 5408 14000
rect 5816 13948 5868 14000
rect 8208 13948 8260 14000
rect 9312 13991 9364 14000
rect 9312 13957 9321 13991
rect 9321 13957 9355 13991
rect 9355 13957 9364 13991
rect 9312 13948 9364 13957
rect 11612 13948 11664 14000
rect 13636 14025 13645 14059
rect 13645 14025 13679 14059
rect 13679 14025 13688 14059
rect 13636 14016 13688 14025
rect 16120 14016 16172 14068
rect 16856 14059 16908 14068
rect 16856 14025 16865 14059
rect 16865 14025 16899 14059
rect 16899 14025 16908 14059
rect 16856 14016 16908 14025
rect 17960 14059 18012 14068
rect 17960 14025 17969 14059
rect 17969 14025 18003 14059
rect 18003 14025 18012 14059
rect 17960 14016 18012 14025
rect 19156 14016 19208 14068
rect 19984 14059 20036 14068
rect 19984 14025 19993 14059
rect 19993 14025 20027 14059
rect 20027 14025 20036 14059
rect 19984 14016 20036 14025
rect 22376 14016 22428 14068
rect 14096 13948 14148 14000
rect 14924 13991 14976 14000
rect 14924 13957 14933 13991
rect 14933 13957 14967 13991
rect 14967 13957 14976 13991
rect 14924 13948 14976 13957
rect 17316 13948 17368 14000
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 10416 13880 10468 13932
rect 12532 13880 12584 13932
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 4436 13812 4488 13864
rect 11152 13812 11204 13864
rect 11520 13812 11572 13864
rect 11980 13812 12032 13864
rect 12716 13812 12768 13864
rect 13636 13812 13688 13864
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 14464 13812 14516 13864
rect 15108 13812 15160 13864
rect 6092 13744 6144 13796
rect 10324 13744 10376 13796
rect 1676 13676 1728 13728
rect 6276 13676 6328 13728
rect 8208 13676 8260 13728
rect 8668 13676 8720 13728
rect 9312 13676 9364 13728
rect 15660 13744 15712 13796
rect 16028 13880 16080 13932
rect 18328 13880 18380 13932
rect 19248 13880 19300 13932
rect 21548 13948 21600 14000
rect 24032 14016 24084 14068
rect 24308 14016 24360 14068
rect 27620 14016 27672 14068
rect 23572 13948 23624 14000
rect 23480 13923 23532 13932
rect 23480 13889 23489 13923
rect 23489 13889 23523 13923
rect 23523 13889 23532 13923
rect 23480 13880 23532 13889
rect 29276 13880 29328 13932
rect 19432 13812 19484 13864
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 22560 13812 22612 13864
rect 13176 13719 13228 13728
rect 13176 13685 13185 13719
rect 13185 13685 13219 13719
rect 13219 13685 13228 13719
rect 13176 13676 13228 13685
rect 13360 13676 13412 13728
rect 14372 13676 14424 13728
rect 14648 13676 14700 13728
rect 21916 13676 21968 13728
rect 22284 13676 22336 13728
rect 38200 13719 38252 13728
rect 38200 13685 38209 13719
rect 38209 13685 38243 13719
rect 38243 13685 38252 13719
rect 38200 13676 38252 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2228 13472 2280 13524
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 2872 13336 2924 13388
rect 4712 13336 4764 13388
rect 7472 13404 7524 13456
rect 5448 13268 5500 13320
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 10692 13472 10744 13524
rect 11888 13472 11940 13524
rect 12900 13472 12952 13524
rect 13452 13472 13504 13524
rect 9036 13336 9088 13388
rect 10784 13336 10836 13388
rect 13360 13404 13412 13456
rect 16028 13404 16080 13456
rect 13728 13336 13780 13388
rect 15200 13336 15252 13388
rect 15568 13336 15620 13388
rect 15844 13336 15896 13388
rect 16764 13379 16816 13388
rect 16764 13345 16773 13379
rect 16773 13345 16807 13379
rect 16807 13345 16816 13379
rect 16764 13336 16816 13345
rect 23388 13472 23440 13524
rect 23572 13472 23624 13524
rect 26148 13472 26200 13524
rect 7288 13268 7340 13277
rect 8300 13268 8352 13320
rect 8484 13268 8536 13320
rect 10692 13268 10744 13320
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 17960 13268 18012 13320
rect 1768 13200 1820 13252
rect 1400 13132 1452 13184
rect 6460 13200 6512 13252
rect 8116 13200 8168 13252
rect 9312 13200 9364 13252
rect 10048 13200 10100 13252
rect 4068 13175 4120 13184
rect 4068 13141 4077 13175
rect 4077 13141 4111 13175
rect 4111 13141 4120 13175
rect 4068 13132 4120 13141
rect 6092 13132 6144 13184
rect 7288 13132 7340 13184
rect 8484 13132 8536 13184
rect 8576 13132 8628 13184
rect 12716 13200 12768 13252
rect 12900 13200 12952 13252
rect 13360 13200 13412 13252
rect 14648 13243 14700 13252
rect 14648 13209 14657 13243
rect 14657 13209 14691 13243
rect 14691 13209 14700 13243
rect 14648 13200 14700 13209
rect 15660 13200 15712 13252
rect 24768 13404 24820 13456
rect 19524 13336 19576 13388
rect 19984 13268 20036 13320
rect 20168 13268 20220 13320
rect 20812 13336 20864 13388
rect 22376 13379 22428 13388
rect 22376 13345 22385 13379
rect 22385 13345 22419 13379
rect 22419 13345 22428 13379
rect 22376 13336 22428 13345
rect 22560 13336 22612 13388
rect 23020 13336 23072 13388
rect 23664 13311 23716 13320
rect 23664 13277 23673 13311
rect 23673 13277 23707 13311
rect 23707 13277 23716 13311
rect 23664 13268 23716 13277
rect 30748 13311 30800 13320
rect 30748 13277 30757 13311
rect 30757 13277 30791 13311
rect 30791 13277 30800 13311
rect 30748 13268 30800 13277
rect 10784 13132 10836 13184
rect 12164 13132 12216 13184
rect 12348 13132 12400 13184
rect 22836 13200 22888 13252
rect 18328 13175 18380 13184
rect 18328 13141 18337 13175
rect 18337 13141 18371 13175
rect 18371 13141 18380 13175
rect 18328 13132 18380 13141
rect 21088 13132 21140 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 8576 12928 8628 12980
rect 9036 12928 9088 12980
rect 3332 12903 3384 12912
rect 3332 12869 3341 12903
rect 3341 12869 3375 12903
rect 3375 12869 3384 12903
rect 3332 12860 3384 12869
rect 3700 12860 3752 12912
rect 6276 12860 6328 12912
rect 6736 12860 6788 12912
rect 2228 12792 2280 12844
rect 1492 12724 1544 12776
rect 2872 12724 2924 12776
rect 6828 12792 6880 12844
rect 7104 12792 7156 12844
rect 7288 12792 7340 12844
rect 10600 12928 10652 12980
rect 11520 12928 11572 12980
rect 11888 12928 11940 12980
rect 12164 12928 12216 12980
rect 12624 12860 12676 12912
rect 12716 12860 12768 12912
rect 14556 12860 14608 12912
rect 3516 12588 3568 12640
rect 4068 12588 4120 12640
rect 5540 12588 5592 12640
rect 6092 12724 6144 12776
rect 10416 12724 10468 12776
rect 10600 12724 10652 12776
rect 12164 12792 12216 12844
rect 13176 12792 13228 12844
rect 15752 12928 15804 12980
rect 21180 12928 21232 12980
rect 22468 12928 22520 12980
rect 22836 12928 22888 12980
rect 15568 12903 15620 12912
rect 15568 12869 15577 12903
rect 15577 12869 15611 12903
rect 15611 12869 15620 12903
rect 15568 12860 15620 12869
rect 15660 12860 15712 12912
rect 18236 12860 18288 12912
rect 19248 12860 19300 12912
rect 19524 12903 19576 12912
rect 19524 12869 19533 12903
rect 19533 12869 19567 12903
rect 19567 12869 19576 12903
rect 19524 12860 19576 12869
rect 20904 12903 20956 12912
rect 20904 12869 20913 12903
rect 20913 12869 20947 12903
rect 20947 12869 20956 12903
rect 20904 12860 20956 12869
rect 21640 12860 21692 12912
rect 22284 12792 22336 12844
rect 8944 12656 8996 12708
rect 9404 12656 9456 12708
rect 11152 12656 11204 12708
rect 12348 12724 12400 12776
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 12716 12767 12768 12776
rect 12716 12733 12725 12767
rect 12725 12733 12759 12767
rect 12759 12733 12768 12767
rect 12716 12724 12768 12733
rect 15476 12767 15528 12776
rect 15476 12733 15485 12767
rect 15485 12733 15519 12767
rect 15519 12733 15528 12767
rect 15476 12724 15528 12733
rect 17500 12767 17552 12776
rect 17500 12733 17509 12767
rect 17509 12733 17543 12767
rect 17543 12733 17552 12767
rect 17500 12724 17552 12733
rect 17684 12767 17736 12776
rect 17684 12733 17693 12767
rect 17693 12733 17727 12767
rect 17727 12733 17736 12767
rect 17684 12724 17736 12733
rect 12900 12699 12952 12708
rect 12900 12665 12909 12699
rect 12909 12665 12943 12699
rect 12943 12665 12952 12699
rect 12900 12656 12952 12665
rect 13176 12656 13228 12708
rect 15200 12656 15252 12708
rect 17316 12699 17368 12708
rect 17316 12665 17325 12699
rect 17325 12665 17359 12699
rect 17359 12665 17368 12699
rect 18328 12724 18380 12776
rect 20628 12724 20680 12776
rect 21088 12724 21140 12776
rect 23112 12724 23164 12776
rect 23388 12724 23440 12776
rect 27620 12792 27672 12844
rect 17316 12656 17368 12665
rect 6092 12588 6144 12640
rect 6368 12588 6420 12640
rect 7932 12588 7984 12640
rect 9312 12588 9364 12640
rect 11704 12588 11756 12640
rect 12348 12588 12400 12640
rect 21088 12588 21140 12640
rect 28080 12588 28132 12640
rect 31668 12588 31720 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 6552 12427 6604 12436
rect 2780 12248 2832 12300
rect 3516 12248 3568 12300
rect 3976 12291 4028 12300
rect 3976 12257 3985 12291
rect 3985 12257 4019 12291
rect 4019 12257 4028 12291
rect 3976 12248 4028 12257
rect 5540 12248 5592 12300
rect 3056 12112 3108 12164
rect 4252 12155 4304 12164
rect 4252 12121 4261 12155
rect 4261 12121 4295 12155
rect 4295 12121 4304 12155
rect 4252 12112 4304 12121
rect 4896 12112 4948 12164
rect 5632 12112 5684 12164
rect 1860 12044 1912 12096
rect 5908 12044 5960 12096
rect 6552 12393 6561 12427
rect 6561 12393 6595 12427
rect 6595 12393 6604 12427
rect 6552 12384 6604 12393
rect 6644 12384 6696 12436
rect 11428 12316 11480 12368
rect 13268 12384 13320 12436
rect 15476 12427 15528 12436
rect 15476 12393 15485 12427
rect 15485 12393 15519 12427
rect 15519 12393 15528 12427
rect 15476 12384 15528 12393
rect 16764 12384 16816 12436
rect 17316 12384 17368 12436
rect 18328 12427 18380 12436
rect 18328 12393 18337 12427
rect 18337 12393 18371 12427
rect 18371 12393 18380 12427
rect 18328 12384 18380 12393
rect 19432 12384 19484 12436
rect 20720 12427 20772 12436
rect 20720 12393 20729 12427
rect 20729 12393 20763 12427
rect 20763 12393 20772 12427
rect 20720 12384 20772 12393
rect 20996 12384 21048 12436
rect 7012 12248 7064 12300
rect 7656 12248 7708 12300
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 8484 12248 8536 12300
rect 11244 12248 11296 12300
rect 11704 12248 11756 12300
rect 11888 12248 11940 12300
rect 6920 12180 6972 12232
rect 9036 12180 9088 12232
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 7748 12112 7800 12164
rect 8392 12044 8444 12096
rect 8852 12044 8904 12096
rect 9312 12112 9364 12164
rect 10508 12112 10560 12164
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 15936 12316 15988 12368
rect 20352 12316 20404 12368
rect 21364 12316 21416 12368
rect 23112 12316 23164 12368
rect 30840 12316 30892 12368
rect 15752 12248 15804 12300
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 15108 12223 15160 12232
rect 15108 12189 15117 12223
rect 15117 12189 15151 12223
rect 15151 12189 15160 12223
rect 15108 12180 15160 12189
rect 16488 12223 16540 12232
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 16488 12180 16540 12189
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 18604 12180 18656 12232
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 22008 12248 22060 12300
rect 20352 12223 20404 12232
rect 20352 12189 20361 12223
rect 20361 12189 20395 12223
rect 20395 12189 20404 12223
rect 20352 12180 20404 12189
rect 20444 12180 20496 12232
rect 21640 12223 21692 12232
rect 21640 12189 21649 12223
rect 21649 12189 21683 12223
rect 21683 12189 21692 12223
rect 21640 12180 21692 12189
rect 23388 12112 23440 12164
rect 12900 12044 12952 12096
rect 13636 12044 13688 12096
rect 14556 12044 14608 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2412 11840 2464 11892
rect 2320 11815 2372 11824
rect 2320 11781 2329 11815
rect 2329 11781 2363 11815
rect 2363 11781 2372 11815
rect 2320 11772 2372 11781
rect 4068 11772 4120 11824
rect 4712 11704 4764 11756
rect 6000 11840 6052 11892
rect 5448 11772 5500 11824
rect 7472 11772 7524 11824
rect 10324 11772 10376 11824
rect 5540 11704 5592 11756
rect 5908 11704 5960 11756
rect 7748 11704 7800 11756
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 9772 11704 9824 11756
rect 10876 11704 10928 11756
rect 13176 11840 13228 11892
rect 15016 11840 15068 11892
rect 15476 11840 15528 11892
rect 16212 11840 16264 11892
rect 17868 11840 17920 11892
rect 18512 11840 18564 11892
rect 20168 11840 20220 11892
rect 20444 11883 20496 11892
rect 20444 11849 20453 11883
rect 20453 11849 20487 11883
rect 20487 11849 20496 11883
rect 20444 11840 20496 11849
rect 20904 11840 20956 11892
rect 23388 11883 23440 11892
rect 23388 11849 23397 11883
rect 23397 11849 23431 11883
rect 23431 11849 23440 11883
rect 23388 11840 23440 11849
rect 36912 11840 36964 11892
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 3608 11568 3660 11620
rect 4160 11636 4212 11688
rect 4712 11568 4764 11620
rect 1676 11500 1728 11552
rect 7840 11568 7892 11620
rect 9956 11636 10008 11688
rect 10692 11636 10744 11688
rect 11060 11636 11112 11688
rect 12440 11704 12492 11756
rect 18144 11772 18196 11824
rect 17132 11704 17184 11756
rect 17592 11704 17644 11756
rect 36820 11772 36872 11824
rect 18696 11704 18748 11756
rect 15016 11679 15068 11688
rect 15016 11645 15025 11679
rect 15025 11645 15059 11679
rect 15059 11645 15068 11679
rect 15016 11636 15068 11645
rect 15200 11679 15252 11688
rect 15200 11645 15209 11679
rect 15209 11645 15243 11679
rect 15243 11645 15252 11679
rect 15200 11636 15252 11645
rect 11152 11568 11204 11620
rect 14280 11568 14332 11620
rect 14740 11568 14792 11620
rect 20444 11704 20496 11756
rect 21088 11704 21140 11756
rect 22744 11747 22796 11756
rect 22744 11713 22753 11747
rect 22753 11713 22787 11747
rect 22787 11713 22796 11747
rect 22744 11704 22796 11713
rect 23296 11704 23348 11756
rect 27436 11747 27488 11756
rect 27436 11713 27445 11747
rect 27445 11713 27479 11747
rect 27479 11713 27488 11747
rect 27436 11704 27488 11713
rect 31668 11704 31720 11756
rect 38292 11747 38344 11756
rect 38292 11713 38301 11747
rect 38301 11713 38335 11747
rect 38335 11713 38344 11747
rect 38292 11704 38344 11713
rect 20260 11568 20312 11620
rect 23664 11568 23716 11620
rect 8300 11500 8352 11552
rect 8392 11500 8444 11552
rect 10416 11500 10468 11552
rect 10692 11500 10744 11552
rect 10876 11500 10928 11552
rect 14372 11500 14424 11552
rect 32864 11500 32916 11552
rect 35348 11500 35400 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 3056 11296 3108 11348
rect 3516 11296 3568 11348
rect 10600 11296 10652 11348
rect 11152 11296 11204 11348
rect 11796 11339 11848 11348
rect 11796 11305 11805 11339
rect 11805 11305 11839 11339
rect 11839 11305 11848 11339
rect 11796 11296 11848 11305
rect 14004 11296 14056 11348
rect 15292 11296 15344 11348
rect 15384 11296 15436 11348
rect 16948 11296 17000 11348
rect 18052 11296 18104 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 19432 11296 19484 11348
rect 20444 11339 20496 11348
rect 20444 11305 20453 11339
rect 20453 11305 20487 11339
rect 20487 11305 20496 11339
rect 20444 11296 20496 11305
rect 2780 11160 2832 11212
rect 6276 11160 6328 11212
rect 7656 11160 7708 11212
rect 8300 11203 8352 11212
rect 8300 11169 8309 11203
rect 8309 11169 8343 11203
rect 8343 11169 8352 11203
rect 11428 11228 11480 11280
rect 13912 11228 13964 11280
rect 19064 11228 19116 11280
rect 8300 11160 8352 11169
rect 3976 11092 4028 11144
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 9404 11092 9456 11144
rect 9496 11092 9548 11144
rect 10232 11092 10284 11144
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 11888 11135 11940 11144
rect 2688 11024 2740 11076
rect 3792 11024 3844 11076
rect 5172 11024 5224 11076
rect 5632 11024 5684 11076
rect 4712 10956 4764 11008
rect 6460 11024 6512 11076
rect 8668 11024 8720 11076
rect 8852 11024 8904 11076
rect 8484 10956 8536 11008
rect 9496 10956 9548 11008
rect 10048 11024 10100 11076
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 14556 11092 14608 11144
rect 17868 11160 17920 11212
rect 16948 11092 17000 11144
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 10876 11024 10928 11076
rect 17132 11024 17184 11076
rect 19984 11092 20036 11144
rect 20260 11135 20312 11144
rect 20260 11101 20269 11135
rect 20269 11101 20303 11135
rect 20303 11101 20312 11135
rect 20260 11092 20312 11101
rect 10968 10956 11020 11008
rect 11152 10956 11204 11008
rect 12072 10956 12124 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 2780 10752 2832 10804
rect 2872 10752 2924 10804
rect 6644 10795 6696 10804
rect 1952 10727 2004 10736
rect 1952 10693 1961 10727
rect 1961 10693 1995 10727
rect 1995 10693 2004 10727
rect 1952 10684 2004 10693
rect 6276 10684 6328 10736
rect 6644 10761 6653 10795
rect 6653 10761 6687 10795
rect 6687 10761 6696 10795
rect 6644 10752 6696 10761
rect 6828 10752 6880 10804
rect 7288 10684 7340 10736
rect 6000 10659 6052 10668
rect 6000 10625 6009 10659
rect 6009 10625 6043 10659
rect 6043 10625 6052 10659
rect 6000 10616 6052 10625
rect 5264 10548 5316 10600
rect 6644 10616 6696 10668
rect 9680 10684 9732 10736
rect 11520 10752 11572 10804
rect 11888 10752 11940 10804
rect 8024 10616 8076 10668
rect 9404 10659 9456 10668
rect 9404 10625 9413 10659
rect 9413 10625 9447 10659
rect 9447 10625 9456 10659
rect 9404 10616 9456 10625
rect 10508 10616 10560 10668
rect 11152 10684 11204 10736
rect 11244 10684 11296 10736
rect 11520 10616 11572 10668
rect 11796 10684 11848 10736
rect 12992 10752 13044 10804
rect 14096 10752 14148 10804
rect 14832 10795 14884 10804
rect 14832 10761 14841 10795
rect 14841 10761 14875 10795
rect 14875 10761 14884 10795
rect 14832 10752 14884 10761
rect 16120 10752 16172 10804
rect 16580 10752 16632 10804
rect 17500 10752 17552 10804
rect 18052 10795 18104 10804
rect 18052 10761 18061 10795
rect 18061 10761 18095 10795
rect 18095 10761 18104 10795
rect 18052 10752 18104 10761
rect 18880 10795 18932 10804
rect 18880 10761 18889 10795
rect 18889 10761 18923 10795
rect 18923 10761 18932 10795
rect 18880 10752 18932 10761
rect 19984 10752 20036 10804
rect 11888 10616 11940 10668
rect 15936 10684 15988 10736
rect 13912 10616 13964 10668
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 14556 10616 14608 10668
rect 16396 10616 16448 10668
rect 17868 10659 17920 10668
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 2412 10412 2464 10464
rect 5632 10412 5684 10464
rect 6092 10412 6144 10464
rect 17684 10548 17736 10600
rect 28080 10616 28132 10668
rect 35348 10616 35400 10668
rect 10416 10480 10468 10532
rect 11796 10480 11848 10532
rect 9496 10412 9548 10464
rect 13268 10412 13320 10464
rect 18880 10412 18932 10464
rect 30104 10455 30156 10464
rect 30104 10421 30113 10455
rect 30113 10421 30147 10455
rect 30147 10421 30156 10455
rect 30104 10412 30156 10421
rect 38200 10455 38252 10464
rect 38200 10421 38209 10455
rect 38209 10421 38243 10455
rect 38243 10421 38252 10455
rect 38200 10412 38252 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1492 10208 1544 10260
rect 6092 10208 6144 10260
rect 6184 10208 6236 10260
rect 8116 10208 8168 10260
rect 9680 10208 9732 10260
rect 10508 10251 10560 10260
rect 6368 10183 6420 10192
rect 2044 10072 2096 10124
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 6368 10149 6377 10183
rect 6377 10149 6411 10183
rect 6411 10149 6420 10183
rect 6368 10140 6420 10149
rect 6644 10140 6696 10192
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 12256 10208 12308 10260
rect 13084 10251 13136 10260
rect 13084 10217 13093 10251
rect 13093 10217 13127 10251
rect 13127 10217 13136 10251
rect 13084 10208 13136 10217
rect 14188 10208 14240 10260
rect 15844 10208 15896 10260
rect 16396 10251 16448 10260
rect 16396 10217 16405 10251
rect 16405 10217 16439 10251
rect 16439 10217 16448 10251
rect 16396 10208 16448 10217
rect 17316 10208 17368 10260
rect 17960 10251 18012 10260
rect 17960 10217 17969 10251
rect 17969 10217 18003 10251
rect 18003 10217 18012 10251
rect 17960 10208 18012 10217
rect 18604 10208 18656 10260
rect 19248 10208 19300 10260
rect 21916 10208 21968 10260
rect 12624 10140 12676 10192
rect 17776 10140 17828 10192
rect 7012 10072 7064 10124
rect 8300 10072 8352 10124
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 10416 10072 10468 10124
rect 3240 9936 3292 9988
rect 3424 9979 3476 9988
rect 3424 9945 3433 9979
rect 3433 9945 3467 9979
rect 3467 9945 3476 9979
rect 3424 9936 3476 9945
rect 3608 9936 3660 9988
rect 2136 9911 2188 9920
rect 2136 9877 2145 9911
rect 2145 9877 2179 9911
rect 2179 9877 2188 9911
rect 2136 9868 2188 9877
rect 3792 9868 3844 9920
rect 5264 9868 5316 9920
rect 7012 9936 7064 9988
rect 8208 9936 8260 9988
rect 10232 10004 10284 10056
rect 11244 10072 11296 10124
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 12808 10004 12860 10056
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 16856 10072 16908 10124
rect 17040 10072 17092 10124
rect 8484 9868 8536 9920
rect 8668 9868 8720 9920
rect 9680 9868 9732 9920
rect 10600 9936 10652 9988
rect 14556 9868 14608 9920
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 17684 10004 17736 10056
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 19524 10004 19576 10056
rect 20444 10004 20496 10056
rect 23756 10004 23808 10056
rect 25412 10047 25464 10056
rect 25412 10013 25421 10047
rect 25421 10013 25455 10047
rect 25455 10013 25464 10047
rect 25412 10004 25464 10013
rect 30104 10004 30156 10056
rect 22744 9936 22796 9988
rect 25596 9936 25648 9988
rect 38016 9868 38068 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4528 9664 4580 9716
rect 4712 9664 4764 9716
rect 8300 9707 8352 9716
rect 2780 9639 2832 9648
rect 2780 9605 2789 9639
rect 2789 9605 2823 9639
rect 2823 9605 2832 9639
rect 2780 9596 2832 9605
rect 3424 9596 3476 9648
rect 6736 9596 6788 9648
rect 7104 9596 7156 9648
rect 7288 9639 7340 9648
rect 7288 9605 7297 9639
rect 7297 9605 7331 9639
rect 7331 9605 7340 9639
rect 7288 9596 7340 9605
rect 2044 9528 2096 9580
rect 5264 9528 5316 9580
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 7472 9528 7524 9580
rect 8300 9673 8309 9707
rect 8309 9673 8343 9707
rect 8343 9673 8352 9707
rect 8300 9664 8352 9673
rect 8392 9664 8444 9716
rect 11244 9664 11296 9716
rect 12532 9664 12584 9716
rect 14924 9664 14976 9716
rect 16856 9707 16908 9716
rect 16856 9673 16865 9707
rect 16865 9673 16899 9707
rect 16899 9673 16908 9707
rect 16856 9664 16908 9673
rect 17408 9664 17460 9716
rect 8116 9596 8168 9648
rect 10600 9639 10652 9648
rect 10600 9605 10609 9639
rect 10609 9605 10643 9639
rect 10643 9605 10652 9639
rect 10600 9596 10652 9605
rect 11152 9639 11204 9648
rect 11152 9605 11161 9639
rect 11161 9605 11195 9639
rect 11195 9605 11204 9639
rect 11152 9596 11204 9605
rect 11980 9596 12032 9648
rect 12072 9596 12124 9648
rect 9680 9528 9732 9580
rect 10232 9528 10284 9580
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 13820 9596 13872 9648
rect 13912 9596 13964 9648
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 14832 9528 14884 9580
rect 16488 9596 16540 9648
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 15936 9528 15988 9580
rect 17684 9528 17736 9580
rect 38108 9528 38160 9580
rect 6184 9460 6236 9512
rect 8760 9460 8812 9512
rect 10692 9460 10744 9512
rect 1676 9324 1728 9376
rect 7564 9392 7616 9444
rect 13360 9392 13412 9444
rect 15568 9392 15620 9444
rect 7840 9324 7892 9376
rect 8208 9324 8260 9376
rect 13544 9324 13596 9376
rect 17592 9324 17644 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 3976 9120 4028 9172
rect 5080 9163 5132 9172
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 7932 9120 7984 9172
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 9772 9163 9824 9172
rect 9772 9129 9781 9163
rect 9781 9129 9815 9163
rect 9815 9129 9824 9163
rect 9772 9120 9824 9129
rect 11612 9120 11664 9172
rect 11796 9120 11848 9172
rect 12716 9120 12768 9172
rect 12900 9120 12952 9172
rect 14648 9120 14700 9172
rect 15660 9163 15712 9172
rect 15660 9129 15669 9163
rect 15669 9129 15703 9163
rect 15703 9129 15712 9163
rect 15660 9120 15712 9129
rect 5356 9052 5408 9104
rect 2136 8984 2188 9036
rect 4620 8984 4672 9036
rect 5080 8984 5132 9036
rect 6000 8984 6052 9036
rect 6184 8984 6236 9036
rect 10140 9052 10192 9104
rect 8300 8984 8352 9036
rect 8484 8984 8536 9036
rect 4160 8916 4212 8968
rect 5448 8916 5500 8968
rect 1768 8848 1820 8900
rect 5540 8848 5592 8900
rect 4068 8780 4120 8832
rect 5632 8780 5684 8832
rect 7288 8848 7340 8900
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 10968 8916 11020 8968
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 11520 8916 11572 8968
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 14188 8984 14240 9036
rect 15016 9027 15068 9036
rect 15016 8993 15025 9027
rect 15025 8993 15059 9027
rect 15059 8993 15068 9027
rect 15016 8984 15068 8993
rect 16488 8959 16540 8968
rect 7564 8848 7616 8900
rect 16488 8925 16497 8959
rect 16497 8925 16531 8959
rect 16531 8925 16540 8959
rect 16488 8916 16540 8925
rect 18236 8916 18288 8968
rect 23020 8916 23072 8968
rect 30840 8959 30892 8968
rect 30840 8925 30849 8959
rect 30849 8925 30883 8959
rect 30883 8925 30892 8959
rect 30840 8916 30892 8925
rect 38016 8959 38068 8968
rect 38016 8925 38025 8959
rect 38025 8925 38059 8959
rect 38059 8925 38068 8959
rect 38016 8916 38068 8925
rect 8852 8780 8904 8832
rect 10324 8823 10376 8832
rect 10324 8789 10333 8823
rect 10333 8789 10367 8823
rect 10367 8789 10376 8823
rect 10324 8780 10376 8789
rect 10416 8780 10468 8832
rect 13360 8780 13412 8832
rect 20352 8848 20404 8900
rect 15476 8780 15528 8832
rect 20168 8780 20220 8832
rect 25504 8780 25556 8832
rect 33048 8780 33100 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 5632 8576 5684 8628
rect 6828 8576 6880 8628
rect 7288 8576 7340 8628
rect 1952 8551 2004 8560
rect 1952 8517 1961 8551
rect 1961 8517 1995 8551
rect 1995 8517 2004 8551
rect 1952 8508 2004 8517
rect 3700 8508 3752 8560
rect 3056 8440 3108 8492
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6368 8440 6420 8492
rect 7288 8440 7340 8492
rect 7472 8440 7524 8492
rect 8024 8576 8076 8628
rect 9220 8576 9272 8628
rect 10048 8576 10100 8628
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 11704 8576 11756 8628
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 15108 8576 15160 8628
rect 15200 8576 15252 8628
rect 8116 8508 8168 8560
rect 2044 8372 2096 8424
rect 3332 8372 3384 8424
rect 5632 8372 5684 8424
rect 8208 8372 8260 8424
rect 1584 8304 1636 8356
rect 6920 8304 6972 8356
rect 9864 8440 9916 8492
rect 10968 8440 11020 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 11888 8508 11940 8560
rect 14556 8440 14608 8492
rect 16488 8508 16540 8560
rect 15476 8483 15528 8492
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15476 8440 15528 8449
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 16304 8440 16356 8492
rect 16764 8304 16816 8356
rect 16856 8304 16908 8356
rect 1952 8236 2004 8288
rect 4620 8236 4672 8288
rect 7380 8236 7432 8288
rect 11244 8236 11296 8288
rect 11612 8236 11664 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1952 8032 2004 8084
rect 3424 8007 3476 8016
rect 3424 7973 3433 8007
rect 3433 7973 3467 8007
rect 3467 7973 3476 8007
rect 3424 7964 3476 7973
rect 2044 7896 2096 7948
rect 4344 8032 4396 8084
rect 4712 7964 4764 8016
rect 7380 8032 7432 8084
rect 10600 8032 10652 8084
rect 4252 7896 4304 7948
rect 5080 7939 5132 7948
rect 5080 7905 5089 7939
rect 5089 7905 5123 7939
rect 5123 7905 5132 7939
rect 5080 7896 5132 7905
rect 9772 7964 9824 8016
rect 5816 7896 5868 7948
rect 6644 7896 6696 7948
rect 7288 7871 7340 7880
rect 1492 7760 1544 7812
rect 2964 7760 3016 7812
rect 4436 7803 4488 7812
rect 4436 7769 4445 7803
rect 4445 7769 4479 7803
rect 4479 7769 4488 7803
rect 4436 7760 4488 7769
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 11612 7871 11664 7880
rect 5264 7760 5316 7812
rect 5816 7760 5868 7812
rect 11152 7760 11204 7812
rect 4712 7692 4764 7744
rect 4988 7692 5040 7744
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 33048 7828 33100 7880
rect 14740 7760 14792 7812
rect 38016 7692 38068 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1584 7488 1636 7540
rect 3148 7488 3200 7540
rect 5172 7488 5224 7540
rect 5448 7488 5500 7540
rect 6644 7531 6696 7540
rect 1952 7352 2004 7404
rect 4160 7420 4212 7472
rect 4988 7420 5040 7472
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 9220 7531 9272 7540
rect 9220 7497 9229 7531
rect 9229 7497 9263 7531
rect 9263 7497 9272 7531
rect 9220 7488 9272 7497
rect 24400 7488 24452 7540
rect 38108 7531 38160 7540
rect 38108 7497 38117 7531
rect 38117 7497 38151 7531
rect 38151 7497 38160 7531
rect 38108 7488 38160 7497
rect 6644 7352 6696 7404
rect 29736 7352 29788 7404
rect 34336 7352 34388 7404
rect 38292 7395 38344 7404
rect 38292 7361 38301 7395
rect 38301 7361 38335 7395
rect 38335 7361 38344 7395
rect 38292 7352 38344 7361
rect 3792 7284 3844 7336
rect 4620 7284 4672 7336
rect 5080 7284 5132 7336
rect 4252 7216 4304 7268
rect 12072 7216 12124 7268
rect 22652 7216 22704 7268
rect 4620 7148 4672 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2228 6944 2280 6996
rect 2688 6851 2740 6860
rect 2688 6817 2697 6851
rect 2697 6817 2731 6851
rect 2731 6817 2740 6851
rect 2688 6808 2740 6817
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 2872 6740 2924 6792
rect 3700 6808 3752 6860
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 5724 6808 5776 6860
rect 6000 6876 6052 6928
rect 7196 6876 7248 6928
rect 9588 6808 9640 6860
rect 10784 6808 10836 6860
rect 14464 6808 14516 6860
rect 21548 6808 21600 6860
rect 4712 6740 4764 6792
rect 3792 6672 3844 6724
rect 5448 6740 5500 6792
rect 14280 6783 14332 6792
rect 3332 6604 3384 6656
rect 4712 6604 4764 6656
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 23388 6740 23440 6792
rect 8760 6672 8812 6724
rect 9312 6715 9364 6724
rect 9312 6681 9321 6715
rect 9321 6681 9355 6715
rect 9355 6681 9364 6715
rect 9312 6672 9364 6681
rect 20812 6672 20864 6724
rect 30564 6740 30616 6792
rect 33048 6740 33100 6792
rect 35624 6740 35676 6792
rect 12808 6604 12860 6656
rect 20076 6604 20128 6656
rect 24492 6604 24544 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2596 6400 2648 6452
rect 2964 6400 3016 6452
rect 3516 6400 3568 6452
rect 3884 6400 3936 6452
rect 4804 6400 4856 6452
rect 8760 6400 8812 6452
rect 9312 6400 9364 6452
rect 2964 6264 3016 6316
rect 3332 6264 3384 6316
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4160 6264 4212 6273
rect 6368 6332 6420 6384
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 4804 6196 4856 6248
rect 8576 6264 8628 6316
rect 13452 6264 13504 6316
rect 30288 6264 30340 6316
rect 11060 6196 11112 6248
rect 11704 6128 11756 6180
rect 6368 6060 6420 6112
rect 16672 6060 16724 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3056 5856 3108 5908
rect 4896 5856 4948 5908
rect 5080 5856 5132 5908
rect 6736 5856 6788 5908
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 15752 5856 15804 5908
rect 3240 5788 3292 5840
rect 9588 5788 9640 5840
rect 6736 5720 6788 5772
rect 2964 5652 3016 5704
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 4068 5652 4120 5704
rect 5908 5652 5960 5704
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 32864 5695 32916 5704
rect 32864 5661 32873 5695
rect 32873 5661 32907 5695
rect 32907 5661 32916 5695
rect 32864 5652 32916 5661
rect 36820 5695 36872 5704
rect 36820 5661 36829 5695
rect 36829 5661 36863 5695
rect 36863 5661 36872 5695
rect 36820 5652 36872 5661
rect 38016 5695 38068 5704
rect 38016 5661 38025 5695
rect 38025 5661 38059 5695
rect 38059 5661 38068 5695
rect 38016 5652 38068 5661
rect 6000 5584 6052 5636
rect 6368 5627 6420 5636
rect 6368 5593 6377 5627
rect 6377 5593 6411 5627
rect 6411 5593 6420 5627
rect 6368 5584 6420 5593
rect 7564 5584 7616 5636
rect 5632 5559 5684 5568
rect 5632 5525 5641 5559
rect 5641 5525 5675 5559
rect 5675 5525 5684 5559
rect 5632 5516 5684 5525
rect 34428 5516 34480 5568
rect 37464 5516 37516 5568
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4620 5312 4672 5364
rect 4988 5355 5040 5364
rect 4988 5321 4997 5355
rect 4997 5321 5031 5355
rect 5031 5321 5040 5355
rect 4988 5312 5040 5321
rect 1676 5015 1728 5024
rect 1676 4981 1685 5015
rect 1685 4981 1719 5015
rect 1719 4981 1728 5015
rect 1676 4972 1728 4981
rect 2872 5176 2924 5228
rect 4344 5176 4396 5228
rect 8484 5244 8536 5296
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 5356 5176 5408 5228
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 20168 5219 20220 5228
rect 20168 5185 20177 5219
rect 20177 5185 20211 5219
rect 20211 5185 20220 5219
rect 20168 5176 20220 5185
rect 25504 5219 25556 5228
rect 25504 5185 25513 5219
rect 25513 5185 25547 5219
rect 25547 5185 25556 5219
rect 25504 5176 25556 5185
rect 25596 5176 25648 5228
rect 37464 5219 37516 5228
rect 37464 5185 37473 5219
rect 37473 5185 37507 5219
rect 37507 5185 37516 5219
rect 37464 5176 37516 5185
rect 7012 5108 7064 5160
rect 6828 5040 6880 5092
rect 27804 5040 27856 5092
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 4344 4972 4396 5024
rect 7564 4972 7616 5024
rect 20076 4972 20128 5024
rect 23296 4972 23348 5024
rect 30012 4972 30064 5024
rect 38016 4972 38068 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1768 4768 1820 4820
rect 3608 4768 3660 4820
rect 6460 4768 6512 4820
rect 5816 4700 5868 4752
rect 3424 4632 3476 4684
rect 6552 4632 6604 4684
rect 7656 4632 7708 4684
rect 1676 4564 1728 4616
rect 3792 4564 3844 4616
rect 2964 4496 3016 4548
rect 5632 4564 5684 4616
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 12624 4564 12676 4616
rect 16764 4564 16816 4616
rect 4620 4471 4672 4480
rect 4620 4437 4629 4471
rect 4629 4437 4663 4471
rect 4663 4437 4672 4471
rect 4620 4428 4672 4437
rect 18604 4428 18656 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 2228 4088 2280 4140
rect 4896 4088 4948 4140
rect 17316 4088 17368 4140
rect 1400 4020 1452 4072
rect 9220 4020 9272 4072
rect 3516 3995 3568 4004
rect 3516 3961 3525 3995
rect 3525 3961 3559 3995
rect 3559 3961 3568 3995
rect 3516 3952 3568 3961
rect 9588 3884 9640 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2412 3680 2464 3732
rect 4712 3680 4764 3732
rect 30748 3680 30800 3732
rect 7748 3612 7800 3664
rect 2964 3476 3016 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 38292 3519 38344 3528
rect 38292 3485 38301 3519
rect 38301 3485 38335 3519
rect 38335 3485 38344 3519
rect 38292 3476 38344 3485
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2780 3068 2832 3120
rect 5264 3136 5316 3188
rect 35624 3136 35676 3188
rect 5540 3068 5592 3120
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 1308 2932 1360 2984
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 37280 3000 37332 3052
rect 38016 3043 38068 3052
rect 38016 3009 38025 3043
rect 38025 3009 38059 3043
rect 38059 3009 38068 3043
rect 38016 3000 38068 3009
rect 6920 2864 6972 2916
rect 6644 2796 6696 2848
rect 9404 2839 9456 2848
rect 9404 2805 9413 2839
rect 9413 2805 9447 2839
rect 9447 2805 9456 2839
rect 9404 2796 9456 2805
rect 38200 2839 38252 2848
rect 38200 2805 38209 2839
rect 38209 2805 38243 2839
rect 38243 2805 38252 2839
rect 38200 2796 38252 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3240 2592 3292 2644
rect 4804 2635 4856 2644
rect 4804 2601 4813 2635
rect 4813 2601 4847 2635
rect 4847 2601 4856 2635
rect 4804 2592 4856 2601
rect 7288 2592 7340 2644
rect 9864 2592 9916 2644
rect 10048 2592 10100 2644
rect 14280 2592 14332 2644
rect 15476 2592 15528 2644
rect 16948 2592 17000 2644
rect 20444 2592 20496 2644
rect 23388 2592 23440 2644
rect 25412 2592 25464 2644
rect 29736 2635 29788 2644
rect 29736 2601 29745 2635
rect 29745 2601 29779 2635
rect 29779 2601 29788 2635
rect 29736 2592 29788 2601
rect 30288 2592 30340 2644
rect 34336 2592 34388 2644
rect 4620 2524 4672 2576
rect 30564 2524 30616 2576
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 34428 2456 34480 2508
rect 2596 2388 2648 2440
rect 4528 2388 4580 2440
rect 5816 2388 5868 2440
rect 7748 2388 7800 2440
rect 9404 2431 9456 2440
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 10324 2388 10376 2440
rect 12256 2388 12308 2440
rect 13544 2388 13596 2440
rect 15476 2388 15528 2440
rect 16764 2388 16816 2440
rect 18604 2431 18656 2440
rect 18604 2397 18613 2431
rect 18613 2397 18647 2431
rect 18647 2397 18656 2431
rect 18604 2388 18656 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 21272 2388 21324 2440
rect 23296 2431 23348 2440
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 24492 2388 24544 2440
rect 26424 2388 26476 2440
rect 27804 2431 27856 2440
rect 27804 2397 27813 2431
rect 27813 2397 27847 2431
rect 27847 2397 27856 2431
rect 27804 2388 27856 2397
rect 29000 2388 29052 2440
rect 30012 2388 30064 2440
rect 32220 2388 32272 2440
rect 34152 2388 34204 2440
rect 35440 2388 35492 2440
rect 38660 2320 38712 2372
rect 20 2252 72 2304
rect 9036 2252 9088 2304
rect 18696 2252 18748 2304
rect 19984 2252 20036 2304
rect 23204 2252 23256 2304
rect 27712 2252 27764 2304
rect 30932 2252 30984 2304
rect 33048 2252 33100 2304
rect 37372 2252 37424 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 2778 39536 2834 39545
rect 2778 39471 2834 39480
rect 676 36922 704 39200
rect 1964 37262 1992 39200
rect 1860 37256 1912 37262
rect 1860 37198 1912 37204
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 1872 36922 1900 37198
rect 2792 37194 2820 39471
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 16224 39222 16528 39250
rect 2962 37496 3018 37505
rect 2962 37431 3018 37440
rect 2976 37262 3004 37431
rect 2964 37256 3016 37262
rect 2964 37198 3016 37204
rect 2780 37188 2832 37194
rect 2780 37130 2832 37136
rect 3896 37126 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4252 37256 4304 37262
rect 4252 37198 4304 37204
rect 3148 37120 3200 37126
rect 3148 37062 3200 37068
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 664 36916 716 36922
rect 664 36858 716 36864
rect 1860 36916 1912 36922
rect 1860 36858 1912 36864
rect 1584 36168 1636 36174
rect 1582 36136 1584 36145
rect 1636 36136 1638 36145
rect 1582 36071 1638 36080
rect 1676 34400 1728 34406
rect 1676 34342 1728 34348
rect 1688 34105 1716 34342
rect 1674 34096 1730 34105
rect 1674 34031 1730 34040
rect 1584 32904 1636 32910
rect 1584 32846 1636 32852
rect 1596 32745 1624 32846
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 3160 32434 3188 37062
rect 3976 36916 4028 36922
rect 3976 36858 4028 36864
rect 3988 35290 4016 36858
rect 4068 36780 4120 36786
rect 4068 36722 4120 36728
rect 3976 35284 4028 35290
rect 3976 35226 4028 35232
rect 4080 34746 4108 36722
rect 4264 36689 4292 37198
rect 5184 37126 5212 39200
rect 7116 37262 7144 39200
rect 8404 37262 8432 39200
rect 10336 37262 10364 39200
rect 11624 37262 11652 39200
rect 12912 37262 12940 39200
rect 5540 37256 5592 37262
rect 5540 37198 5592 37204
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 10324 37256 10376 37262
rect 10324 37198 10376 37204
rect 11612 37256 11664 37262
rect 11612 37198 11664 37204
rect 12900 37256 12952 37262
rect 12900 37198 12952 37204
rect 5172 37120 5224 37126
rect 5172 37062 5224 37068
rect 4250 36680 4306 36689
rect 4250 36615 4306 36624
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 5552 35834 5580 37198
rect 6552 37188 6604 37194
rect 6552 37130 6604 37136
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5908 35692 5960 35698
rect 5908 35634 5960 35640
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 34740 4120 34746
rect 4068 34682 4120 34688
rect 3976 34604 4028 34610
rect 3976 34546 4028 34552
rect 3148 32428 3200 32434
rect 3148 32370 3200 32376
rect 3988 30938 4016 34546
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4620 32768 4672 32774
rect 4620 32710 4672 32716
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3976 30932 4028 30938
rect 3976 30874 4028 30880
rect 1584 30728 1636 30734
rect 1582 30696 1584 30705
rect 4068 30728 4120 30734
rect 1636 30696 1638 30705
rect 4068 30670 4120 30676
rect 1582 30631 1638 30640
rect 2964 30252 3016 30258
rect 2964 30194 3016 30200
rect 2228 30184 2280 30190
rect 2228 30126 2280 30132
rect 1676 29504 1728 29510
rect 1676 29446 1728 29452
rect 1688 29345 1716 29446
rect 1674 29336 1730 29345
rect 1674 29271 1730 29280
rect 1584 29164 1636 29170
rect 1584 29106 1636 29112
rect 1596 27985 1624 29106
rect 2240 28082 2268 30126
rect 2596 29708 2648 29714
rect 2596 29650 2648 29656
rect 2320 29096 2372 29102
rect 2320 29038 2372 29044
rect 2228 28076 2280 28082
rect 2228 28018 2280 28024
rect 1582 27976 1638 27985
rect 1582 27911 1638 27920
rect 2044 27872 2096 27878
rect 2044 27814 2096 27820
rect 1768 27328 1820 27334
rect 1768 27270 1820 27276
rect 20 26988 72 26994
rect 20 26930 72 26936
rect 32 17785 60 26930
rect 1582 25936 1638 25945
rect 1582 25871 1584 25880
rect 1636 25871 1638 25880
rect 1584 25842 1636 25848
rect 1308 25764 1360 25770
rect 1308 25706 1360 25712
rect 18 17776 74 17785
rect 18 17711 74 17720
rect 1320 14006 1348 25706
rect 1676 24608 1728 24614
rect 1674 24576 1676 24585
rect 1728 24576 1730 24585
rect 1674 24511 1730 24520
rect 1492 24200 1544 24206
rect 1492 24142 1544 24148
rect 1400 21888 1452 21894
rect 1400 21830 1452 21836
rect 1412 21078 1440 21830
rect 1400 21072 1452 21078
rect 1400 21014 1452 21020
rect 1308 14000 1360 14006
rect 1308 13942 1360 13948
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1412 4078 1440 13126
rect 1504 12866 1532 24142
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 1596 22545 1624 22578
rect 1582 22536 1638 22545
rect 1582 22471 1638 22480
rect 1674 21176 1730 21185
rect 1674 21111 1730 21120
rect 1688 20602 1716 21111
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1688 16794 1716 18158
rect 1780 17610 1808 27270
rect 1860 26784 1912 26790
rect 1860 26726 1912 26732
rect 1872 26353 1900 26726
rect 1858 26344 1914 26353
rect 1858 26279 1914 26288
rect 1952 26308 2004 26314
rect 1952 26250 2004 26256
rect 1860 25696 1912 25702
rect 1860 25638 1912 25644
rect 1872 25294 1900 25638
rect 1860 25288 1912 25294
rect 1860 25230 1912 25236
rect 1860 24676 1912 24682
rect 1860 24618 1912 24624
rect 1872 23866 1900 24618
rect 1860 23860 1912 23866
rect 1860 23802 1912 23808
rect 1860 23316 1912 23322
rect 1860 23258 1912 23264
rect 1872 22778 1900 23258
rect 1860 22772 1912 22778
rect 1860 22714 1912 22720
rect 1860 21888 1912 21894
rect 1860 21830 1912 21836
rect 1768 17604 1820 17610
rect 1768 17546 1820 17552
rect 1872 17490 1900 21830
rect 1964 18834 1992 26250
rect 2056 21622 2084 27814
rect 2240 27470 2268 28018
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 2240 25906 2268 27406
rect 2332 27402 2360 29038
rect 2504 28484 2556 28490
rect 2504 28426 2556 28432
rect 2320 27396 2372 27402
rect 2320 27338 2372 27344
rect 2332 26382 2360 27338
rect 2516 26994 2544 28426
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2504 26784 2556 26790
rect 2504 26726 2556 26732
rect 2320 26376 2372 26382
rect 2320 26318 2372 26324
rect 2228 25900 2280 25906
rect 2228 25842 2280 25848
rect 2136 25152 2188 25158
rect 2136 25094 2188 25100
rect 2148 24206 2176 25094
rect 2240 24206 2268 25842
rect 2332 24290 2360 26318
rect 2412 25288 2464 25294
rect 2412 25230 2464 25236
rect 2424 24818 2452 25230
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2424 24410 2452 24754
rect 2412 24404 2464 24410
rect 2412 24346 2464 24352
rect 2332 24262 2452 24290
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2228 23180 2280 23186
rect 2228 23122 2280 23128
rect 2136 23044 2188 23050
rect 2136 22986 2188 22992
rect 2148 22778 2176 22986
rect 2136 22772 2188 22778
rect 2136 22714 2188 22720
rect 2240 22642 2268 23122
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 2136 22092 2188 22098
rect 2240 22080 2268 22578
rect 2320 22432 2372 22438
rect 2320 22374 2372 22380
rect 2188 22052 2268 22080
rect 2136 22034 2188 22040
rect 2044 21616 2096 21622
rect 2044 21558 2096 21564
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 2056 19922 2084 21082
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2148 19802 2176 21422
rect 2240 21418 2268 22052
rect 2228 21412 2280 21418
rect 2228 21354 2280 21360
rect 2240 21146 2268 21354
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 2056 19774 2176 19802
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 2056 18222 2084 19774
rect 2332 19666 2360 22374
rect 2148 19638 2360 19666
rect 2044 18216 2096 18222
rect 1950 18184 2006 18193
rect 2044 18158 2096 18164
rect 1950 18119 2006 18128
rect 1780 17462 1900 17490
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1582 16416 1638 16425
rect 1582 16351 1638 16360
rect 1596 16250 1624 16351
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1688 14482 1716 16730
rect 1780 15026 1808 17462
rect 1964 16114 1992 18119
rect 2148 17270 2176 19638
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 2136 17264 2188 17270
rect 2136 17206 2188 17212
rect 2042 16280 2098 16289
rect 2042 16215 2098 16224
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 2056 15162 2084 16215
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1780 14906 1808 14962
rect 1780 14878 1992 14906
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1688 14074 1716 14418
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 13394 1624 13806
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1504 12838 1624 12866
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1504 10266 1532 12718
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1504 7818 1532 10202
rect 1596 8362 1624 12838
rect 1688 11558 1716 13670
rect 1768 13252 1820 13258
rect 1768 13194 1820 13200
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11354 1716 11494
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1780 11234 1808 13194
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1688 11206 1808 11234
rect 1688 9382 1716 11206
rect 1872 9674 1900 12038
rect 1964 11098 1992 14878
rect 2240 13530 2268 19450
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2332 15910 2360 19314
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2056 11234 2084 11630
rect 2056 11206 2176 11234
rect 1964 11070 2084 11098
rect 1950 10976 2006 10985
rect 1950 10911 2006 10920
rect 1964 10742 1992 10911
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 2056 10130 2084 11070
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1872 9646 1992 9674
rect 1768 9512 1820 9518
rect 1766 9480 1768 9489
rect 1820 9480 1822 9489
rect 1766 9415 1822 9424
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 9178 1716 9318
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 1596 7546 1624 8191
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4865 1716 4966
rect 1674 4856 1730 4865
rect 1780 4826 1808 8842
rect 1964 8673 1992 9646
rect 2056 9586 2084 10066
rect 2148 9926 2176 11206
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2148 9042 2176 9862
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 1950 8664 2006 8673
rect 1950 8599 2006 8608
rect 1964 8566 1992 8599
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 2044 8424 2096 8430
rect 2148 8378 2176 8978
rect 2096 8372 2176 8378
rect 2044 8366 2176 8372
rect 2056 8350 2176 8366
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1964 8090 1992 8230
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1964 7410 1992 8026
rect 2148 7970 2176 8350
rect 2056 7954 2176 7970
rect 2044 7948 2176 7954
rect 2096 7942 2176 7948
rect 2044 7890 2096 7896
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1964 6798 1992 7346
rect 2240 7002 2268 12786
rect 2332 11830 2360 14962
rect 2424 11898 2452 24262
rect 2516 22094 2544 26726
rect 2608 23730 2636 29650
rect 2976 29646 3004 30194
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 2976 29102 3004 29582
rect 3608 29572 3660 29578
rect 3608 29514 3660 29520
rect 2964 29096 3016 29102
rect 2964 29038 3016 29044
rect 2976 28558 3004 29038
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 2596 23724 2648 23730
rect 2596 23666 2648 23672
rect 2596 23520 2648 23526
rect 2596 23462 2648 23468
rect 2608 22438 2636 23462
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2516 22066 2636 22094
rect 2608 21962 2636 22066
rect 2596 21956 2648 21962
rect 2596 21898 2648 21904
rect 2700 19786 2728 27814
rect 2872 27328 2924 27334
rect 2872 27270 2924 27276
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2792 19825 2820 23598
rect 2884 20466 2912 27270
rect 2976 26382 3004 28494
rect 3516 27328 3568 27334
rect 3516 27270 3568 27276
rect 3148 26784 3200 26790
rect 3148 26726 3200 26732
rect 2964 26376 3016 26382
rect 2964 26318 3016 26324
rect 2976 24342 3004 26318
rect 3056 25220 3108 25226
rect 3056 25162 3108 25168
rect 3068 24818 3096 25162
rect 3056 24812 3108 24818
rect 3056 24754 3108 24760
rect 2964 24336 3016 24342
rect 2964 24278 3016 24284
rect 2976 23730 3004 24278
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 3054 23624 3110 23633
rect 3054 23559 3056 23568
rect 3108 23559 3110 23568
rect 3056 23530 3108 23536
rect 2964 22228 3016 22234
rect 2964 22170 3016 22176
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2778 19816 2834 19825
rect 2688 19780 2740 19786
rect 2778 19751 2834 19760
rect 2688 19722 2740 19728
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2884 15570 2912 15982
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2792 14618 2820 14758
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2778 14512 2834 14521
rect 2778 14447 2834 14456
rect 2792 12434 2820 14447
rect 2884 13394 2912 15506
rect 2976 14414 3004 22170
rect 3160 20534 3188 26726
rect 3240 25696 3292 25702
rect 3240 25638 3292 25644
rect 3252 24818 3280 25638
rect 3240 24812 3292 24818
rect 3240 24754 3292 24760
rect 3332 24064 3384 24070
rect 3332 24006 3384 24012
rect 3344 23497 3372 24006
rect 3330 23488 3386 23497
rect 3330 23423 3386 23432
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3240 21616 3292 21622
rect 3240 21558 3292 21564
rect 3148 20528 3200 20534
rect 3148 20470 3200 20476
rect 3054 18728 3110 18737
rect 3054 18663 3056 18672
rect 3108 18663 3110 18672
rect 3056 18634 3108 18640
rect 3068 14550 3096 18634
rect 3252 18426 3280 21558
rect 3344 19378 3372 22918
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 3436 20398 3464 22714
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3436 20058 3464 20198
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 3148 17264 3200 17270
rect 3148 17206 3200 17212
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2884 12782 2912 13330
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2792 12406 2912 12434
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2320 11824 2372 11830
rect 2318 11792 2320 11801
rect 2372 11792 2374 11801
rect 2318 11727 2374 11736
rect 2686 11248 2742 11257
rect 2792 11218 2820 12242
rect 2686 11183 2742 11192
rect 2780 11212 2832 11218
rect 2700 11082 2728 11183
rect 2780 11154 2832 11160
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2792 10810 2820 11154
rect 2884 10810 2912 12406
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3068 11354 3096 12106
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1674 4791 1730 4800
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1688 4146 1716 4558
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 2240 3058 2268 4082
rect 2424 3738 2452 10406
rect 2792 9654 2820 10746
rect 2870 10568 2926 10577
rect 2870 10503 2926 10512
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2884 7426 2912 10503
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2608 7398 2912 7426
rect 2608 6458 2636 7398
rect 2686 6896 2742 6905
rect 2686 6831 2688 6840
rect 2740 6831 2742 6840
rect 2688 6802 2740 6808
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2778 6216 2834 6225
rect 2778 6151 2834 6160
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2792 3126 2820 6151
rect 2884 5234 2912 6734
rect 2976 6458 3004 7754
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2976 5710 3004 6258
rect 3068 5914 3096 8434
rect 3160 7546 3188 17206
rect 3344 17134 3372 19314
rect 3436 18170 3464 19654
rect 3528 18358 3556 27270
rect 3620 27130 3648 29514
rect 3884 29028 3936 29034
rect 3884 28970 3936 28976
rect 3608 27124 3660 27130
rect 3608 27066 3660 27072
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 3804 26042 3832 26930
rect 3792 26036 3844 26042
rect 3792 25978 3844 25984
rect 3700 25356 3752 25362
rect 3700 25298 3752 25304
rect 3608 25152 3660 25158
rect 3608 25094 3660 25100
rect 3620 24750 3648 25094
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3608 22500 3660 22506
rect 3608 22442 3660 22448
rect 3516 18352 3568 18358
rect 3516 18294 3568 18300
rect 3436 18142 3556 18170
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3436 17678 3464 18022
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3252 15706 3280 15982
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3252 9994 3280 14282
rect 3344 12918 3372 16390
rect 3436 14521 3464 17478
rect 3422 14512 3478 14521
rect 3422 14447 3478 14456
rect 3528 14006 3556 18142
rect 3620 16522 3648 22442
rect 3712 21554 3740 25298
rect 3896 23866 3924 28970
rect 4080 28762 4108 30670
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29170 4660 32710
rect 5920 30938 5948 35634
rect 6184 32224 6236 32230
rect 6184 32166 6236 32172
rect 5908 30932 5960 30938
rect 5908 30874 5960 30880
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 5000 29170 5028 29582
rect 4620 29164 4672 29170
rect 4620 29106 4672 29112
rect 4988 29164 5040 29170
rect 4988 29106 5040 29112
rect 5080 29096 5132 29102
rect 5078 29064 5080 29073
rect 5132 29064 5134 29073
rect 5078 28999 5134 29008
rect 5356 29028 5408 29034
rect 5356 28970 5408 28976
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 4896 28552 4948 28558
rect 4896 28494 4948 28500
rect 4068 28076 4120 28082
rect 4068 28018 4120 28024
rect 3976 27872 4028 27878
rect 3976 27814 4028 27820
rect 3884 23860 3936 23866
rect 3884 23802 3936 23808
rect 3884 23724 3936 23730
rect 3884 23666 3936 23672
rect 3896 23118 3924 23666
rect 3884 23112 3936 23118
rect 3884 23054 3936 23060
rect 3792 22704 3844 22710
rect 3792 22646 3844 22652
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3804 20777 3832 22646
rect 3896 22030 3924 23054
rect 3988 22094 4016 27814
rect 4080 27470 4108 28018
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 4080 27062 4108 27406
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4066 26344 4122 26353
rect 4066 26279 4068 26288
rect 4120 26279 4122 26288
rect 4068 26250 4120 26256
rect 4344 26240 4396 26246
rect 4344 26182 4396 26188
rect 4356 25974 4384 26182
rect 4344 25968 4396 25974
rect 4344 25910 4396 25916
rect 4620 25696 4672 25702
rect 4620 25638 4672 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 4080 22234 4108 25434
rect 4632 24818 4660 25638
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4252 24404 4304 24410
rect 4252 24346 4304 24352
rect 4264 23730 4292 24346
rect 4724 24274 4752 26726
rect 4816 26586 4844 26930
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4816 25906 4844 26318
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4712 24268 4764 24274
rect 4712 24210 4764 24216
rect 4344 23792 4396 23798
rect 4342 23760 4344 23769
rect 4396 23760 4398 23769
rect 4252 23724 4304 23730
rect 4342 23695 4398 23704
rect 4712 23724 4764 23730
rect 4252 23666 4304 23672
rect 4712 23666 4764 23672
rect 4620 23656 4672 23662
rect 4620 23598 4672 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 22642 4660 23598
rect 4724 23118 4752 23666
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 22228 4120 22234
rect 4068 22170 4120 22176
rect 3988 22066 4108 22094
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 3790 20768 3846 20777
rect 3790 20703 3846 20712
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3988 19718 4016 20538
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3698 19544 3754 19553
rect 3698 19479 3754 19488
rect 3712 19378 3740 19479
rect 4080 19446 4108 22066
rect 4528 22092 4580 22098
rect 4528 22034 4580 22040
rect 4252 21956 4304 21962
rect 4252 21898 4304 21904
rect 4264 21690 4292 21898
rect 4252 21684 4304 21690
rect 4252 21626 4304 21632
rect 4540 21434 4568 22034
rect 4540 21418 4660 21434
rect 4540 21412 4672 21418
rect 4540 21406 4620 21412
rect 4620 21354 4672 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4160 21072 4212 21078
rect 4160 21014 4212 21020
rect 4172 20534 4200 21014
rect 4160 20528 4212 20534
rect 4160 20470 4212 20476
rect 4632 20398 4660 21354
rect 4724 21162 4752 22918
rect 4816 21962 4844 25842
rect 4908 24818 4936 28494
rect 4988 27872 5040 27878
rect 4988 27814 5040 27820
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4908 24410 4936 24754
rect 4896 24404 4948 24410
rect 4896 24346 4948 24352
rect 5000 24290 5028 27814
rect 5080 26784 5132 26790
rect 5080 26726 5132 26732
rect 4908 24262 5028 24290
rect 4804 21956 4856 21962
rect 4804 21898 4856 21904
rect 4724 21134 4844 21162
rect 4712 21072 4764 21078
rect 4712 21014 4764 21020
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 3884 19440 3936 19446
rect 3884 19382 3936 19388
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3712 17610 3740 19314
rect 3792 18080 3844 18086
rect 3792 18022 3844 18028
rect 3700 17604 3752 17610
rect 3700 17546 3752 17552
rect 3804 17542 3832 18022
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3896 17490 3924 19382
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 17678 4016 19246
rect 4172 19156 4200 19790
rect 4632 19786 4660 20334
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4080 19128 4200 19156
rect 4080 18952 4108 19128
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4080 18924 4200 18952
rect 4172 18086 4200 18924
rect 4632 18834 4660 19722
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4448 18426 4476 18702
rect 4436 18420 4488 18426
rect 4436 18362 4488 18368
rect 4724 18358 4752 21014
rect 4816 19718 4844 21134
rect 4908 21078 4936 24262
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 5000 23730 5028 24142
rect 4988 23724 5040 23730
rect 4988 23666 5040 23672
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 5000 23050 5028 23462
rect 4988 23044 5040 23050
rect 4988 22986 5040 22992
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 4896 21072 4948 21078
rect 4896 21014 4948 21020
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4908 19990 4936 20878
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4816 17746 4844 18770
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 4620 17604 4672 17610
rect 4620 17546 4672 17552
rect 4632 17513 4660 17546
rect 4618 17504 4674 17513
rect 3804 17270 3832 17478
rect 3896 17462 4016 17490
rect 3792 17264 3844 17270
rect 3792 17206 3844 17212
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3608 16516 3660 16522
rect 3608 16458 3660 16464
rect 3896 16250 3924 17070
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 3608 15564 3660 15570
rect 3608 15506 3660 15512
rect 3620 15026 3648 15506
rect 3884 15428 3936 15434
rect 3884 15370 3936 15376
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3712 14385 3740 15098
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3698 14376 3754 14385
rect 3698 14311 3754 14320
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3804 13682 3832 15030
rect 3620 13654 3832 13682
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3528 12306 3556 12582
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3620 11778 3648 13654
rect 3790 13560 3846 13569
rect 3790 13495 3846 13504
rect 3700 12912 3752 12918
rect 3700 12854 3752 12860
rect 3344 11750 3648 11778
rect 3240 9988 3292 9994
rect 3240 9930 3292 9936
rect 3238 9616 3294 9625
rect 3238 9551 3294 9560
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3252 5846 3280 9551
rect 3344 8430 3372 11750
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3436 9654 3464 9930
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3422 8120 3478 8129
rect 3422 8055 3478 8064
rect 3436 8022 3464 8055
rect 3424 8016 3476 8022
rect 3424 7958 3476 7964
rect 3332 6792 3384 6798
rect 3330 6760 3332 6769
rect 3384 6760 3386 6769
rect 3330 6695 3386 6704
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3344 6322 3372 6598
rect 3528 6458 3556 11290
rect 3620 9994 3648 11562
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3712 8650 3740 12854
rect 3804 11082 3832 13495
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3620 8622 3740 8650
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 2872 5228 2924 5234
rect 2924 5188 3004 5216
rect 2872 5170 2924 5176
rect 2976 4554 3004 5188
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2976 3534 3004 4490
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 32 800 60 2246
rect 1320 800 1348 2926
rect 3252 2650 3280 5646
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3436 4690 3464 4966
rect 3620 4826 3648 8622
rect 3700 8560 3752 8566
rect 3700 8502 3752 8508
rect 3712 6866 3740 8502
rect 3804 7342 3832 9862
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3804 6730 3832 7278
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3804 4622 3832 6666
rect 3896 6458 3924 15370
rect 3988 12434 4016 17462
rect 4618 17439 4674 17448
rect 4816 17202 4844 17682
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4080 16658 4108 16934
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4528 16516 4580 16522
rect 4528 16458 4580 16464
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 15366 4108 16390
rect 4540 16114 4568 16458
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4448 13870 4476 14554
rect 4632 14521 4660 16730
rect 4816 16658 4844 17138
rect 4908 16794 4936 17138
rect 5000 16969 5028 22578
rect 5092 17610 5120 26726
rect 5172 26240 5224 26246
rect 5172 26182 5224 26188
rect 5184 25294 5212 26182
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 5172 24812 5224 24818
rect 5172 24754 5224 24760
rect 5184 24274 5212 24754
rect 5172 24268 5224 24274
rect 5172 24210 5224 24216
rect 5172 24132 5224 24138
rect 5172 24074 5224 24080
rect 5184 23050 5212 24074
rect 5276 23866 5304 25094
rect 5368 24274 5396 28970
rect 5632 27328 5684 27334
rect 5632 27270 5684 27276
rect 5908 27328 5960 27334
rect 5908 27270 5960 27276
rect 6092 27328 6144 27334
rect 6092 27270 6144 27276
rect 5448 26920 5500 26926
rect 5448 26862 5500 26868
rect 5460 24886 5488 26862
rect 5540 25696 5592 25702
rect 5540 25638 5592 25644
rect 5448 24880 5500 24886
rect 5448 24822 5500 24828
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 5264 23860 5316 23866
rect 5264 23802 5316 23808
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 5276 23361 5304 23598
rect 5460 23594 5488 24686
rect 5552 24274 5580 25638
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 5356 23588 5408 23594
rect 5356 23530 5408 23536
rect 5448 23588 5500 23594
rect 5448 23530 5500 23536
rect 5262 23352 5318 23361
rect 5262 23287 5318 23296
rect 5264 23180 5316 23186
rect 5264 23122 5316 23128
rect 5172 23044 5224 23050
rect 5172 22986 5224 22992
rect 5276 22710 5304 23122
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 5172 22568 5224 22574
rect 5172 22510 5224 22516
rect 5184 20942 5212 22510
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 5184 20058 5212 20402
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5170 19000 5226 19009
rect 5170 18935 5226 18944
rect 5184 18698 5212 18935
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 4986 16960 5042 16969
rect 4986 16895 5042 16904
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4908 16538 4936 16730
rect 4816 16510 4936 16538
rect 4710 16144 4766 16153
rect 4710 16079 4766 16088
rect 4618 14512 4674 14521
rect 4618 14447 4674 14456
rect 4632 14414 4660 14447
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4724 14074 4752 16079
rect 4816 14414 4844 16510
rect 5276 16266 5304 22170
rect 5368 21962 5396 23530
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5460 22234 5488 23054
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5446 22128 5502 22137
rect 5552 22098 5580 23190
rect 5446 22063 5502 22072
rect 5540 22092 5592 22098
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 5354 21176 5410 21185
rect 5354 21111 5356 21120
rect 5408 21111 5410 21120
rect 5356 21082 5408 21088
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5368 18358 5396 20878
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5368 17649 5396 17750
rect 5354 17640 5410 17649
rect 5354 17575 5410 17584
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5368 16697 5396 16934
rect 5354 16688 5410 16697
rect 5354 16623 5410 16632
rect 5000 16238 5304 16266
rect 4894 16144 4950 16153
rect 4894 16079 4950 16088
rect 4908 16046 4936 16079
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4894 15600 4950 15609
rect 4894 15535 4950 15544
rect 4908 15502 4936 15535
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4896 15088 4948 15094
rect 4896 15030 4948 15036
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4436 13864 4488 13870
rect 4436 13806 4488 13812
rect 4908 13682 4936 15030
rect 4816 13654 4936 13682
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 4080 13025 4108 13126
rect 4066 13016 4122 13025
rect 4066 12951 4122 12960
rect 4068 12640 4120 12646
rect 4066 12608 4068 12617
rect 4120 12608 4122 12617
rect 4066 12543 4122 12552
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3988 12406 4108 12434
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3988 11150 4016 12242
rect 4080 11914 4108 12406
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4264 12073 4292 12106
rect 4250 12064 4306 12073
rect 4250 11999 4306 12008
rect 4080 11886 4200 11914
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3974 10840 4030 10849
rect 3974 10775 4030 10784
rect 3988 9178 4016 10775
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 4080 8838 4108 11766
rect 4172 11694 4200 11886
rect 4724 11762 4752 13330
rect 4712 11756 4764 11762
rect 4632 11716 4712 11744
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10248 4660 11716
rect 4712 11698 4764 11704
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4724 11393 4752 11562
rect 4710 11384 4766 11393
rect 4710 11319 4766 11328
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4540 10220 4660 10248
rect 4540 9722 4568 10220
rect 4724 10146 4752 10950
rect 4632 10130 4752 10146
rect 4620 10124 4752 10130
rect 4672 10118 4752 10124
rect 4620 10066 4672 10072
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9042 4660 10066
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4172 8378 4200 8910
rect 4080 8350 4200 8378
rect 4080 7970 4108 8350
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4080 7942 4200 7970
rect 4172 7478 4200 7942
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4172 7290 4200 7414
rect 4264 7410 4292 7890
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4356 7290 4384 8026
rect 4434 7848 4490 7857
rect 4434 7783 4436 7792
rect 4488 7783 4490 7792
rect 4436 7754 4488 7760
rect 4632 7342 4660 8230
rect 4724 8022 4752 9658
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4080 7262 4200 7290
rect 4264 7274 4384 7290
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4252 7268 4384 7274
rect 4080 6882 4108 7262
rect 4304 7262 4384 7268
rect 4252 7210 4304 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4080 6854 4200 6882
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 4172 6322 4200 6854
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4172 6202 4200 6258
rect 4080 6174 4200 6202
rect 4080 5710 4108 6174
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4632 5370 4660 7142
rect 4724 6798 4752 7686
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4356 5030 4384 5170
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 3514 4040 3570 4049
rect 3514 3975 3516 3984
rect 3568 3975 3570 3984
rect 3516 3946 3568 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3528 2825 3556 2994
rect 3514 2816 3570 2825
rect 3514 2751 3570 2760
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2608 800 2636 2382
rect 3988 1465 4016 3470
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2582 4660 4422
rect 4724 3738 4752 6598
rect 4816 6458 4844 13654
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4816 2650 4844 6190
rect 4908 5914 4936 12106
rect 5000 7750 5028 16238
rect 5080 16176 5132 16182
rect 5080 16118 5132 16124
rect 5092 9178 5120 16118
rect 5264 15428 5316 15434
rect 5264 15370 5316 15376
rect 5276 15337 5304 15370
rect 5262 15328 5318 15337
rect 5262 15263 5318 15272
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5276 14550 5304 14826
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5460 14090 5488 22063
rect 5540 22034 5592 22040
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5552 20262 5580 20470
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5538 19000 5594 19009
rect 5538 18935 5594 18944
rect 5552 15434 5580 18935
rect 5644 18698 5672 27270
rect 5920 26450 5948 27270
rect 6104 26450 6132 27270
rect 5908 26444 5960 26450
rect 5908 26386 5960 26392
rect 6092 26444 6144 26450
rect 6092 26386 6144 26392
rect 5908 25764 5960 25770
rect 5908 25706 5960 25712
rect 5816 25288 5868 25294
rect 5816 25230 5868 25236
rect 5828 24954 5856 25230
rect 5816 24948 5868 24954
rect 5816 24890 5868 24896
rect 5722 24848 5778 24857
rect 5722 24783 5778 24792
rect 5816 24812 5868 24818
rect 5736 19786 5764 24783
rect 5816 24754 5868 24760
rect 5828 24206 5856 24754
rect 5816 24200 5868 24206
rect 5816 24142 5868 24148
rect 5920 23497 5948 25706
rect 6092 24948 6144 24954
rect 6092 24890 6144 24896
rect 6000 24608 6052 24614
rect 6000 24550 6052 24556
rect 5906 23488 5962 23497
rect 5906 23423 5962 23432
rect 6012 22522 6040 24550
rect 6104 23322 6132 24890
rect 6196 24274 6224 32166
rect 6276 30728 6328 30734
rect 6276 30670 6328 30676
rect 6288 27130 6316 30670
rect 6564 30258 6592 37130
rect 14844 37126 14872 39200
rect 16132 39114 16160 39200
rect 16224 39114 16252 39222
rect 16132 39086 16252 39114
rect 15200 37256 15252 37262
rect 15200 37198 15252 37204
rect 7196 37120 7248 37126
rect 7196 37062 7248 37068
rect 8300 37120 8352 37126
rect 8300 37062 8352 37068
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 10876 37120 10928 37126
rect 10876 37062 10928 37068
rect 14740 37120 14792 37126
rect 14740 37062 14792 37068
rect 14832 37120 14884 37126
rect 14832 37062 14884 37068
rect 7208 36553 7236 37062
rect 7194 36544 7250 36553
rect 7194 36479 7250 36488
rect 6644 36032 6696 36038
rect 6644 35974 6696 35980
rect 6552 30252 6604 30258
rect 6552 30194 6604 30200
rect 6656 28082 6684 35974
rect 6736 35080 6788 35086
rect 6736 35022 6788 35028
rect 6748 30326 6776 35022
rect 8312 30734 8340 37062
rect 10336 33998 10364 37062
rect 10888 34066 10916 37062
rect 14752 34610 14780 37062
rect 15212 34746 15240 37198
rect 16500 37108 16528 39222
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 20626 39200 20682 39800
rect 22558 39200 22614 39800
rect 23846 39200 23902 39800
rect 25778 39200 25834 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 31574 39200 31630 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 16580 37120 16632 37126
rect 16500 37080 16580 37108
rect 16580 37062 16632 37068
rect 16868 35834 16896 37198
rect 18064 37126 18092 39200
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 18236 37256 18288 37262
rect 18236 37198 18288 37204
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 16856 35828 16908 35834
rect 16856 35770 16908 35776
rect 17040 35692 17092 35698
rect 17040 35634 17092 35640
rect 16488 35080 16540 35086
rect 16488 35022 16540 35028
rect 15200 34740 15252 34746
rect 15200 34682 15252 34688
rect 12072 34604 12124 34610
rect 12072 34546 12124 34552
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 15660 34604 15712 34610
rect 15660 34546 15712 34552
rect 10876 34060 10928 34066
rect 10876 34002 10928 34008
rect 10324 33992 10376 33998
rect 10324 33934 10376 33940
rect 8392 33856 8444 33862
rect 8392 33798 8444 33804
rect 10232 33856 10284 33862
rect 10232 33798 10284 33804
rect 8300 30728 8352 30734
rect 8300 30670 8352 30676
rect 8208 30592 8260 30598
rect 8208 30534 8260 30540
rect 6736 30320 6788 30326
rect 6736 30262 6788 30268
rect 7748 30048 7800 30054
rect 7748 29990 7800 29996
rect 7472 29572 7524 29578
rect 7472 29514 7524 29520
rect 6644 28076 6696 28082
rect 6644 28018 6696 28024
rect 7104 27532 7156 27538
rect 7104 27474 7156 27480
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6276 27124 6328 27130
rect 6276 27066 6328 27072
rect 6288 26586 6316 27066
rect 6276 26580 6328 26586
rect 6276 26522 6328 26528
rect 6840 25974 6868 27338
rect 6828 25968 6880 25974
rect 6828 25910 6880 25916
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 6828 25832 6880 25838
rect 6828 25774 6880 25780
rect 6460 25696 6512 25702
rect 6460 25638 6512 25644
rect 6472 25294 6500 25638
rect 6460 25288 6512 25294
rect 6460 25230 6512 25236
rect 6840 25226 6868 25774
rect 6276 25220 6328 25226
rect 6276 25162 6328 25168
rect 6828 25220 6880 25226
rect 6828 25162 6880 25168
rect 6288 24290 6316 25162
rect 6552 25152 6604 25158
rect 6552 25094 6604 25100
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6564 24562 6592 25094
rect 6564 24534 6684 24562
rect 6184 24268 6236 24274
rect 6288 24262 6500 24290
rect 6184 24210 6236 24216
rect 6276 24200 6328 24206
rect 6276 24142 6328 24148
rect 6092 23316 6144 23322
rect 6092 23258 6144 23264
rect 6184 22976 6236 22982
rect 6184 22918 6236 22924
rect 6196 22710 6224 22918
rect 6184 22704 6236 22710
rect 6184 22646 6236 22652
rect 5920 22494 6040 22522
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5828 22273 5856 22374
rect 5814 22264 5870 22273
rect 5814 22199 5870 22208
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5736 18834 5764 19246
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 5632 18692 5684 18698
rect 5632 18634 5684 18640
rect 5736 18290 5764 18770
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 5276 14062 5488 14090
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5092 7954 5120 8978
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 5184 7546 5212 11018
rect 5276 10606 5304 14062
rect 5356 14000 5408 14006
rect 5356 13942 5408 13948
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5276 9926 5304 10542
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5276 7818 5304 9522
rect 5368 9110 5396 13942
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 11830 5488 13262
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12306 5580 12582
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5446 11520 5502 11529
rect 5446 11455 5502 11464
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5460 8974 5488 11455
rect 5552 9081 5580 11698
rect 5644 11082 5672 12106
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 10305 5672 10406
rect 5630 10296 5686 10305
rect 5630 10231 5686 10240
rect 5538 9072 5594 9081
rect 5538 9007 5594 9016
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5276 7698 5304 7754
rect 5276 7670 5396 7698
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5000 5370 5028 7414
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5092 5914 5120 7278
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4908 4146 4936 5170
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5276 3194 5304 6258
rect 5368 5234 5396 7670
rect 5460 7546 5488 8910
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5460 6798 5488 7482
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5552 3126 5580 8842
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5644 8634 5672 8774
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5630 8528 5686 8537
rect 5630 8463 5686 8472
rect 5644 8430 5672 8463
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5736 6866 5764 14282
rect 5828 14006 5856 21830
rect 5920 20874 5948 22494
rect 6288 21894 6316 24142
rect 6368 23656 6420 23662
rect 6368 23598 6420 23604
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 5908 20868 5960 20874
rect 5908 20810 5960 20816
rect 6196 20058 6224 21490
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 6288 20210 6316 20402
rect 6380 20398 6408 23598
rect 6472 21622 6500 24262
rect 6656 24138 6684 24534
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6748 22710 6776 25094
rect 6736 22704 6788 22710
rect 6736 22646 6788 22652
rect 6840 22556 6868 25162
rect 7024 23798 7052 25842
rect 7012 23792 7064 23798
rect 7012 23734 7064 23740
rect 7024 23610 7052 23734
rect 6932 23582 7052 23610
rect 6932 22710 6960 23582
rect 6920 22704 6972 22710
rect 7116 22658 7144 27474
rect 7288 27464 7340 27470
rect 7288 27406 7340 27412
rect 7300 26994 7328 27406
rect 7288 26988 7340 26994
rect 7288 26930 7340 26936
rect 6920 22646 6972 22652
rect 6748 22528 6868 22556
rect 7024 22630 7144 22658
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6460 21616 6512 21622
rect 6460 21558 6512 21564
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6288 20182 6408 20210
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6288 19922 6316 19994
rect 6380 19922 6408 20182
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 5920 19446 5948 19654
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 6380 18902 6408 19858
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6104 18222 6132 18838
rect 6472 18714 6500 21558
rect 6656 19334 6684 21830
rect 6196 18686 6500 18714
rect 6564 19306 6684 19334
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6090 18048 6146 18057
rect 6090 17983 6146 17992
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5920 12434 5948 16458
rect 6000 15428 6052 15434
rect 6000 15370 6052 15376
rect 5828 12406 5948 12434
rect 5828 7954 5856 12406
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11762 5948 12038
rect 6012 11898 6040 15370
rect 6104 13802 6132 17983
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6104 12782 6132 13126
rect 6092 12776 6144 12782
rect 6090 12744 6092 12753
rect 6144 12744 6146 12753
rect 6090 12679 6146 12688
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5998 11248 6054 11257
rect 5998 11183 6054 11192
rect 6012 10674 6040 11183
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6104 10554 6132 12582
rect 5920 10526 6132 10554
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 4622 5672 5510
rect 5828 4758 5856 7754
rect 5920 5710 5948 10526
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 10266 6132 10406
rect 6196 10266 6224 18686
rect 6366 17640 6422 17649
rect 6366 17575 6368 17584
rect 6420 17575 6422 17584
rect 6368 17546 6420 17552
rect 6564 17066 6592 19306
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6656 17202 6684 18158
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6552 16040 6604 16046
rect 6550 16008 6552 16017
rect 6604 16008 6606 16017
rect 6550 15943 6606 15952
rect 6460 14952 6512 14958
rect 6512 14900 6592 14906
rect 6460 14894 6592 14900
rect 6472 14878 6592 14894
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6366 14784 6422 14793
rect 6288 13734 6316 14758
rect 6366 14719 6422 14728
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6288 12434 6316 12854
rect 6380 12646 6408 14719
rect 6460 13252 6512 13258
rect 6460 13194 6512 13200
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6288 12406 6408 12434
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6288 10742 6316 11154
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6380 10198 6408 12406
rect 6472 11234 6500 13194
rect 6564 12442 6592 14878
rect 6656 12442 6684 16934
rect 6748 15638 6776 22528
rect 7024 22094 7052 22630
rect 7104 22500 7156 22506
rect 7104 22442 7156 22448
rect 6932 22066 7052 22094
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6840 20806 6868 21830
rect 6932 21026 6960 22066
rect 7116 21350 7144 22442
rect 7300 22166 7328 26930
rect 7380 25900 7432 25906
rect 7380 25842 7432 25848
rect 7392 25294 7420 25842
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7392 24070 7420 25230
rect 7380 24064 7432 24070
rect 7380 24006 7432 24012
rect 7288 22160 7340 22166
rect 7288 22102 7340 22108
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 6932 20998 7052 21026
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6840 16590 6868 20742
rect 6918 20632 6974 20641
rect 6918 20567 6920 20576
rect 6972 20567 6974 20576
rect 6920 20538 6972 20544
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6932 18766 6960 19994
rect 7024 19922 7052 20998
rect 7116 20466 7144 21286
rect 7300 20806 7328 22102
rect 7484 21622 7512 29514
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7668 26246 7696 26862
rect 7656 26240 7708 26246
rect 7656 26182 7708 26188
rect 7668 26042 7696 26182
rect 7656 26036 7708 26042
rect 7656 25978 7708 25984
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7472 21616 7524 21622
rect 7472 21558 7524 21564
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7288 20800 7340 20806
rect 7288 20742 7340 20748
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7484 20398 7512 20878
rect 7472 20392 7524 20398
rect 7286 20360 7342 20369
rect 7472 20334 7524 20340
rect 7286 20295 7288 20304
rect 7340 20295 7342 20304
rect 7288 20266 7340 20272
rect 7484 20262 7512 20334
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7392 19990 7420 20198
rect 7380 19984 7432 19990
rect 7380 19926 7432 19932
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7116 19174 7144 19654
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 7208 18426 7236 19110
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7104 17536 7156 17542
rect 7010 17504 7066 17513
rect 7104 17478 7156 17484
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7010 17439 7066 17448
rect 7024 17270 7052 17439
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 6840 16250 6868 16526
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6748 14464 6776 15574
rect 6840 14906 6868 16186
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6932 15881 6960 15914
rect 6918 15872 6974 15881
rect 6918 15807 6974 15816
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6932 15094 6960 15438
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6840 14878 6960 14906
rect 6748 14436 6868 14464
rect 6840 14074 6868 14436
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6932 13954 6960 14878
rect 7024 14482 7052 16662
rect 7116 15910 7144 17478
rect 7208 17202 7236 17478
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7300 15586 7328 19314
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7392 17134 7420 17682
rect 7484 17678 7512 18158
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7392 16046 7420 17070
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7208 15558 7328 15586
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 6748 13926 6960 13954
rect 6748 12918 6776 13926
rect 6918 13696 6974 13705
rect 6918 13631 6974 13640
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6472 11206 6592 11234
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6196 9042 6224 9454
rect 6366 9072 6422 9081
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6184 9036 6236 9042
rect 6366 9007 6422 9016
rect 6184 8978 6236 8984
rect 6012 8498 6040 8978
rect 6380 8498 6408 9007
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 6012 5642 6040 6870
rect 6380 6390 6408 8434
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5642 6408 6054
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6472 4826 6500 11018
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 6564 4690 6592 11206
rect 6642 10840 6698 10849
rect 6642 10775 6644 10784
rect 6696 10775 6698 10784
rect 6644 10746 6696 10752
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6656 10198 6684 10610
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6748 9654 6776 12854
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6840 11801 6868 12786
rect 6932 12238 6960 13631
rect 7208 12866 7236 15558
rect 7472 15496 7524 15502
rect 7286 15464 7342 15473
rect 7472 15438 7524 15444
rect 7286 15399 7288 15408
rect 7340 15399 7342 15408
rect 7288 15370 7340 15376
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7392 14482 7420 14758
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7300 13190 7328 13262
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7208 12850 7328 12866
rect 7104 12844 7156 12850
rect 7208 12844 7340 12850
rect 7208 12838 7288 12844
rect 7104 12786 7156 12792
rect 7288 12786 7340 12792
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6826 11792 6882 11801
rect 6826 11727 6882 11736
rect 6840 10810 6868 11727
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 7024 10130 7052 12242
rect 7116 10792 7144 12786
rect 7116 10764 7236 10792
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 7546 6684 7890
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 6656 2854 6684 7346
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6748 5914 6776 6258
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6748 5778 6776 5850
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6840 5098 6868 8570
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6932 2922 6960 8298
rect 7024 5166 7052 9930
rect 7104 9648 7156 9654
rect 7102 9616 7104 9625
rect 7156 9616 7158 9625
rect 7102 9551 7158 9560
rect 7208 6934 7236 10764
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7300 9654 7328 10678
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7300 8634 7328 8842
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7300 8498 7328 8570
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7392 8294 7420 14282
rect 7484 13462 7512 15438
rect 7472 13456 7524 13462
rect 7472 13398 7524 13404
rect 7472 11824 7524 11830
rect 7470 11792 7472 11801
rect 7524 11792 7526 11801
rect 7470 11727 7526 11736
rect 7576 9602 7604 24346
rect 7668 23798 7696 25094
rect 7760 24410 7788 29990
rect 8024 29504 8076 29510
rect 8024 29446 8076 29452
rect 7932 27872 7984 27878
rect 7932 27814 7984 27820
rect 7840 25152 7892 25158
rect 7840 25094 7892 25100
rect 7852 24818 7880 25094
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7944 24750 7972 27814
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 7760 24138 7788 24346
rect 7852 24138 7880 24550
rect 7748 24132 7800 24138
rect 7748 24074 7800 24080
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 7656 23792 7708 23798
rect 7656 23734 7708 23740
rect 7932 22772 7984 22778
rect 7932 22714 7984 22720
rect 7656 22432 7708 22438
rect 7656 22374 7708 22380
rect 7668 19281 7696 22374
rect 7944 22137 7972 22714
rect 7930 22128 7986 22137
rect 7930 22063 7986 22072
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7654 19272 7710 19281
rect 7654 19207 7710 19216
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7668 18873 7696 19110
rect 7654 18864 7710 18873
rect 7654 18799 7710 18808
rect 7656 17264 7708 17270
rect 7656 17206 7708 17212
rect 7668 12306 7696 17206
rect 7760 16046 7788 20742
rect 7840 20528 7892 20534
rect 7840 20470 7892 20476
rect 7852 20398 7880 20470
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7852 17814 7880 18702
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7852 16182 7880 17478
rect 7944 17218 7972 22063
rect 8036 20233 8064 29446
rect 8220 26518 8248 30534
rect 8208 26512 8260 26518
rect 8208 26454 8260 26460
rect 8220 26382 8248 26454
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8404 25906 8432 33798
rect 9128 30864 9180 30870
rect 9128 30806 9180 30812
rect 9140 27470 9168 30806
rect 9864 29708 9916 29714
rect 9864 29650 9916 29656
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9220 27328 9272 27334
rect 9220 27270 9272 27276
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8116 25424 8168 25430
rect 8116 25366 8168 25372
rect 8128 22642 8156 25366
rect 8588 25294 8616 26862
rect 9048 26382 9076 26930
rect 9036 26376 9088 26382
rect 9036 26318 9088 26324
rect 8668 25696 8720 25702
rect 8668 25638 8720 25644
rect 8576 25288 8628 25294
rect 8496 25248 8576 25276
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8208 24132 8260 24138
rect 8208 24074 8260 24080
rect 8220 23662 8248 24074
rect 8208 23656 8260 23662
rect 8208 23598 8260 23604
rect 8300 23248 8352 23254
rect 8300 23190 8352 23196
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8220 22778 8248 23054
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8206 22264 8262 22273
rect 8206 22199 8262 22208
rect 8220 21570 8248 22199
rect 8312 21690 8340 23190
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 8220 21542 8340 21570
rect 8208 20868 8260 20874
rect 8208 20810 8260 20816
rect 8022 20224 8078 20233
rect 8022 20159 8078 20168
rect 8220 19854 8248 20810
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8128 18834 8156 19450
rect 8220 18873 8248 19790
rect 8206 18864 8262 18873
rect 8116 18828 8168 18834
rect 8206 18799 8262 18808
rect 8116 18770 8168 18776
rect 8312 18426 8340 21542
rect 8404 19802 8432 24754
rect 8496 23610 8524 25248
rect 8576 25230 8628 25236
rect 8680 24750 8708 25638
rect 8760 25288 8812 25294
rect 8760 25230 8812 25236
rect 8772 24954 8800 25230
rect 8760 24948 8812 24954
rect 8760 24890 8812 24896
rect 8668 24744 8720 24750
rect 8668 24686 8720 24692
rect 8576 24132 8628 24138
rect 8576 24074 8628 24080
rect 8588 23730 8616 24074
rect 8680 23798 8708 24686
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8956 24342 8984 24550
rect 8944 24336 8996 24342
rect 8944 24278 8996 24284
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 8668 23792 8720 23798
rect 8668 23734 8720 23740
rect 8758 23760 8814 23769
rect 8576 23724 8628 23730
rect 8758 23695 8814 23704
rect 8576 23666 8628 23672
rect 8496 23582 8708 23610
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8496 23186 8524 23462
rect 8484 23180 8536 23186
rect 8484 23122 8536 23128
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8496 21486 8524 21626
rect 8484 21480 8536 21486
rect 8484 21422 8536 21428
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8496 20874 8524 21286
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 8404 19774 8524 19802
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19514 8432 19654
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8208 18352 8260 18358
rect 8114 18320 8170 18329
rect 8208 18294 8260 18300
rect 8114 18255 8170 18264
rect 8128 18222 8156 18255
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8128 18057 8156 18158
rect 8114 18048 8170 18057
rect 8114 17983 8170 17992
rect 7944 17190 8064 17218
rect 7840 16176 7892 16182
rect 7840 16118 7892 16124
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7930 15192 7986 15201
rect 7930 15127 7986 15136
rect 7944 15026 7972 15127
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7852 14550 7880 14894
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7760 11880 7788 12106
rect 7668 11852 7788 11880
rect 7668 11218 7696 11852
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7472 9580 7524 9586
rect 7576 9574 7696 9602
rect 7472 9522 7524 9528
rect 7484 8786 7512 9522
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 8906 7604 9386
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7484 8758 7604 8786
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7484 8401 7512 8434
rect 7470 8392 7526 8401
rect 7470 8327 7526 8336
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7392 8090 7420 8230
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 7300 2650 7328 7822
rect 7576 5642 7604 8758
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7576 5030 7604 5578
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7668 4690 7696 9574
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7760 3670 7788 11698
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7852 11529 7880 11562
rect 7838 11520 7894 11529
rect 7838 11455 7894 11464
rect 7838 11112 7894 11121
rect 7838 11047 7894 11056
rect 7852 9382 7880 11047
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7944 9178 7972 12582
rect 8036 12306 8064 17190
rect 8220 16454 8248 18294
rect 8496 17610 8524 19774
rect 8588 17882 8616 23462
rect 8680 19281 8708 23582
rect 8772 20534 8800 23695
rect 8864 21486 8892 24006
rect 8956 23526 8984 24278
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8956 22817 8984 22918
rect 8942 22808 8998 22817
rect 8942 22743 8998 22752
rect 8956 22710 8984 22743
rect 8944 22704 8996 22710
rect 8944 22646 8996 22652
rect 9048 22234 9076 26318
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 9140 23730 9168 24550
rect 9128 23724 9180 23730
rect 9128 23666 9180 23672
rect 9232 23050 9260 27270
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9784 25838 9812 26182
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9496 25220 9548 25226
rect 9496 25162 9548 25168
rect 9312 25152 9364 25158
rect 9312 25094 9364 25100
rect 9324 24954 9352 25094
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9324 23866 9352 24142
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9416 23798 9444 24006
rect 9404 23792 9456 23798
rect 9404 23734 9456 23740
rect 9404 23520 9456 23526
rect 9404 23462 9456 23468
rect 9220 23044 9272 23050
rect 9220 22986 9272 22992
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 9036 22228 9088 22234
rect 9036 22170 9088 22176
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 8864 20806 8892 20878
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8760 20528 8812 20534
rect 8760 20470 8812 20476
rect 8758 20224 8814 20233
rect 8758 20159 8814 20168
rect 8772 19786 8800 20159
rect 8864 19922 8892 20742
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8760 19780 8812 19786
rect 8760 19722 8812 19728
rect 8666 19272 8722 19281
rect 8666 19207 8722 19216
rect 8680 18902 8708 19207
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8956 18630 8984 22034
rect 9140 21962 9168 22714
rect 9220 22228 9272 22234
rect 9220 22170 9272 22176
rect 9128 21956 9180 21962
rect 9128 21898 9180 21904
rect 9140 21350 9168 21898
rect 9232 21570 9260 22170
rect 9312 22160 9364 22166
rect 9310 22128 9312 22137
rect 9364 22128 9366 22137
rect 9310 22063 9366 22072
rect 9232 21542 9352 21570
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 9140 20942 9168 21286
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 9048 20058 9076 20402
rect 9140 20262 9168 20878
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9140 19922 9168 20198
rect 9232 20058 9260 21422
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9048 19768 9076 19858
rect 9048 19740 9168 19768
rect 9034 19408 9090 19417
rect 9034 19343 9090 19352
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8772 17898 8800 18362
rect 8944 18352 8996 18358
rect 8944 18294 8996 18300
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8668 17876 8720 17882
rect 8772 17870 8892 17898
rect 8668 17818 8720 17824
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8576 17604 8628 17610
rect 8576 17546 8628 17552
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8114 16144 8170 16153
rect 8114 16079 8170 16088
rect 8128 16046 8156 16079
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8220 15910 8248 16390
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8128 13258 8156 14282
rect 8220 14006 8248 15846
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 8036 8634 8064 10610
rect 8114 10296 8170 10305
rect 8114 10231 8116 10240
rect 8168 10231 8170 10240
rect 8116 10202 8168 10208
rect 8220 9994 8248 13670
rect 8312 13326 8340 17546
rect 8496 15473 8524 17546
rect 8588 16289 8616 17546
rect 8680 17338 8708 17818
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8574 16280 8630 16289
rect 8772 16266 8800 17750
rect 8864 16590 8892 17870
rect 8956 17649 8984 18294
rect 8942 17640 8998 17649
rect 8942 17575 8998 17584
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8956 16726 8984 17274
rect 8944 16720 8996 16726
rect 8944 16662 8996 16668
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8574 16215 8630 16224
rect 8680 16238 8800 16266
rect 8482 15464 8538 15473
rect 8482 15399 8538 15408
rect 8496 15366 8524 15399
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8404 14414 8432 15302
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8588 14074 8616 14214
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8390 13968 8446 13977
rect 8390 13903 8446 13912
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8404 12102 8432 13903
rect 8680 13734 8708 16238
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8484 13320 8536 13326
rect 8482 13288 8484 13297
rect 8536 13288 8538 13297
rect 8482 13223 8538 13232
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8496 12306 8524 13126
rect 8588 12986 8616 13126
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8496 11880 8524 12242
rect 8496 11852 8616 11880
rect 8482 11792 8538 11801
rect 8482 11727 8538 11736
rect 8300 11552 8352 11558
rect 8392 11552 8444 11558
rect 8300 11494 8352 11500
rect 8390 11520 8392 11529
rect 8444 11520 8446 11529
rect 8312 11218 8340 11494
rect 8390 11455 8446 11464
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8496 11014 8524 11727
rect 8588 11257 8616 11852
rect 8574 11248 8630 11257
rect 8574 11183 8630 11192
rect 8588 11150 8616 11183
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8588 10130 8616 11086
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8312 9722 8340 10066
rect 8680 9926 8708 11018
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8116 9648 8168 9654
rect 8114 9616 8116 9625
rect 8168 9616 8170 9625
rect 8114 9551 8170 9560
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8114 8664 8170 8673
rect 8024 8628 8076 8634
rect 8114 8599 8170 8608
rect 8024 8570 8076 8576
rect 8128 8566 8156 8599
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8220 8430 8248 9318
rect 8312 9042 8340 9658
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8208 8424 8260 8430
rect 8404 8401 8432 9658
rect 8496 9178 8524 9862
rect 8772 9518 8800 16118
rect 8944 15632 8996 15638
rect 8944 15574 8996 15580
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8864 14958 8892 15438
rect 8956 15434 8984 15574
rect 8944 15428 8996 15434
rect 8944 15370 8996 15376
rect 9048 15094 9076 19343
rect 9140 17202 9168 19740
rect 9218 19680 9274 19689
rect 9218 19615 9274 19624
rect 9232 18834 9260 19615
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9218 17368 9274 17377
rect 9218 17303 9274 17312
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9232 16998 9260 17303
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9140 16794 9168 16934
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9324 16658 9352 21542
rect 9416 17270 9444 23462
rect 9508 20806 9536 25162
rect 9692 24818 9720 25638
rect 9772 25424 9824 25430
rect 9772 25366 9824 25372
rect 9784 25158 9812 25366
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 9876 24698 9904 29650
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9968 26382 9996 26726
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 10244 25906 10272 33798
rect 12084 29850 12112 34546
rect 15672 33658 15700 34546
rect 16120 34536 16172 34542
rect 16120 34478 16172 34484
rect 15660 33652 15712 33658
rect 15660 33594 15712 33600
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 12164 33380 12216 33386
rect 12164 33322 12216 33328
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 12072 26376 12124 26382
rect 12072 26318 12124 26324
rect 10980 25906 11008 26318
rect 11060 26308 11112 26314
rect 11060 26250 11112 26256
rect 11888 26308 11940 26314
rect 11888 26250 11940 26256
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 10048 25832 10100 25838
rect 10048 25774 10100 25780
rect 10060 25498 10088 25774
rect 10048 25492 10100 25498
rect 10048 25434 10100 25440
rect 10336 25158 10364 25842
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10322 24848 10378 24857
rect 9956 24812 10008 24818
rect 10322 24783 10324 24792
rect 9956 24754 10008 24760
rect 10376 24783 10378 24792
rect 10324 24754 10376 24760
rect 9692 24670 9904 24698
rect 9586 22808 9642 22817
rect 9586 22743 9588 22752
rect 9640 22743 9642 22752
rect 9588 22714 9640 22720
rect 9586 22672 9642 22681
rect 9586 22607 9588 22616
rect 9640 22607 9642 22616
rect 9588 22578 9640 22584
rect 9588 22092 9640 22098
rect 9692 22094 9720 24670
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9876 24410 9904 24550
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 9784 22574 9812 24346
rect 9968 23594 9996 24754
rect 10428 24698 10456 25434
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10336 24670 10456 24698
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 9954 23080 10010 23089
rect 9864 23044 9916 23050
rect 9954 23015 10010 23024
rect 9864 22986 9916 22992
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 9876 22438 9904 22986
rect 9968 22642 9996 23015
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 9772 22432 9824 22438
rect 9770 22400 9772 22409
rect 9864 22432 9916 22438
rect 9824 22400 9826 22409
rect 9864 22374 9916 22380
rect 9770 22335 9826 22344
rect 9692 22066 9904 22094
rect 9588 22034 9640 22040
rect 9600 21418 9628 22034
rect 9588 21412 9640 21418
rect 9588 21354 9640 21360
rect 9876 20874 9904 22066
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9680 20800 9732 20806
rect 10060 20754 10088 24210
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10152 22642 10180 24006
rect 10336 23322 10364 24670
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10324 23316 10376 23322
rect 10324 23258 10376 23264
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10140 21616 10192 21622
rect 10138 21584 10140 21593
rect 10192 21584 10194 21593
rect 10336 21554 10364 23258
rect 10428 22030 10456 24550
rect 10612 23186 10640 25094
rect 11072 24274 11100 26250
rect 11612 25900 11664 25906
rect 11612 25842 11664 25848
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 11164 24993 11192 25094
rect 11150 24984 11206 24993
rect 11150 24919 11206 24928
rect 11152 24744 11204 24750
rect 11152 24686 11204 24692
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10968 23588 11020 23594
rect 10968 23530 11020 23536
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10980 22574 11008 23530
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 11072 22710 11100 23462
rect 11164 23186 11192 24686
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 11256 23066 11284 24550
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11164 23038 11284 23066
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10138 21519 10194 21528
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 9680 20742 9732 20748
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9586 20360 9642 20369
rect 9508 19417 9536 20334
rect 9586 20295 9642 20304
rect 9600 20262 9628 20295
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9692 19446 9720 20742
rect 9784 20726 10088 20754
rect 10230 20768 10286 20777
rect 9680 19440 9732 19446
rect 9494 19408 9550 19417
rect 9680 19382 9732 19388
rect 9494 19343 9550 19352
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9600 19281 9628 19314
rect 9680 19304 9732 19310
rect 9586 19272 9642 19281
rect 9680 19246 9732 19252
rect 9586 19207 9642 19216
rect 9588 19168 9640 19174
rect 9586 19136 9588 19145
rect 9640 19136 9642 19145
rect 9586 19071 9642 19080
rect 9496 18760 9548 18766
rect 9494 18728 9496 18737
rect 9548 18728 9550 18737
rect 9494 18663 9550 18672
rect 9692 18222 9720 19246
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9508 16794 9536 17138
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9232 16266 9260 16526
rect 9232 16238 9352 16266
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9140 15910 9168 16050
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 9036 15088 9088 15094
rect 9034 15056 9036 15065
rect 9088 15056 9090 15065
rect 9034 14991 9090 15000
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9048 13938 9076 14418
rect 9140 14346 9168 15846
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9048 13394 9076 13874
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 9048 12986 9076 13330
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8864 11082 8892 12038
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8537 8524 8978
rect 8864 8838 8892 11018
rect 8956 10169 8984 12650
rect 9048 12238 9076 12922
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9048 11744 9076 12174
rect 9128 11756 9180 11762
rect 9048 11716 9128 11744
rect 9128 11698 9180 11704
rect 8942 10160 8998 10169
rect 8942 10095 8998 10104
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 9232 8634 9260 14894
rect 9324 14006 9352 16238
rect 9404 15904 9456 15910
rect 9402 15872 9404 15881
rect 9456 15872 9458 15881
rect 9402 15807 9458 15816
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9324 13734 9352 13942
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9324 12646 9352 13194
rect 9416 12714 9444 14282
rect 9508 13569 9536 16526
rect 9784 16182 9812 20726
rect 10230 20703 10286 20712
rect 10244 20602 10272 20703
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 9862 20496 9918 20505
rect 10336 20482 10364 21490
rect 9862 20431 9864 20440
rect 9916 20431 9918 20440
rect 10244 20454 10364 20482
rect 9864 20402 9916 20408
rect 9954 19816 10010 19825
rect 9954 19751 10010 19760
rect 9968 19514 9996 19751
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9772 16176 9824 16182
rect 9678 16144 9734 16153
rect 9772 16118 9824 16124
rect 9678 16079 9734 16088
rect 9692 16046 9720 16079
rect 9680 16040 9732 16046
rect 9876 16017 9904 19314
rect 10138 18728 10194 18737
rect 10138 18663 10194 18672
rect 10048 18352 10100 18358
rect 9968 18312 10048 18340
rect 9968 18222 9996 18312
rect 10048 18294 10100 18300
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9680 15982 9732 15988
rect 9862 16008 9918 16017
rect 9862 15943 9918 15952
rect 10152 15688 10180 18663
rect 10244 18426 10272 20454
rect 10324 19780 10376 19786
rect 10324 19722 10376 19728
rect 10336 19378 10364 19722
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10598 19272 10654 19281
rect 10598 19207 10600 19216
rect 10652 19207 10654 19216
rect 10600 19178 10652 19184
rect 10598 18728 10654 18737
rect 10598 18663 10600 18672
rect 10652 18663 10654 18672
rect 10600 18634 10652 18640
rect 10796 18630 10824 22442
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10888 18850 10916 19722
rect 10980 19378 11008 22510
rect 11164 22094 11192 23038
rect 11244 22094 11296 22098
rect 11164 22092 11296 22094
rect 11164 22066 11244 22092
rect 11244 22034 11296 22040
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11072 20398 11100 20878
rect 11348 20398 11376 24142
rect 11532 23662 11560 24210
rect 11624 23866 11652 25842
rect 11704 25764 11756 25770
rect 11704 25706 11756 25712
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11716 23730 11744 25706
rect 11796 24948 11848 24954
rect 11796 24890 11848 24896
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11520 23656 11572 23662
rect 11520 23598 11572 23604
rect 11428 22704 11480 22710
rect 11428 22646 11480 22652
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 10968 19372 11020 19378
rect 11348 19334 11376 20334
rect 10968 19314 11020 19320
rect 11256 19306 11376 19334
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 10888 18822 11008 18850
rect 11072 18834 11100 19110
rect 11150 18864 11206 18873
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10704 18358 10732 18566
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10888 18290 10916 18702
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10244 17338 10272 17478
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 9876 15660 10180 15688
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9494 13560 9550 13569
rect 9494 13495 9550 13504
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 8482 8528 8538 8537
rect 8482 8463 8538 8472
rect 8208 8366 8260 8372
rect 8390 8392 8446 8401
rect 8390 8327 8446 8336
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7944 5234 7972 5646
rect 8496 5302 8524 7686
rect 9218 7576 9274 7585
rect 9218 7511 9220 7520
rect 9272 7511 9274 7520
rect 9220 7482 9272 7488
rect 9324 6848 9352 12106
rect 9404 11144 9456 11150
rect 9496 11144 9548 11150
rect 9404 11086 9456 11092
rect 9494 11112 9496 11121
rect 9548 11112 9550 11121
rect 9416 10674 9444 11086
rect 9494 11047 9550 11056
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9508 10470 9536 10950
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9600 6866 9628 14214
rect 9692 10742 9720 15302
rect 9876 14822 9904 15660
rect 10244 15586 10272 16118
rect 10336 15978 10364 18158
rect 10598 17776 10654 17785
rect 10598 17711 10654 17720
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10520 17513 10548 17546
rect 10506 17504 10562 17513
rect 10506 17439 10562 17448
rect 10612 17134 10640 17711
rect 10888 17678 10916 18226
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10888 17202 10916 17614
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10520 15638 10548 16458
rect 10060 15558 10272 15586
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 10060 14618 10088 15558
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9968 12434 9996 14282
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 10060 12889 10088 13194
rect 10046 12880 10102 12889
rect 10046 12815 10102 12824
rect 9876 12406 9996 12434
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9692 10441 9720 10678
rect 9678 10432 9734 10441
rect 9678 10367 9734 10376
rect 9678 10296 9734 10305
rect 9678 10231 9680 10240
rect 9732 10231 9734 10240
rect 9680 10202 9732 10208
rect 9680 9920 9732 9926
rect 9678 9888 9680 9897
rect 9732 9888 9734 9897
rect 9678 9823 9734 9832
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 8974 9720 9522
rect 9784 9178 9812 11698
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9876 8650 9904 12406
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9784 8622 9904 8650
rect 9784 8022 9812 8622
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9232 6820 9352 6848
rect 9588 6860 9640 6866
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8772 6458 8800 6666
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8588 5914 8616 6258
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7944 4622 7972 5170
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 9232 4078 9260 6820
rect 9588 6802 9640 6808
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9324 6458 9352 6666
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9600 5846 9628 6802
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 9600 3058 9628 3878
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 9416 2446 9444 2790
rect 9876 2650 9904 8434
rect 9968 5914 9996 11630
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10060 8634 10088 11018
rect 10152 9110 10180 15370
rect 10416 15360 10468 15366
rect 10322 15328 10378 15337
rect 10468 15308 10640 15314
rect 10416 15302 10640 15308
rect 10428 15286 10640 15302
rect 10322 15263 10378 15272
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10244 14793 10272 14826
rect 10230 14784 10286 14793
rect 10230 14719 10286 14728
rect 10336 13802 10364 15263
rect 10506 15056 10562 15065
rect 10506 14991 10508 15000
rect 10560 14991 10562 15000
rect 10508 14962 10560 14968
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10428 13841 10456 13874
rect 10414 13832 10470 13841
rect 10324 13796 10376 13802
rect 10414 13767 10470 13776
rect 10324 13738 10376 13744
rect 10336 11830 10364 13738
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10336 11370 10364 11766
rect 10428 11558 10456 12718
rect 10520 12170 10548 14758
rect 10612 14521 10640 15286
rect 10598 14512 10654 14521
rect 10598 14447 10600 14456
rect 10652 14447 10654 14456
rect 10600 14418 10652 14424
rect 10612 14387 10640 14418
rect 10704 13530 10732 17070
rect 10888 16658 10916 17138
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10980 16538 11008 18822
rect 11060 18828 11112 18834
rect 11150 18799 11152 18808
rect 11060 18770 11112 18776
rect 11204 18799 11206 18808
rect 11152 18770 11204 18776
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10796 16510 11008 16538
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10796 13394 10824 16510
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 15978 10916 16390
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10888 14618 10916 15914
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10782 13288 10838 13297
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10612 12782 10640 12922
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10704 12434 10732 13262
rect 10782 13223 10838 13232
rect 10796 13190 10824 13223
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10612 12406 10732 12434
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10336 11342 10456 11370
rect 10612 11354 10640 12406
rect 10888 11762 10916 14418
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10692 11688 10744 11694
rect 10980 11642 11008 15030
rect 11072 14958 11100 18158
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11060 14816 11112 14822
rect 11058 14784 11060 14793
rect 11112 14784 11114 14793
rect 11058 14719 11114 14728
rect 11164 13870 11192 17546
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11150 12744 11206 12753
rect 11150 12679 11152 12688
rect 11204 12679 11206 12688
rect 11152 12650 11204 12656
rect 11256 12306 11284 19306
rect 11440 17746 11468 22646
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 11612 21004 11664 21010
rect 11612 20946 11664 20952
rect 11624 20466 11652 20946
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11716 17814 11744 22034
rect 11808 19922 11836 24890
rect 11900 24800 11928 26250
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 11992 24954 12020 25638
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 11980 24812 12032 24818
rect 11900 24772 11980 24800
rect 11980 24754 12032 24760
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 11900 22574 11928 24346
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11992 23662 12020 24006
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 11992 22506 12020 23598
rect 11980 22500 12032 22506
rect 11980 22442 12032 22448
rect 11888 22092 11940 22098
rect 12084 22094 12112 26318
rect 11888 22034 11940 22040
rect 11992 22066 12112 22094
rect 11900 21418 11928 22034
rect 11888 21412 11940 21418
rect 11888 21354 11940 21360
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 11886 19408 11942 19417
rect 11886 19343 11888 19352
rect 11940 19343 11942 19352
rect 11888 19314 11940 19320
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11612 17060 11664 17066
rect 11612 17002 11664 17008
rect 11624 16658 11652 17002
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11610 16552 11666 16561
rect 11716 16538 11744 16730
rect 11666 16510 11744 16538
rect 11610 16487 11612 16496
rect 11664 16487 11666 16496
rect 11612 16458 11664 16464
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 11532 14890 11560 15370
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 11624 14482 11652 15642
rect 11716 15162 11744 16050
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11520 14272 11572 14278
rect 11518 14240 11520 14249
rect 11572 14240 11574 14249
rect 11518 14175 11574 14184
rect 11334 14104 11390 14113
rect 11624 14090 11652 14418
rect 11334 14039 11390 14048
rect 11440 14062 11652 14090
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 10692 11630 10744 11636
rect 10704 11558 10732 11630
rect 10796 11614 11008 11642
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10232 11144 10284 11150
rect 10230 11112 10232 11121
rect 10324 11144 10376 11150
rect 10284 11112 10286 11121
rect 10324 11086 10376 11092
rect 10230 11047 10286 11056
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10244 9586 10272 9998
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10336 8838 10364 11086
rect 10428 10538 10456 11342
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10520 10266 10548 10610
rect 10598 10432 10654 10441
rect 10598 10367 10654 10376
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10414 10160 10470 10169
rect 10414 10095 10416 10104
rect 10468 10095 10470 10104
rect 10416 10066 10468 10072
rect 10612 9994 10640 10367
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 8634 10456 8774
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10612 8090 10640 9590
rect 10704 9518 10732 11494
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10796 6866 10824 11614
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10966 11520 11022 11529
rect 10888 11082 10916 11494
rect 10966 11455 11022 11464
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10980 11014 11008 11455
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10980 8498 11008 8910
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 11072 6254 11100 11630
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11164 11354 11192 11562
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11242 11112 11298 11121
rect 11242 11047 11298 11056
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10742 11192 10950
rect 11256 10742 11284 11047
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11348 10266 11376 14039
rect 11440 12374 11468 14062
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11532 12986 11560 13806
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11428 11280 11480 11286
rect 11426 11248 11428 11257
rect 11480 11248 11482 11257
rect 11426 11183 11482 11192
rect 11532 10810 11560 12174
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11256 9722 11284 10066
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11164 7818 11192 9590
rect 11532 8974 11560 10610
rect 11624 9178 11652 13942
rect 11704 12640 11756 12646
rect 11702 12608 11704 12617
rect 11756 12608 11758 12617
rect 11702 12543 11758 12552
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11256 8294 11284 8910
rect 11716 8634 11744 12242
rect 11808 11354 11836 18702
rect 11992 17270 12020 22066
rect 12070 21992 12126 22001
rect 12070 21927 12072 21936
rect 12124 21927 12126 21936
rect 12072 21898 12124 21904
rect 12176 21010 12204 33322
rect 13556 31754 13584 33458
rect 13464 31726 13584 31754
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 12256 27328 12308 27334
rect 12256 27270 12308 27276
rect 12268 26382 12296 27270
rect 12636 27033 12664 27406
rect 12622 27024 12678 27033
rect 12622 26959 12624 26968
rect 12676 26959 12678 26968
rect 12624 26930 12676 26936
rect 12440 26852 12492 26858
rect 12440 26794 12492 26800
rect 12256 26376 12308 26382
rect 12452 26330 12480 26794
rect 12256 26318 12308 26324
rect 12360 26302 12480 26330
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12360 26042 12388 26302
rect 12348 26036 12400 26042
rect 12348 25978 12400 25984
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12452 25702 12480 25910
rect 12348 25696 12400 25702
rect 12348 25638 12400 25644
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 12360 24342 12388 25638
rect 12348 24336 12400 24342
rect 12348 24278 12400 24284
rect 12544 23322 12572 26318
rect 12900 26308 12952 26314
rect 12900 26250 12952 26256
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12636 24857 12664 25842
rect 12728 25294 12756 26182
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12622 24848 12678 24857
rect 12622 24783 12678 24792
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12544 22234 12572 23258
rect 12728 22642 12756 24346
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12268 21690 12296 21898
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12360 20806 12388 21966
rect 12820 21554 12848 25774
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12360 20602 12388 20742
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 12084 19310 12112 19994
rect 12728 19689 12756 20402
rect 12714 19680 12770 19689
rect 12714 19615 12770 19624
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18970 12480 19110
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11992 17082 12020 17206
rect 11900 17054 12020 17082
rect 11900 15609 11928 17054
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11992 16794 12020 16934
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11978 16008 12034 16017
rect 11978 15943 11980 15952
rect 12032 15943 12034 15952
rect 11980 15914 12032 15920
rect 11886 15600 11942 15609
rect 11886 15535 11942 15544
rect 11900 13530 11928 15535
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 14113 12020 14214
rect 11978 14104 12034 14113
rect 11978 14039 12034 14048
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11900 12306 11928 12922
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11886 11384 11942 11393
rect 11796 11348 11848 11354
rect 11886 11319 11942 11328
rect 11796 11290 11848 11296
rect 11900 11150 11928 11319
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11900 10810 11928 11086
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11808 10538 11836 10678
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11796 10532 11848 10538
rect 11796 10474 11848 10480
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11808 9178 11836 9998
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11900 8566 11928 10610
rect 11992 9654 12020 13806
rect 12084 11014 12112 15370
rect 12176 15178 12204 17546
rect 12360 16998 12388 18566
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12360 15570 12388 16934
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12176 15150 12388 15178
rect 12176 14482 12204 15150
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12176 14249 12204 14282
rect 12162 14240 12218 14249
rect 12162 14175 12218 14184
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12176 12986 12204 13126
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12176 12753 12204 12786
rect 12162 12744 12218 12753
rect 12162 12679 12218 12688
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12176 9674 12204 12679
rect 12268 10266 12296 15030
rect 12360 14618 12388 15150
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12360 12782 12388 13126
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12348 12640 12400 12646
rect 12346 12608 12348 12617
rect 12400 12608 12402 12617
rect 12346 12543 12402 12552
rect 12452 11762 12480 18906
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12636 17746 12664 18294
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12636 16425 12664 16458
rect 12622 16416 12678 16425
rect 12622 16351 12678 16360
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12530 13968 12586 13977
rect 12530 13903 12532 13912
rect 12584 13903 12586 13912
rect 12532 13874 12584 13880
rect 12636 12918 12664 14486
rect 12728 13870 12756 19615
rect 12912 19009 12940 26250
rect 13004 25362 13032 30194
rect 13360 26784 13412 26790
rect 13360 26726 13412 26732
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 13188 25498 13216 25842
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 12992 25356 13044 25362
rect 12992 25298 13044 25304
rect 13004 24886 13032 25298
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 13096 23186 13124 25094
rect 13372 24886 13400 26726
rect 13464 25106 13492 31726
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13544 26512 13596 26518
rect 13544 26454 13596 26460
rect 13556 25226 13584 26454
rect 13544 25220 13596 25226
rect 13544 25162 13596 25168
rect 13464 25078 13584 25106
rect 13360 24880 13412 24886
rect 13266 24848 13322 24857
rect 13360 24822 13412 24828
rect 13266 24783 13322 24792
rect 13176 23520 13228 23526
rect 13176 23462 13228 23468
rect 13084 23180 13136 23186
rect 13084 23122 13136 23128
rect 13188 23050 13216 23462
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 13004 22438 13032 22714
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 12898 19000 12954 19009
rect 13004 18970 13032 19858
rect 13096 18970 13124 22578
rect 13280 22094 13308 24783
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13464 23866 13492 24006
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13556 23186 13584 25078
rect 13648 24818 13676 26726
rect 14280 26444 14332 26450
rect 14280 26386 14332 26392
rect 14464 26444 14516 26450
rect 14464 26386 14516 26392
rect 13728 26240 13780 26246
rect 13728 26182 13780 26188
rect 13740 25974 13768 26182
rect 13728 25968 13780 25974
rect 13728 25910 13780 25916
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13636 24064 13688 24070
rect 13636 24006 13688 24012
rect 13648 23798 13676 24006
rect 13636 23792 13688 23798
rect 13636 23734 13688 23740
rect 13832 23662 13860 25638
rect 14188 24132 14240 24138
rect 14188 24074 14240 24080
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13924 23730 13952 24006
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13820 23656 13872 23662
rect 14004 23656 14056 23662
rect 13820 23598 13872 23604
rect 13924 23604 14004 23610
rect 13924 23598 14056 23604
rect 13924 23582 14044 23598
rect 13924 23526 13952 23582
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 14108 23186 14136 23462
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 14004 23180 14056 23186
rect 14004 23122 14056 23128
rect 14096 23180 14148 23186
rect 14096 23122 14148 23128
rect 13728 23112 13780 23118
rect 13556 23060 13728 23066
rect 13556 23054 13780 23060
rect 13556 23038 13768 23054
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13188 22066 13308 22094
rect 12898 18935 12954 18944
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12820 17610 12848 18090
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12728 12918 12756 13194
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12346 11656 12402 11665
rect 12346 11591 12402 11600
rect 12360 11150 12388 11591
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12544 9722 12572 12718
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12636 10198 12664 12174
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12084 9654 12204 9674
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 12072 9648 12204 9654
rect 12124 9646 12204 9648
rect 12072 9590 12124 9596
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 7886 11652 8230
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11716 6186 11744 8434
rect 12084 7274 12112 9590
rect 12728 9178 12756 12718
rect 12820 10062 12848 17546
rect 13188 17542 13216 22066
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13268 21480 13320 21486
rect 13372 21457 13400 21490
rect 13268 21422 13320 21428
rect 13358 21448 13414 21457
rect 13280 20262 13308 21422
rect 13358 21383 13414 21392
rect 13372 20641 13400 21383
rect 13358 20632 13414 20641
rect 13358 20567 13414 20576
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13268 19304 13320 19310
rect 13266 19272 13268 19281
rect 13320 19272 13322 19281
rect 13266 19207 13322 19216
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 13096 16697 13124 17138
rect 13082 16688 13138 16697
rect 13082 16623 13138 16632
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13096 15552 13124 16390
rect 13004 15524 13124 15552
rect 13004 15026 13032 15524
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12912 14550 12940 14894
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12912 13530 12940 14350
rect 13004 13938 13032 14962
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12912 12714 12940 13194
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12912 9674 12940 12038
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13004 10810 13032 11086
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13096 10266 13124 14894
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13188 12850 13216 13670
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13188 11898 13216 12650
rect 13280 12442 13308 18770
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13372 18057 13400 18702
rect 13464 18358 13492 22170
rect 13556 22166 13584 23038
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13544 22160 13596 22166
rect 13544 22102 13596 22108
rect 13636 22092 13688 22098
rect 13636 22034 13688 22040
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13556 20942 13584 21830
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 19446 13584 20198
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13648 19310 13676 22034
rect 13740 20262 13768 22510
rect 13832 21962 13860 22646
rect 13820 21956 13872 21962
rect 13820 21898 13872 21904
rect 14016 21554 14044 23122
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13912 21072 13964 21078
rect 13912 21014 13964 21020
rect 13924 20874 13952 21014
rect 13912 20868 13964 20874
rect 13912 20810 13964 20816
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14016 20466 14044 20810
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13740 19514 13768 20198
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13820 18692 13872 18698
rect 13820 18634 13872 18640
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13358 18048 13414 18057
rect 13358 17983 13414 17992
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17134 13492 17478
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13464 15722 13492 17070
rect 13556 15910 13584 17546
rect 13832 16454 13860 18634
rect 14016 17921 14044 20402
rect 14002 17912 14058 17921
rect 14002 17847 14058 17856
rect 14108 17762 14136 22918
rect 14200 21962 14228 24074
rect 14292 22982 14320 26386
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14384 22098 14412 25094
rect 14476 24206 14504 26386
rect 14556 25492 14608 25498
rect 14556 25434 14608 25440
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 14188 21956 14240 21962
rect 14188 21898 14240 21904
rect 14476 21706 14504 24142
rect 14568 23730 14596 25434
rect 14660 24342 14688 29582
rect 15384 29572 15436 29578
rect 15384 29514 15436 29520
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 14740 25696 14792 25702
rect 14740 25638 14792 25644
rect 14648 24336 14700 24342
rect 14648 24278 14700 24284
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 14568 23322 14596 23666
rect 14660 23594 14688 24278
rect 14752 23730 14780 25638
rect 14844 24138 14872 26726
rect 15108 26308 15160 26314
rect 15108 26250 15160 26256
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 15028 24682 15056 25230
rect 15016 24676 15068 24682
rect 15016 24618 15068 24624
rect 14832 24132 14884 24138
rect 14832 24074 14884 24080
rect 14740 23724 14792 23730
rect 14740 23666 14792 23672
rect 14924 23656 14976 23662
rect 14924 23598 14976 23604
rect 14648 23588 14700 23594
rect 14648 23530 14700 23536
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14648 22092 14700 22098
rect 14844 22094 14872 22986
rect 14936 22778 14964 23598
rect 15120 23118 15148 26250
rect 15212 25362 15240 26726
rect 15200 25356 15252 25362
rect 15200 25298 15252 25304
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15304 22438 15332 22646
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 14844 22066 15056 22094
rect 14648 22034 14700 22040
rect 14660 22001 14688 22034
rect 14646 21992 14702 22001
rect 14556 21956 14608 21962
rect 14646 21927 14702 21936
rect 14556 21898 14608 21904
rect 14384 21678 14504 21706
rect 14384 21468 14412 21678
rect 14464 21616 14516 21622
rect 14462 21584 14464 21593
rect 14516 21584 14518 21593
rect 14462 21519 14518 21528
rect 14384 21440 14504 21468
rect 14186 21040 14242 21049
rect 14186 20975 14242 20984
rect 14200 20602 14228 20975
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14292 20534 14320 20878
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14384 19990 14412 20878
rect 14476 20505 14504 21440
rect 14568 21418 14596 21898
rect 14556 21412 14608 21418
rect 14556 21354 14608 21360
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14844 20505 14872 20538
rect 14462 20496 14518 20505
rect 14462 20431 14518 20440
rect 14830 20496 14886 20505
rect 14936 20466 14964 21286
rect 15028 20806 15056 22066
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 15120 20874 15148 21966
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 14830 20431 14886 20440
rect 14924 20460 14976 20466
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14292 19514 14320 19790
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14384 19378 14412 19450
rect 14476 19378 14504 20431
rect 14924 20402 14976 20408
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14568 19360 14596 19790
rect 14648 19372 14700 19378
rect 14568 19332 14648 19360
rect 14568 19258 14596 19332
rect 14648 19314 14700 19320
rect 14016 17734 14136 17762
rect 14476 19230 14596 19258
rect 14016 17134 14044 17734
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 14016 16726 14044 17070
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13740 16046 13768 16186
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13464 15694 13584 15722
rect 13360 14884 13412 14890
rect 13360 14826 13412 14832
rect 13372 14482 13400 14826
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13372 13462 13400 13670
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13280 10062 13308 10406
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 12820 9646 12940 9674
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 8634 12664 8910
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12820 6662 12848 9646
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12912 9178 12940 9522
rect 13372 9450 13400 13194
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13358 8936 13414 8945
rect 13358 8871 13414 8880
rect 13372 8838 13400 8871
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 13464 6322 13492 13466
rect 13556 9382 13584 15694
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13832 14958 13860 15506
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13648 14074 13676 14486
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13648 12102 13676 13806
rect 13740 13394 13768 14758
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11257 13676 12038
rect 13634 11248 13690 11257
rect 13634 11183 13690 11192
rect 13832 9654 13860 14214
rect 13924 11286 13952 15982
rect 14016 11354 14044 15982
rect 14108 14006 14136 17614
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14200 15570 14228 16526
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 15706 14320 15846
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14186 15464 14242 15473
rect 14186 15399 14242 15408
rect 14200 15094 14228 15399
rect 14292 15094 14320 15642
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13910 11112 13966 11121
rect 13910 11047 13966 11056
rect 13924 10674 13952 11047
rect 14108 10810 14136 13806
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13924 9897 13952 10610
rect 14200 10266 14228 14350
rect 14384 13734 14412 16662
rect 14476 14090 14504 19230
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14844 17270 14872 18702
rect 15028 17746 15056 20742
rect 15212 20448 15240 22374
rect 15396 22094 15424 29514
rect 15660 28552 15712 28558
rect 15660 28494 15712 28500
rect 15476 26920 15528 26926
rect 15476 26862 15528 26868
rect 15488 24818 15516 26862
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15580 26382 15608 26726
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15488 22710 15516 23462
rect 15672 22982 15700 28494
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15752 27328 15804 27334
rect 15752 27270 15804 27276
rect 15764 24818 15792 27270
rect 15856 26042 15884 28018
rect 15936 27872 15988 27878
rect 15936 27814 15988 27820
rect 15948 27470 15976 27814
rect 15936 27464 15988 27470
rect 15936 27406 15988 27412
rect 16028 26240 16080 26246
rect 16028 26182 16080 26188
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 15936 25900 15988 25906
rect 15936 25842 15988 25848
rect 15948 24954 15976 25842
rect 16040 25294 16068 26182
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15936 23180 15988 23186
rect 15936 23122 15988 23128
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15948 22094 15976 23122
rect 16132 22098 16160 34478
rect 16500 29850 16528 35022
rect 17052 31482 17080 35634
rect 18156 35290 18184 37198
rect 18144 35284 18196 35290
rect 18144 35226 18196 35232
rect 18248 35222 18276 37198
rect 19352 37126 19380 39200
rect 20640 37210 20668 39200
rect 22572 37262 22600 39200
rect 20720 37256 20772 37262
rect 20640 37204 20720 37210
rect 20640 37198 20772 37204
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 22928 37256 22980 37262
rect 22928 37198 22980 37204
rect 19984 37188 20036 37194
rect 20640 37182 20760 37198
rect 19984 37130 20036 37136
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 18236 35216 18288 35222
rect 18236 35158 18288 35164
rect 17500 35080 17552 35086
rect 17500 35022 17552 35028
rect 17040 31476 17092 31482
rect 17040 31418 17092 31424
rect 16672 31340 16724 31346
rect 16672 31282 16724 31288
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16304 28552 16356 28558
rect 16304 28494 16356 28500
rect 16316 28082 16344 28494
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 16684 27606 16712 31282
rect 17132 30252 17184 30258
rect 17132 30194 17184 30200
rect 17040 29640 17092 29646
rect 17040 29582 17092 29588
rect 16948 27872 17000 27878
rect 16948 27814 17000 27820
rect 16672 27600 16724 27606
rect 16672 27542 16724 27548
rect 16684 27130 16712 27542
rect 16672 27124 16724 27130
rect 16672 27066 16724 27072
rect 16960 26994 16988 27814
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16212 26240 16264 26246
rect 16212 26182 16264 26188
rect 16224 25362 16252 26182
rect 16396 25764 16448 25770
rect 16396 25706 16448 25712
rect 16488 25764 16540 25770
rect 16488 25706 16540 25712
rect 16212 25356 16264 25362
rect 16212 25298 16264 25304
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16316 23089 16344 24142
rect 16302 23080 16358 23089
rect 16302 23015 16358 23024
rect 15396 22066 15608 22094
rect 15948 22066 16068 22094
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15384 20460 15436 20466
rect 15212 20420 15384 20448
rect 15384 20402 15436 20408
rect 15488 20262 15516 20742
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15580 19310 15608 22066
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15672 21010 15700 21422
rect 15856 21049 15884 21490
rect 15842 21040 15898 21049
rect 15660 21004 15712 21010
rect 15842 20975 15898 20984
rect 15660 20946 15712 20952
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15580 18834 15608 19246
rect 15672 19242 15700 20810
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 15660 19236 15712 19242
rect 15660 19178 15712 19184
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15764 18426 15792 19722
rect 15856 19514 15884 19722
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 15304 17678 15332 18158
rect 14924 17672 14976 17678
rect 14922 17640 14924 17649
rect 15292 17672 15344 17678
rect 14976 17640 14978 17649
rect 15292 17614 15344 17620
rect 14922 17575 14978 17584
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 14832 17264 14884 17270
rect 14832 17206 14884 17212
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15396 16794 15424 17070
rect 15488 16794 15516 17138
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14568 15706 14596 15914
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14660 15042 14688 15642
rect 15108 15428 15160 15434
rect 14568 15014 14688 15042
rect 15028 15388 15108 15416
rect 14568 14958 14596 15014
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14568 14278 14596 14554
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14476 14062 14596 14090
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14292 12238 14320 12271
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14292 10674 14320 11562
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11150 14412 11494
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 13910 9888 13966 9897
rect 13910 9823 13966 9832
rect 13924 9654 13952 9823
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 14200 9042 14228 9522
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14476 6866 14504 13806
rect 14568 12918 14596 14062
rect 14660 13734 14688 14418
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 11150 14596 12038
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14568 9926 14596 10610
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14568 8498 14596 9862
rect 14660 9178 14688 13194
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 14752 11529 14780 11562
rect 14738 11520 14794 11529
rect 14738 11455 14794 11464
rect 14738 11112 14794 11121
rect 14738 11047 14794 11056
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14752 7818 14780 11047
rect 14844 10810 14872 14894
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14936 10146 14964 13942
rect 15028 11898 15056 15388
rect 15108 15370 15160 15376
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15120 14618 15148 14758
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15120 13870 15148 14554
rect 15212 14550 15240 16458
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15198 14376 15254 14385
rect 15198 14311 15200 14320
rect 15252 14311 15254 14320
rect 15200 14282 15252 14288
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15212 12714 15240 13330
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 14844 10118 14964 10146
rect 14844 9586 14872 10118
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14936 9722 14964 9998
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 15028 9042 15056 11630
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 15120 8634 15148 12174
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15212 8634 15240 11630
rect 15304 11354 15332 15370
rect 15396 11354 15424 16458
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15488 14550 15516 15506
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15580 13394 15608 17546
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15672 13802 15700 14350
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15672 12918 15700 13194
rect 15764 12986 15792 18158
rect 15948 16590 15976 20742
rect 16040 20602 16068 22066
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16040 20058 16068 20538
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16408 19786 16436 25706
rect 16500 24410 16528 25706
rect 16764 25696 16816 25702
rect 16764 25638 16816 25644
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16488 24404 16540 24410
rect 16488 24346 16540 24352
rect 16592 24138 16620 24686
rect 16684 24206 16712 25230
rect 16776 24818 16804 25638
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16868 24750 16896 25638
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16580 21072 16632 21078
rect 16684 21060 16712 24142
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16776 22574 16804 22986
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 17052 22506 17080 29582
rect 17040 22500 17092 22506
rect 17040 22442 17092 22448
rect 17144 22001 17172 30194
rect 17512 29850 17540 35022
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 17592 33312 17644 33318
rect 17592 33254 17644 33260
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17604 28778 17632 33254
rect 17512 28750 17632 28778
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17236 26450 17264 26862
rect 17224 26444 17276 26450
rect 17224 26386 17276 26392
rect 17130 21992 17186 22001
rect 17130 21927 17186 21936
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 16868 21554 16896 21626
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 17132 21616 17184 21622
rect 17132 21558 17184 21564
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16632 21032 16712 21060
rect 16580 21014 16632 21020
rect 16868 21010 16896 21286
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 16500 19990 16528 20946
rect 16960 20058 16988 21558
rect 17144 21146 17172 21558
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17236 20448 17264 26386
rect 17512 25906 17540 28750
rect 17684 28416 17736 28422
rect 17684 28358 17736 28364
rect 17696 27470 17724 28358
rect 18696 28212 18748 28218
rect 18696 28154 18748 28160
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17592 26512 17644 26518
rect 17592 26454 17644 26460
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17604 24274 17632 26454
rect 17696 26382 17724 26726
rect 18156 26586 18184 26862
rect 18144 26580 18196 26586
rect 18144 26522 18196 26528
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 18156 25498 18184 26522
rect 18708 25838 18736 28154
rect 18800 26450 18828 33798
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19996 33522 20024 37130
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 20076 34672 20128 34678
rect 20076 34614 20128 34620
rect 19984 33516 20036 33522
rect 19984 33458 20036 33464
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18880 26784 18932 26790
rect 18880 26726 18932 26732
rect 18788 26444 18840 26450
rect 18788 26386 18840 26392
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 18144 25492 18196 25498
rect 18144 25434 18196 25440
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17696 24614 17724 24754
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17684 24608 17736 24614
rect 17684 24550 17736 24556
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17408 24132 17460 24138
rect 17408 24074 17460 24080
rect 17420 23730 17448 24074
rect 17788 24070 17816 24550
rect 17880 24274 17908 24686
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17788 23254 17816 24006
rect 17776 23248 17828 23254
rect 17776 23190 17828 23196
rect 17316 23112 17368 23118
rect 17314 23080 17316 23089
rect 17368 23080 17370 23089
rect 17880 23066 17908 24210
rect 17972 24206 18000 25094
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 18144 23520 18196 23526
rect 18248 23474 18276 25230
rect 18420 24812 18472 24818
rect 18524 24800 18552 25638
rect 18892 25362 18920 26726
rect 18880 25356 18932 25362
rect 18880 25298 18932 25304
rect 18984 25294 19012 31758
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 20088 28762 20116 34614
rect 20732 34610 20760 37062
rect 22940 34678 22968 37198
rect 23860 37126 23888 39200
rect 24768 37256 24820 37262
rect 24768 37198 24820 37204
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 24780 34746 24808 37198
rect 25792 37126 25820 39200
rect 27080 37262 27108 39200
rect 27068 37256 27120 37262
rect 27068 37198 27120 37204
rect 27436 37256 27488 37262
rect 27436 37198 27488 37204
rect 25780 37120 25832 37126
rect 25780 37062 25832 37068
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 24768 34740 24820 34746
rect 24768 34682 24820 34688
rect 22928 34672 22980 34678
rect 22928 34614 22980 34620
rect 20720 34604 20772 34610
rect 20720 34546 20772 34552
rect 21272 34604 21324 34610
rect 21272 34546 21324 34552
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 20352 34536 20404 34542
rect 20352 34478 20404 34484
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 19064 28552 19116 28558
rect 19064 28494 19116 28500
rect 18972 25288 19024 25294
rect 18972 25230 19024 25236
rect 18696 24880 18748 24886
rect 18696 24822 18748 24828
rect 18472 24772 18552 24800
rect 18420 24754 18472 24760
rect 18196 23468 18276 23474
rect 18144 23462 18276 23468
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 18156 23446 18276 23462
rect 18248 23186 18276 23446
rect 18340 23186 18368 23462
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18328 23180 18380 23186
rect 18328 23122 18380 23128
rect 17314 23015 17370 23024
rect 17604 23038 17908 23066
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17420 22710 17448 22918
rect 17408 22704 17460 22710
rect 17408 22646 17460 22652
rect 17408 22568 17460 22574
rect 17408 22510 17460 22516
rect 17316 20460 17368 20466
rect 17236 20420 17316 20448
rect 17316 20402 17368 20408
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 17038 19816 17094 19825
rect 16396 19780 16448 19786
rect 17038 19751 17040 19760
rect 16396 19722 16448 19728
rect 17092 19751 17094 19760
rect 17224 19780 17276 19786
rect 17040 19722 17092 19728
rect 17224 19722 17276 19728
rect 16408 19689 16436 19722
rect 16394 19680 16450 19689
rect 16394 19615 16450 19624
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15488 12442 15516 12718
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15488 11898 15516 12378
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15580 9450 15608 12854
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15672 9178 15700 9522
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15488 8498 15516 8774
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10060 2650 10088 5646
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 12636 2514 12664 4558
rect 14292 2650 14320 6734
rect 15764 5914 15792 12242
rect 15856 10266 15884 13330
rect 15948 12374 15976 16118
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 16040 14550 16068 15982
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 16132 14074 16160 19382
rect 17236 18834 17264 19722
rect 17328 19553 17356 20402
rect 17314 19544 17370 19553
rect 17314 19479 17370 19488
rect 17316 19372 17368 19378
rect 17420 19360 17448 22510
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17512 21690 17540 21966
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17368 19332 17448 19360
rect 17316 19314 17368 19320
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16592 18426 16620 18634
rect 16580 18420 16632 18426
rect 16580 18362 16632 18368
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17270 16528 18022
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16684 16998 16712 18634
rect 17328 18358 17356 19314
rect 17604 18442 17632 23038
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17682 20496 17738 20505
rect 17682 20431 17684 20440
rect 17736 20431 17738 20440
rect 17684 20402 17736 20408
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17420 18414 17632 18442
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16396 16720 16448 16726
rect 16396 16662 16448 16668
rect 16408 16182 16436 16662
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16040 13462 16068 13874
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15948 9586 15976 10678
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 16040 8498 16068 13398
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16132 10810 16160 13262
rect 16224 11898 16252 15982
rect 16408 15570 16436 16118
rect 16500 15910 16528 16526
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16592 15706 16620 15982
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16684 15473 16712 16050
rect 16776 15502 16804 18226
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16764 15496 16816 15502
rect 16670 15464 16726 15473
rect 16764 15438 16816 15444
rect 16670 15399 16726 15408
rect 16684 15026 16712 15399
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 12434 16436 14214
rect 16316 12406 16436 12434
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16316 8498 16344 12406
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16408 10266 16436 10610
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16500 9654 16528 12174
rect 16592 10810 16620 14350
rect 16776 13394 16804 15098
rect 16868 14074 16896 18158
rect 17052 17785 17080 18158
rect 17038 17776 17094 17785
rect 17038 17711 17094 17720
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 16960 16561 16988 17614
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17236 16794 17264 17138
rect 17328 17066 17356 17614
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 16946 16552 17002 16561
rect 16946 16487 17002 16496
rect 16960 16454 16988 16487
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 17420 15688 17448 18414
rect 17592 18352 17644 18358
rect 17592 18294 17644 18300
rect 17328 15660 17448 15688
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16776 12442 16804 13330
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16500 8566 16528 8910
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16684 6118 16712 12174
rect 16960 11354 16988 15030
rect 17328 14414 17356 15660
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17328 14006 17356 14350
rect 17420 14346 17448 15370
rect 17604 15162 17632 18294
rect 17696 17066 17724 19790
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17788 17882 17816 19246
rect 17880 18290 17908 22646
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 17972 21894 18000 22578
rect 18052 22568 18104 22574
rect 18052 22510 18104 22516
rect 18064 21962 18092 22510
rect 18432 22098 18460 22578
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 18052 21956 18104 21962
rect 18052 21898 18104 21904
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18156 21457 18184 21490
rect 18142 21448 18198 21457
rect 18142 21383 18198 21392
rect 18156 20466 18184 21383
rect 18340 20777 18368 21898
rect 18432 21486 18460 22034
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18326 20768 18382 20777
rect 18326 20703 18382 20712
rect 18524 20602 18552 24772
rect 18708 24410 18736 24822
rect 18788 24744 18840 24750
rect 18788 24686 18840 24692
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17788 17082 17816 17478
rect 18064 17218 18092 20334
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18144 18148 18196 18154
rect 18144 18090 18196 18096
rect 18156 17542 18184 18090
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 17880 17202 18092 17218
rect 17868 17196 18092 17202
rect 17920 17190 18092 17196
rect 17868 17138 17920 17144
rect 17960 17128 18012 17134
rect 17788 17066 17908 17082
rect 17960 17070 18012 17076
rect 17684 17060 17736 17066
rect 17788 17060 17920 17066
rect 17788 17054 17868 17060
rect 17684 17002 17736 17008
rect 17868 17002 17920 17008
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17696 14498 17724 15982
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17788 14618 17816 15302
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17328 12442 17356 12650
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17132 12232 17184 12238
rect 17130 12200 17132 12209
rect 17316 12232 17368 12238
rect 17184 12200 17186 12209
rect 17316 12174 17368 12180
rect 17130 12135 17186 12144
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16868 9722 16896 10066
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16856 8356 16908 8362
rect 16856 8298 16908 8304
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15488 2650 15516 5646
rect 16776 4622 16804 8298
rect 16868 5234 16896 8298
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16960 2650 16988 11086
rect 17144 11082 17172 11698
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17038 10296 17094 10305
rect 17328 10266 17356 12174
rect 17038 10231 17094 10240
rect 17316 10260 17368 10266
rect 17052 10130 17080 10231
rect 17316 10202 17368 10208
rect 17420 10146 17448 14282
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 10810 17540 12718
rect 17604 11762 17632 14486
rect 17696 14470 17816 14498
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17696 10962 17724 12718
rect 17604 10934 17724 10962
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17328 10118 17448 10146
rect 17328 4146 17356 10118
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17420 9722 17448 9998
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17604 9382 17632 10934
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17696 10062 17724 10542
rect 17788 10198 17816 14470
rect 17880 11898 17908 14894
rect 17972 14074 18000 17070
rect 18064 15450 18092 17190
rect 18156 15978 18184 17478
rect 18248 16522 18276 19994
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18432 19310 18460 19450
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18340 18737 18368 18838
rect 18326 18728 18382 18737
rect 18326 18663 18382 18672
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 18340 16153 18368 16458
rect 18326 16144 18382 16153
rect 18326 16079 18382 16088
rect 18432 16046 18460 19246
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18524 17814 18552 18158
rect 18512 17808 18564 17814
rect 18512 17750 18564 17756
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18064 15422 18276 15450
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17880 10674 17908 11154
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17972 10266 18000 13262
rect 18064 11354 18092 15030
rect 18156 11830 18184 15302
rect 18248 14958 18276 15422
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18340 13938 18368 15642
rect 18418 14784 18474 14793
rect 18418 14719 18474 14728
rect 18432 14482 18460 14719
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18616 14278 18644 22510
rect 18800 22438 18828 24686
rect 18972 24064 19024 24070
rect 18972 24006 19024 24012
rect 18984 23798 19012 24006
rect 18972 23792 19024 23798
rect 18972 23734 19024 23740
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18788 22432 18840 22438
rect 18788 22374 18840 22380
rect 18696 22092 18748 22098
rect 18800 22094 18828 22374
rect 18892 22234 18920 22918
rect 18880 22228 18932 22234
rect 18880 22170 18932 22176
rect 18880 22094 18932 22098
rect 18800 22092 18932 22094
rect 18800 22066 18880 22092
rect 18696 22034 18748 22040
rect 18880 22034 18932 22040
rect 18708 21962 18736 22034
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18984 21622 19012 21830
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 19076 21162 19104 28494
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19340 26240 19392 26246
rect 19340 26182 19392 26188
rect 19352 25906 19380 26182
rect 19444 26042 19472 26862
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 20088 26042 20116 26930
rect 19432 26036 19484 26042
rect 20076 26036 20128 26042
rect 19484 25996 19564 26024
rect 19432 25978 19484 25984
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19536 25838 19564 25996
rect 20076 25978 20128 25984
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 19536 25294 19564 25774
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23662 19472 24006
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23798 20024 24686
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20088 24138 20116 24550
rect 20076 24132 20128 24138
rect 20076 24074 20128 24080
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19260 22778 19288 23054
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19260 22409 19288 22578
rect 19246 22400 19302 22409
rect 19246 22335 19302 22344
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 19352 21486 19380 21966
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 18984 21134 19104 21162
rect 18788 20868 18840 20874
rect 18984 20856 19012 21134
rect 19064 21072 19116 21078
rect 19064 21014 19116 21020
rect 18840 20828 19012 20856
rect 18788 20810 18840 20816
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18708 16658 18736 20402
rect 19076 19514 19104 21014
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19352 20602 19380 20946
rect 19996 20874 20024 21830
rect 20180 21690 20208 21966
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20076 21412 20128 21418
rect 20076 21354 20128 21360
rect 20088 21078 20116 21354
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 20088 20602 20116 20742
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 20180 19854 20208 19926
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18800 16590 18828 19246
rect 19444 18986 19472 19314
rect 19352 18970 19472 18986
rect 19352 18964 19484 18970
rect 19352 18958 19432 18964
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18892 18222 18920 18702
rect 19352 18426 19380 18958
rect 19432 18906 19484 18912
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18800 14550 18828 14826
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18892 14414 18920 16390
rect 18984 15570 19012 16594
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18064 10810 18092 11086
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 9586 17724 9998
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 18248 8974 18276 12854
rect 18340 12782 18368 13126
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18340 12442 18368 12718
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18524 11898 18552 14214
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18616 10266 18644 12174
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18708 11354 18736 11698
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18892 10810 18920 12174
rect 19076 11286 19104 14894
rect 19168 14074 19196 17070
rect 19444 17066 19472 18770
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 18702
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19996 17746 20024 18362
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20088 17202 20116 19654
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 19432 17060 19484 17066
rect 19432 17002 19484 17008
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15162 20116 15642
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 20180 15094 20208 19790
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20272 19378 20300 19654
rect 20364 19378 20392 34478
rect 21284 30326 21312 34546
rect 21272 30320 21324 30326
rect 21272 30262 21324 30268
rect 24688 29850 24716 34546
rect 27172 31822 27200 37062
rect 27448 34746 27476 37198
rect 29012 37126 29040 39200
rect 30300 37210 30328 39200
rect 30380 37256 30432 37262
rect 30300 37204 30380 37210
rect 30300 37198 30432 37204
rect 31588 37210 31616 39200
rect 33520 37262 33548 39200
rect 34808 37262 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 36740 37262 36768 39200
rect 37186 38176 37242 38185
rect 37186 38111 37242 38120
rect 31760 37256 31812 37262
rect 31588 37204 31760 37210
rect 31588 37198 31812 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 36728 37256 36780 37262
rect 36728 37198 36780 37204
rect 29368 37188 29420 37194
rect 30300 37182 30420 37198
rect 31588 37182 31800 37198
rect 33968 37188 34020 37194
rect 29368 37130 29420 37136
rect 33968 37130 34020 37136
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 27436 34740 27488 34746
rect 27436 34682 27488 34688
rect 29380 33522 29408 37130
rect 30472 37120 30524 37126
rect 30472 37062 30524 37068
rect 32312 37120 32364 37126
rect 32312 37062 32364 37068
rect 30288 36916 30340 36922
rect 30288 36858 30340 36864
rect 30300 33998 30328 36858
rect 30288 33992 30340 33998
rect 30288 33934 30340 33940
rect 29368 33516 29420 33522
rect 29368 33458 29420 33464
rect 27160 31816 27212 31822
rect 27160 31758 27212 31764
rect 27252 30048 27304 30054
rect 27252 29990 27304 29996
rect 29184 30048 29236 30054
rect 29184 29990 29236 29996
rect 24676 29844 24728 29850
rect 24676 29786 24728 29792
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20456 23730 20484 26522
rect 20628 26308 20680 26314
rect 20628 26250 20680 26256
rect 20640 26042 20668 26250
rect 20628 26036 20680 26042
rect 20628 25978 20680 25984
rect 20536 25696 20588 25702
rect 20536 25638 20588 25644
rect 20548 24818 20576 25638
rect 20732 24818 20760 27814
rect 20904 25152 20956 25158
rect 20904 25094 20956 25100
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20812 24676 20864 24682
rect 20812 24618 20864 24624
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 20548 23322 20576 23802
rect 20536 23316 20588 23322
rect 20536 23258 20588 23264
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20732 22710 20760 23054
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20824 22574 20852 24618
rect 20916 24274 20944 25094
rect 21088 24744 21140 24750
rect 21088 24686 21140 24692
rect 21100 24274 21128 24686
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19444 14414 19472 14758
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19260 13938 19288 14214
rect 19444 13954 19472 14350
rect 19996 14346 20024 14758
rect 20272 14618 20300 15438
rect 20352 15428 20404 15434
rect 20456 15416 20484 22374
rect 21192 21554 21220 22578
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21284 21078 21312 21898
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21272 21072 21324 21078
rect 21272 21014 21324 21020
rect 21180 20936 21232 20942
rect 21180 20878 21232 20884
rect 21192 20602 21220 20878
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21376 20466 21404 21490
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20732 18086 20760 18566
rect 20824 18290 20852 19654
rect 21008 18970 21036 19790
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20548 15706 20576 17546
rect 20732 17270 20760 18022
rect 20916 17746 20944 18702
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20916 17270 20944 17682
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 21008 16998 21036 18702
rect 21100 18329 21128 20334
rect 21376 19922 21404 20402
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21192 19378 21220 19450
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21086 18320 21142 18329
rect 21086 18255 21142 18264
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20640 16182 20668 16390
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20404 15388 20484 15416
rect 20352 15370 20404 15376
rect 20456 14618 20484 15388
rect 20916 15162 20944 16118
rect 21192 15570 21220 19314
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 18290 21312 19110
rect 21468 18970 21496 22578
rect 21928 22098 21956 23462
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 21824 21956 21876 21962
rect 21824 21898 21876 21904
rect 21836 21690 21864 21898
rect 21824 21684 21876 21690
rect 21824 21626 21876 21632
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21560 18902 21588 21490
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 21928 21010 21956 21422
rect 23400 21078 23428 29582
rect 25412 29504 25464 29510
rect 25412 29446 25464 29452
rect 24032 25900 24084 25906
rect 24032 25842 24084 25848
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23388 21072 23440 21078
rect 23388 21014 23440 21020
rect 21916 21004 21968 21010
rect 21916 20946 21968 20952
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 21548 18896 21600 18902
rect 21548 18838 21600 18844
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21284 17202 21312 17478
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14074 20024 14282
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19248 13932 19300 13938
rect 19444 13926 19564 13954
rect 19248 13874 19300 13880
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18892 10062 18920 10406
rect 19260 10266 19288 12854
rect 19444 12442 19472 13806
rect 19536 13394 19564 13926
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19536 12186 19564 12854
rect 19996 12434 20024 13262
rect 19996 12406 20116 12434
rect 19444 12158 19564 12186
rect 19444 11354 19472 12158
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10810 20024 11086
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19522 10704 19578 10713
rect 19522 10639 19524 10648
rect 19576 10639 19578 10648
rect 19524 10610 19576 10616
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19536 10062 19564 10610
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 20088 6662 20116 12406
rect 20180 11898 20208 13262
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20732 12730 20760 14350
rect 20824 13394 20852 14894
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20640 12594 20668 12718
rect 20732 12702 20852 12730
rect 20640 12566 20760 12594
rect 20732 12442 20760 12566
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20352 12368 20404 12374
rect 20352 12310 20404 12316
rect 20364 12238 20392 12310
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 20272 11150 20300 11562
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20364 8906 20392 12174
rect 20456 11898 20484 12174
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20456 11354 20484 11698
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 20180 5234 20208 8774
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 18616 2446 18644 4422
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20088 2446 20116 4966
rect 20456 2650 20484 9998
rect 20824 6730 20852 12702
rect 20916 11898 20944 12854
rect 21008 12442 21036 13806
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12782 21128 13126
rect 21192 12986 21220 14962
rect 21284 14618 21312 15370
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 21100 11762 21128 12582
rect 21376 12374 21404 18158
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21468 16590 21496 17546
rect 21560 16590 21588 18838
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 21456 15972 21508 15978
rect 21456 15914 21508 15920
rect 21468 15570 21496 15914
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21560 14822 21588 16050
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21468 14278 21496 14554
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 21560 14006 21588 14350
rect 21548 14000 21600 14006
rect 21548 13942 21600 13948
rect 21652 13852 21680 16662
rect 21744 14482 21772 17070
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21560 13824 21680 13852
rect 21836 13841 21864 16934
rect 22020 16522 22048 20402
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22112 19242 22140 19654
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 22204 17338 22232 19314
rect 22296 18222 22324 20198
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22388 17882 22416 18362
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22480 17762 22508 20946
rect 22836 20868 22888 20874
rect 22836 20810 22888 20816
rect 22848 20602 22876 20810
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23584 20602 23612 20742
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23676 20466 23704 21286
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 24044 19922 24072 25842
rect 25424 24342 25452 29446
rect 25412 24336 25464 24342
rect 25412 24278 25464 24284
rect 27264 24206 27292 29990
rect 27252 24200 27304 24206
rect 27252 24142 27304 24148
rect 25320 21548 25372 21554
rect 25320 21490 25372 21496
rect 24584 20392 24636 20398
rect 24584 20334 24636 20340
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 23112 19780 23164 19786
rect 23112 19722 23164 19728
rect 23124 19378 23152 19722
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22664 18290 22692 18566
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 23124 17882 23152 19314
rect 24044 18834 24072 19858
rect 24596 19854 24624 20334
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 24768 19304 24820 19310
rect 24768 19246 24820 19252
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24688 18834 24716 19110
rect 24780 18902 24808 19246
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24768 18896 24820 18902
rect 24768 18838 24820 18844
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23400 18426 23428 18634
rect 24688 18426 24716 18770
rect 24768 18692 24820 18698
rect 24768 18634 24820 18640
rect 24780 18426 24808 18634
rect 24872 18630 24900 19110
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 22388 17746 22508 17762
rect 24780 17746 24808 18022
rect 24964 17882 24992 18226
rect 25056 18154 25084 19246
rect 25240 19242 25268 19654
rect 25228 19236 25280 19242
rect 25228 19178 25280 19184
rect 25332 18834 25360 21490
rect 29000 21344 29052 21350
rect 29000 21286 29052 21292
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25412 19848 25464 19854
rect 25412 19790 25464 19796
rect 25424 18970 25452 19790
rect 25516 19378 25544 20198
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25884 18970 25912 19246
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 25320 18828 25372 18834
rect 25320 18770 25372 18776
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25044 18148 25096 18154
rect 25044 18090 25096 18096
rect 24952 17876 25004 17882
rect 24952 17818 25004 17824
rect 22376 17740 22508 17746
rect 22428 17734 22508 17740
rect 24768 17740 24820 17746
rect 22376 17682 22428 17688
rect 24768 17682 24820 17688
rect 25148 17678 25176 18634
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 22664 17338 22692 17614
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 23584 16794 23612 17614
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23860 16658 23888 17614
rect 25136 17264 25188 17270
rect 25136 17206 25188 17212
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 24136 16794 24164 16934
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 22664 16538 22692 16594
rect 22008 16516 22060 16522
rect 22664 16510 22784 16538
rect 22008 16458 22060 16464
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22664 16250 22692 16390
rect 22756 16250 22784 16510
rect 23768 16250 23796 16594
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 21822 13832 21878 13841
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21560 6866 21588 13824
rect 21822 13767 21878 13776
rect 21928 13734 21956 15982
rect 22204 15706 22232 15982
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22480 15366 22508 15982
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22572 15638 22600 15846
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22664 15450 22692 16186
rect 24308 16040 24360 16046
rect 24360 16000 24440 16028
rect 24308 15982 24360 15988
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 22664 15434 22784 15450
rect 22664 15428 22796 15434
rect 22664 15422 22744 15428
rect 22744 15370 22796 15376
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 23124 14958 23152 15506
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23296 14952 23348 14958
rect 23584 14906 23612 14962
rect 23676 14958 23704 15302
rect 23296 14894 23348 14900
rect 23308 14414 23336 14894
rect 23400 14878 23612 14906
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22388 14074 22416 14214
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22006 13832 22062 13841
rect 22006 13767 22062 13776
rect 21916 13728 21968 13734
rect 21916 13670 21968 13676
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 21652 12238 21680 12854
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21928 10266 21956 13670
rect 22020 12306 22048 13767
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22296 12850 22324 13670
rect 22388 13394 22416 14010
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22480 12986 22508 14350
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22572 13394 22600 13806
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 22664 7274 22692 14350
rect 23400 13530 23428 14878
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23492 13938 23520 14350
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23492 13841 23520 13874
rect 23478 13832 23534 13841
rect 23478 13767 23534 13776
rect 23584 13530 23612 13942
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 22836 13252 22888 13258
rect 22836 13194 22888 13200
rect 22848 12986 22876 13194
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22756 9994 22784 11698
rect 22744 9988 22796 9994
rect 22744 9930 22796 9936
rect 23032 8974 23060 13330
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23124 12374 23152 12718
rect 23400 12434 23428 12718
rect 23308 12406 23428 12434
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23308 11762 23336 12406
rect 23388 12164 23440 12170
rect 23388 12106 23440 12112
rect 23400 11898 23428 12106
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23676 11626 23704 13262
rect 23664 11620 23716 11626
rect 23664 11562 23716 11568
rect 23768 10062 23796 15914
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23860 15162 23888 15302
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 24044 14074 24072 15438
rect 24308 14544 24360 14550
rect 24308 14486 24360 14492
rect 24320 14074 24348 14486
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 23756 10056 23808 10062
rect 23756 9998 23808 10004
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 24412 7546 24440 16000
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 22652 7268 22704 7274
rect 22652 7210 22704 7216
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 23296 5024 23348 5030
rect 23296 4966 23348 4972
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 23308 2446 23336 4966
rect 23400 2650 23428 6734
rect 24504 6662 24532 17070
rect 24596 16794 24624 17070
rect 25148 16794 25176 17206
rect 25332 17134 25360 18770
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 25608 17678 25636 18226
rect 25596 17672 25648 17678
rect 25596 17614 25648 17620
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 25504 17536 25556 17542
rect 25504 17478 25556 17484
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 25136 16788 25188 16794
rect 25136 16730 25188 16736
rect 25516 16658 25544 17478
rect 26160 17202 26188 17614
rect 26252 17338 26280 18226
rect 26620 17882 26648 18702
rect 29012 18358 29040 21286
rect 29196 20058 29224 29990
rect 30484 29646 30512 37062
rect 32324 30190 32352 37062
rect 33232 35488 33284 35494
rect 33232 35430 33284 35436
rect 33244 34610 33272 35430
rect 33232 34604 33284 34610
rect 33232 34546 33284 34552
rect 33140 34536 33192 34542
rect 33140 34478 33192 34484
rect 32312 30184 32364 30190
rect 32312 30126 32364 30132
rect 30472 29640 30524 29646
rect 30472 29582 30524 29588
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 29736 26988 29788 26994
rect 29736 26930 29788 26936
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 29748 19990 29776 26930
rect 30484 22574 30512 29446
rect 33152 26234 33180 34478
rect 33508 33516 33560 33522
rect 33508 33458 33560 33464
rect 33232 32428 33284 32434
rect 33232 32370 33284 32376
rect 33244 27130 33272 32370
rect 33324 30252 33376 30258
rect 33324 30194 33376 30200
rect 33336 28762 33364 30194
rect 33520 30122 33548 33458
rect 33980 32570 34008 37130
rect 34888 37120 34940 37126
rect 34888 37062 34940 37068
rect 35900 37120 35952 37126
rect 35900 37062 35952 37068
rect 34900 36922 34928 37062
rect 34888 36916 34940 36922
rect 34888 36858 34940 36864
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35348 35080 35400 35086
rect 35348 35022 35400 35028
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 33968 32564 34020 32570
rect 33968 32506 34020 32512
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 33784 31952 33836 31958
rect 33784 31894 33836 31900
rect 33508 30116 33560 30122
rect 33508 30058 33560 30064
rect 33324 28756 33376 28762
rect 33324 28698 33376 28704
rect 33324 28552 33376 28558
rect 33324 28494 33376 28500
rect 33232 27124 33284 27130
rect 33232 27066 33284 27072
rect 33152 26206 33272 26234
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 30472 22568 30524 22574
rect 30472 22510 30524 22516
rect 32220 21888 32272 21894
rect 32220 21830 32272 21836
rect 32232 20942 32260 21830
rect 33152 21690 33180 24142
rect 33244 23186 33272 26206
rect 33232 23180 33284 23186
rect 33232 23122 33284 23128
rect 33336 22438 33364 28494
rect 33796 28082 33824 31894
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30938 35388 35022
rect 35348 30932 35400 30938
rect 35348 30874 35400 30880
rect 33876 30728 33928 30734
rect 33876 30670 33928 30676
rect 33784 28076 33836 28082
rect 33784 28018 33836 28024
rect 33888 26042 33916 30670
rect 35912 30326 35940 37062
rect 36728 36576 36780 36582
rect 36728 36518 36780 36524
rect 35900 30320 35952 30326
rect 35900 30262 35952 30268
rect 35440 30048 35492 30054
rect 35440 29990 35492 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35452 28558 35480 29990
rect 36740 29646 36768 36518
rect 37200 36378 37228 38111
rect 37556 36780 37608 36786
rect 37556 36722 37608 36728
rect 37372 36576 37424 36582
rect 37372 36518 37424 36524
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 37384 36174 37412 36518
rect 37372 36168 37424 36174
rect 37372 36110 37424 36116
rect 36728 29640 36780 29646
rect 36728 29582 36780 29588
rect 35440 28552 35492 28558
rect 35440 28494 35492 28500
rect 34060 28416 34112 28422
rect 34060 28358 34112 28364
rect 34072 28218 34100 28358
rect 34060 28212 34112 28218
rect 34060 28154 34112 28160
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35348 26988 35400 26994
rect 35348 26930 35400 26936
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 33876 26036 33928 26042
rect 33876 25978 33928 25984
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34808 23730 34836 25094
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24410 35388 26930
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 36096 25498 36124 26318
rect 36084 25492 36136 25498
rect 36084 25434 36136 25440
rect 35624 25288 35676 25294
rect 35624 25230 35676 25236
rect 35348 24404 35400 24410
rect 35348 24346 35400 24352
rect 34796 23724 34848 23730
rect 34796 23666 34848 23672
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 33324 22432 33376 22438
rect 33324 22374 33376 22380
rect 33140 21684 33192 21690
rect 33140 21626 33192 21632
rect 34532 21554 34560 23462
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34520 21548 34572 21554
rect 34520 21490 34572 21496
rect 35636 21418 35664 25230
rect 37568 24818 37596 36722
rect 38028 35698 38056 39200
rect 38200 37120 38252 37126
rect 38200 37062 38252 37068
rect 38212 36825 38240 37062
rect 39316 36854 39344 39200
rect 39304 36848 39356 36854
rect 38198 36816 38254 36825
rect 39304 36790 39356 36796
rect 38198 36751 38254 36760
rect 38016 35692 38068 35698
rect 38016 35634 38068 35640
rect 38200 34944 38252 34950
rect 38200 34886 38252 34892
rect 38212 34785 38240 34886
rect 38198 34776 38254 34785
rect 38198 34711 38254 34720
rect 38198 33416 38254 33425
rect 38198 33351 38200 33360
rect 38252 33351 38254 33360
rect 38200 33322 38252 33328
rect 38292 31816 38344 31822
rect 38292 31758 38344 31764
rect 38304 31385 38332 31758
rect 38290 31376 38346 31385
rect 38290 31311 38346 31320
rect 38292 30252 38344 30258
rect 38292 30194 38344 30200
rect 38304 30025 38332 30194
rect 38290 30016 38346 30025
rect 38290 29951 38346 29960
rect 38016 29164 38068 29170
rect 38016 29106 38068 29112
rect 38028 26586 38056 29106
rect 38200 29028 38252 29034
rect 38200 28970 38252 28976
rect 38212 28665 38240 28970
rect 38198 28656 38254 28665
rect 38198 28591 38254 28600
rect 38200 26784 38252 26790
rect 38200 26726 38252 26732
rect 38212 26625 38240 26726
rect 38198 26616 38254 26625
rect 38016 26580 38068 26586
rect 38198 26551 38254 26560
rect 38016 26522 38068 26528
rect 38292 25288 38344 25294
rect 38290 25256 38292 25265
rect 38344 25256 38346 25265
rect 38290 25191 38346 25200
rect 37556 24812 37608 24818
rect 37556 24754 37608 24760
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 38304 23225 38332 23666
rect 38290 23216 38346 23225
rect 38290 23151 38346 23160
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38304 21865 38332 21966
rect 38290 21856 38346 21865
rect 38290 21791 38346 21800
rect 35624 21412 35676 21418
rect 35624 21354 35676 21360
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32128 20800 32180 20806
rect 32128 20742 32180 20748
rect 29736 19984 29788 19990
rect 29736 19926 29788 19932
rect 32140 19446 32168 20742
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 38292 19848 38344 19854
rect 38290 19816 38292 19825
rect 38344 19816 38346 19825
rect 38290 19751 38346 19760
rect 35532 19712 35584 19718
rect 35532 19654 35584 19660
rect 32128 19440 32180 19446
rect 32128 19382 32180 19388
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 29000 18352 29052 18358
rect 29000 18294 29052 18300
rect 35544 18290 35572 19654
rect 38292 18760 38344 18766
rect 38292 18702 38344 18708
rect 38304 18465 38332 18702
rect 38290 18456 38346 18465
rect 38290 18391 38346 18400
rect 35532 18284 35584 18290
rect 35532 18226 35584 18232
rect 34244 18080 34296 18086
rect 34244 18022 34296 18028
rect 26608 17876 26660 17882
rect 26608 17818 26660 17824
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 33796 17202 33824 17478
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 33784 17196 33836 17202
rect 33784 17138 33836 17144
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25056 16250 25084 16526
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 26160 16114 26188 17138
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 27172 16590 27200 16934
rect 34256 16726 34284 18022
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 17604 34848 17610
rect 34796 17546 34848 17552
rect 34244 16720 34296 16726
rect 34244 16662 34296 16668
rect 34808 16590 34836 17546
rect 38198 17096 38254 17105
rect 38198 17031 38200 17040
rect 38252 17031 38254 17040
rect 38200 17002 38252 17008
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 38108 16652 38160 16658
rect 38108 16594 38160 16600
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 34796 16584 34848 16590
rect 34796 16526 34848 16532
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 24596 15502 24624 16050
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 38120 15706 38148 16594
rect 38108 15700 38160 15706
rect 38108 15642 38160 15648
rect 27436 15632 27488 15638
rect 27436 15574 27488 15580
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24584 15088 24636 15094
rect 24584 15030 24636 15036
rect 24596 14618 24624 15030
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24780 14278 24808 14962
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 25240 14414 25268 14554
rect 26148 14544 26200 14550
rect 26148 14486 26200 14492
rect 25228 14408 25280 14414
rect 25228 14350 25280 14356
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24780 13462 24808 14214
rect 26160 13530 26188 14486
rect 26148 13524 26200 13530
rect 26148 13466 26200 13472
rect 24768 13456 24820 13462
rect 24768 13398 24820 13404
rect 27448 11762 27476 15574
rect 38292 15496 38344 15502
rect 38292 15438 38344 15444
rect 38304 15065 38332 15438
rect 38290 15056 38346 15065
rect 38290 14991 38346 15000
rect 29276 14816 29328 14822
rect 29276 14758 29328 14764
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27632 12850 27660 14010
rect 29288 13938 29316 14758
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 36912 14408 36964 14414
rect 36912 14350 36964 14356
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 30748 13320 30800 13326
rect 30748 13262 30800 13268
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 28080 12640 28132 12646
rect 28080 12582 28132 12588
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 28092 10674 28120 12582
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30116 10062 30144 10406
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 24492 6656 24544 6662
rect 24492 6598 24544 6604
rect 25424 2650 25452 9998
rect 25596 9988 25648 9994
rect 25596 9930 25648 9936
rect 25504 8832 25556 8838
rect 25504 8774 25556 8780
rect 25516 5234 25544 8774
rect 25608 5234 25636 9930
rect 29736 7404 29788 7410
rect 29736 7346 29788 7352
rect 25504 5228 25556 5234
rect 25504 5170 25556 5176
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 27804 5092 27856 5098
rect 27804 5034 27856 5040
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 27816 2446 27844 5034
rect 29748 2650 29776 7346
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30012 5024 30064 5030
rect 30012 4966 30064 4972
rect 29736 2644 29788 2650
rect 29736 2586 29788 2592
rect 30024 2446 30052 4966
rect 30300 2650 30328 6258
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 30576 2582 30604 6734
rect 30760 3738 30788 13262
rect 31668 12640 31720 12646
rect 31668 12582 31720 12588
rect 30840 12368 30892 12374
rect 30840 12310 30892 12316
rect 30852 8974 30880 12310
rect 31680 11762 31708 12582
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 36924 11898 36952 14350
rect 38200 13728 38252 13734
rect 38198 13696 38200 13705
rect 38252 13696 38254 13705
rect 38198 13631 38254 13640
rect 36912 11892 36964 11898
rect 36912 11834 36964 11840
rect 36820 11824 36872 11830
rect 36820 11766 36872 11772
rect 31668 11756 31720 11762
rect 31668 11698 31720 11704
rect 32864 11552 32916 11558
rect 32864 11494 32916 11500
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 30840 8968 30892 8974
rect 30840 8910 30892 8916
rect 32876 5710 32904 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35360 10674 35388 11494
rect 35348 10668 35400 10674
rect 35348 10610 35400 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33060 7886 33088 8774
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 33048 6792 33100 6798
rect 33048 6734 33100 6740
rect 32864 5704 32916 5710
rect 32864 5646 32916 5652
rect 30748 3732 30800 3738
rect 30748 3674 30800 3680
rect 30564 2576 30616 2582
rect 30564 2518 30616 2524
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 27804 2440 27856 2446
rect 27804 2382 27856 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 3974 1456 4030 1465
rect 3974 1391 4030 1400
rect 4540 800 4568 2382
rect 5828 800 5856 2382
rect 7760 800 7788 2382
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9048 800 9076 2246
rect 10336 800 10364 2382
rect 12268 800 12296 2382
rect 13556 800 13584 2382
rect 15488 800 15516 2382
rect 16776 800 16804 2382
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 18708 800 18736 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2246
rect 21284 800 21312 2382
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 23216 800 23244 2246
rect 24504 800 24532 2382
rect 26436 800 26464 2382
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27724 800 27752 2246
rect 29012 800 29040 2382
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 30944 800 30972 2246
rect 32232 800 32260 2382
rect 33060 2310 33088 6734
rect 34348 2650 34376 7346
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34428 5568 34480 5574
rect 34428 5510 34480 5516
rect 34336 2644 34388 2650
rect 34336 2586 34388 2592
rect 34440 2514 34468 5510
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35636 3194 35664 6734
rect 36832 5710 36860 11766
rect 38292 11756 38344 11762
rect 38292 11698 38344 11704
rect 38304 11665 38332 11698
rect 38290 11656 38346 11665
rect 38290 11591 38346 11600
rect 38200 10464 38252 10470
rect 38200 10406 38252 10412
rect 38212 10305 38240 10406
rect 38198 10296 38254 10305
rect 38198 10231 38254 10240
rect 38016 9920 38068 9926
rect 38016 9862 38068 9868
rect 38028 8974 38056 9862
rect 38108 9580 38160 9586
rect 38108 9522 38160 9528
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38016 7744 38068 7750
rect 38016 7686 38068 7692
rect 38028 5710 38056 7686
rect 38120 7546 38148 9522
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38108 7540 38160 7546
rect 38108 7482 38160 7488
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 38304 6905 38332 7346
rect 38290 6896 38346 6905
rect 38290 6831 38346 6840
rect 36820 5704 36872 5710
rect 36820 5646 36872 5652
rect 38016 5704 38068 5710
rect 38016 5646 38068 5652
rect 37464 5568 37516 5574
rect 38200 5568 38252 5574
rect 37464 5510 37516 5516
rect 38198 5536 38200 5545
rect 38252 5536 38254 5545
rect 37476 5234 37504 5510
rect 38198 5471 38254 5480
rect 37464 5228 37516 5234
rect 37464 5170 37516 5176
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 35624 3188 35676 3194
rect 35624 3130 35676 3136
rect 38028 3058 38056 4966
rect 38292 3528 38344 3534
rect 38290 3496 38292 3505
rect 38344 3496 38346 3505
rect 38290 3431 38346 3440
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 38016 3052 38068 3058
rect 38016 2994 38068 3000
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34428 2508 34480 2514
rect 34428 2450 34480 2456
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 33048 2304 33100 2310
rect 33048 2246 33100 2252
rect 34164 800 34192 2382
rect 35452 800 35480 2382
rect 18 200 74 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 7746 200 7802 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 12254 200 12310 800
rect 13542 200 13598 800
rect 15474 200 15530 800
rect 16762 200 16818 800
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 26422 200 26478 800
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 37292 105 37320 2994
rect 38200 2848 38252 2854
rect 38200 2790 38252 2796
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 37384 800 37412 2246
rect 38212 2145 38240 2790
rect 38660 2372 38712 2378
rect 38660 2314 38712 2320
rect 38198 2136 38254 2145
rect 38198 2071 38254 2080
rect 38672 800 38700 2314
rect 37370 200 37426 800
rect 38658 200 38714 800
rect 37278 96 37334 105
rect 37278 31 37334 40
<< via2 >>
rect 2778 39480 2834 39536
rect 2962 37440 3018 37496
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1582 36116 1584 36136
rect 1584 36116 1636 36136
rect 1636 36116 1638 36136
rect 1582 36080 1638 36116
rect 1674 34040 1730 34096
rect 1582 32680 1638 32736
rect 4250 36624 4306 36680
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 1582 30676 1584 30696
rect 1584 30676 1636 30696
rect 1636 30676 1638 30696
rect 1582 30640 1638 30676
rect 1674 29280 1730 29336
rect 1582 27920 1638 27976
rect 1582 25900 1638 25936
rect 1582 25880 1584 25900
rect 1584 25880 1636 25900
rect 1636 25880 1638 25900
rect 18 17720 74 17776
rect 1674 24556 1676 24576
rect 1676 24556 1728 24576
rect 1728 24556 1730 24576
rect 1674 24520 1730 24556
rect 1582 22480 1638 22536
rect 1674 21120 1730 21176
rect 1858 26288 1914 26344
rect 1950 18128 2006 18184
rect 1582 16360 1638 16416
rect 2042 16224 2098 16280
rect 1950 10920 2006 10976
rect 1766 9460 1768 9480
rect 1768 9460 1820 9480
rect 1820 9460 1822 9480
rect 1766 9424 1822 9460
rect 1582 8200 1638 8256
rect 1674 4800 1730 4856
rect 1950 8608 2006 8664
rect 3054 23588 3110 23624
rect 3054 23568 3056 23588
rect 3056 23568 3108 23588
rect 3108 23568 3110 23588
rect 2778 19760 2834 19816
rect 2778 14456 2834 14512
rect 3330 23432 3386 23488
rect 3054 18692 3110 18728
rect 3054 18672 3056 18692
rect 3056 18672 3108 18692
rect 3108 18672 3110 18692
rect 2318 11772 2320 11792
rect 2320 11772 2372 11792
rect 2372 11772 2374 11792
rect 2318 11736 2374 11772
rect 2686 11192 2742 11248
rect 2870 10512 2926 10568
rect 2686 6860 2742 6896
rect 2686 6840 2688 6860
rect 2688 6840 2740 6860
rect 2740 6840 2742 6860
rect 2778 6160 2834 6216
rect 3422 14456 3478 14512
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 5078 29044 5080 29064
rect 5080 29044 5132 29064
rect 5132 29044 5134 29064
rect 5078 29008 5134 29044
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4066 26308 4122 26344
rect 4066 26288 4068 26308
rect 4068 26288 4120 26308
rect 4120 26288 4122 26308
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4342 23740 4344 23760
rect 4344 23740 4396 23760
rect 4396 23740 4398 23760
rect 4342 23704 4398 23740
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3790 20712 3846 20768
rect 3698 19488 3754 19544
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 3698 14320 3754 14376
rect 3790 13504 3846 13560
rect 3238 9560 3294 9616
rect 3422 8064 3478 8120
rect 3330 6740 3332 6760
rect 3332 6740 3384 6760
rect 3384 6740 3386 6760
rect 3330 6704 3386 6740
rect 4618 17448 4674 17504
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 5262 23296 5318 23352
rect 5170 18944 5226 19000
rect 4986 16904 5042 16960
rect 4710 16088 4766 16144
rect 4618 14456 4674 14512
rect 5446 22072 5502 22128
rect 5354 21140 5410 21176
rect 5354 21120 5356 21140
rect 5356 21120 5408 21140
rect 5408 21120 5410 21140
rect 5354 17584 5410 17640
rect 5354 16632 5410 16688
rect 4894 16088 4950 16144
rect 4894 15544 4950 15600
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4066 12960 4122 13016
rect 4066 12588 4068 12608
rect 4068 12588 4120 12608
rect 4120 12588 4122 12608
rect 4066 12552 4122 12588
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4250 12008 4306 12064
rect 3974 10784 4030 10840
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4710 11328 4766 11384
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4434 7812 4490 7848
rect 4434 7792 4436 7812
rect 4436 7792 4488 7812
rect 4488 7792 4490 7812
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3514 4004 3570 4040
rect 3514 3984 3516 4004
rect 3516 3984 3568 4004
rect 3568 3984 3570 4004
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3514 2760 3570 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5262 15272 5318 15328
rect 5538 18944 5594 19000
rect 5722 24792 5778 24848
rect 5906 23432 5962 23488
rect 7194 36488 7250 36544
rect 5814 22208 5870 22264
rect 5446 11464 5502 11520
rect 5630 10240 5686 10296
rect 5538 9016 5594 9072
rect 5630 8472 5686 8528
rect 6090 17992 6146 18048
rect 6090 12724 6092 12744
rect 6092 12724 6144 12744
rect 6144 12724 6146 12744
rect 6090 12688 6146 12724
rect 5998 11192 6054 11248
rect 6366 17604 6422 17640
rect 6366 17584 6368 17604
rect 6368 17584 6420 17604
rect 6420 17584 6422 17604
rect 6550 15988 6552 16008
rect 6552 15988 6604 16008
rect 6604 15988 6606 16008
rect 6550 15952 6606 15988
rect 6366 14728 6422 14784
rect 6918 20596 6974 20632
rect 6918 20576 6920 20596
rect 6920 20576 6972 20596
rect 6972 20576 6974 20596
rect 7286 20324 7342 20360
rect 7286 20304 7288 20324
rect 7288 20304 7340 20324
rect 7340 20304 7342 20324
rect 7010 17448 7066 17504
rect 6918 15816 6974 15872
rect 6918 13640 6974 13696
rect 6366 9016 6422 9072
rect 6642 10804 6698 10840
rect 6642 10784 6644 10804
rect 6644 10784 6696 10804
rect 6696 10784 6698 10804
rect 7286 15428 7342 15464
rect 7286 15408 7288 15428
rect 7288 15408 7340 15428
rect 7340 15408 7342 15428
rect 6826 11736 6882 11792
rect 7102 9596 7104 9616
rect 7104 9596 7156 9616
rect 7156 9596 7158 9616
rect 7102 9560 7158 9596
rect 7470 11772 7472 11792
rect 7472 11772 7524 11792
rect 7524 11772 7526 11792
rect 7470 11736 7526 11772
rect 7930 22072 7986 22128
rect 7654 19216 7710 19272
rect 7654 18808 7710 18864
rect 8206 22208 8262 22264
rect 8022 20168 8078 20224
rect 8206 18808 8262 18864
rect 8758 23704 8814 23760
rect 8114 18264 8170 18320
rect 8114 17992 8170 18048
rect 7930 15136 7986 15192
rect 7470 8336 7526 8392
rect 7838 11464 7894 11520
rect 7838 11056 7894 11112
rect 8942 22752 8998 22808
rect 8758 20168 8814 20224
rect 8666 19216 8722 19272
rect 9310 22108 9312 22128
rect 9312 22108 9364 22128
rect 9364 22108 9366 22128
rect 9310 22072 9366 22108
rect 9034 19352 9090 19408
rect 8114 16088 8170 16144
rect 8114 10260 8170 10296
rect 8114 10240 8116 10260
rect 8116 10240 8168 10260
rect 8168 10240 8170 10260
rect 8574 16224 8630 16280
rect 8942 17584 8998 17640
rect 8482 15408 8538 15464
rect 8390 13912 8446 13968
rect 8482 13268 8484 13288
rect 8484 13268 8536 13288
rect 8536 13268 8538 13288
rect 8482 13232 8538 13268
rect 8482 11736 8538 11792
rect 8390 11500 8392 11520
rect 8392 11500 8444 11520
rect 8444 11500 8446 11520
rect 8390 11464 8446 11500
rect 8574 11192 8630 11248
rect 8114 9596 8116 9616
rect 8116 9596 8168 9616
rect 8168 9596 8170 9616
rect 8114 9560 8170 9596
rect 8114 8608 8170 8664
rect 9218 19624 9274 19680
rect 9218 17312 9274 17368
rect 10322 24812 10378 24848
rect 10322 24792 10324 24812
rect 10324 24792 10376 24812
rect 10376 24792 10378 24812
rect 9586 22772 9642 22808
rect 9586 22752 9588 22772
rect 9588 22752 9640 22772
rect 9640 22752 9642 22772
rect 9586 22636 9642 22672
rect 9586 22616 9588 22636
rect 9588 22616 9640 22636
rect 9640 22616 9642 22636
rect 9954 23024 10010 23080
rect 9770 22380 9772 22400
rect 9772 22380 9824 22400
rect 9824 22380 9826 22400
rect 9770 22344 9826 22380
rect 10138 21564 10140 21584
rect 10140 21564 10192 21584
rect 10192 21564 10194 21584
rect 10138 21528 10194 21564
rect 11150 24928 11206 24984
rect 9586 20304 9642 20360
rect 9494 19352 9550 19408
rect 9586 19216 9642 19272
rect 9586 19116 9588 19136
rect 9588 19116 9640 19136
rect 9640 19116 9642 19136
rect 9586 19080 9642 19116
rect 9494 18708 9496 18728
rect 9496 18708 9548 18728
rect 9548 18708 9550 18728
rect 9494 18672 9550 18708
rect 9034 15036 9036 15056
rect 9036 15036 9088 15056
rect 9088 15036 9090 15056
rect 9034 15000 9090 15036
rect 8942 10104 8998 10160
rect 9402 15852 9404 15872
rect 9404 15852 9456 15872
rect 9456 15852 9458 15872
rect 9402 15816 9458 15852
rect 10230 20712 10286 20768
rect 9862 20460 9918 20496
rect 9862 20440 9864 20460
rect 9864 20440 9916 20460
rect 9916 20440 9918 20460
rect 9954 19760 10010 19816
rect 9678 16088 9734 16144
rect 10138 18672 10194 18728
rect 9862 15952 9918 16008
rect 10598 19236 10654 19272
rect 10598 19216 10600 19236
rect 10600 19216 10652 19236
rect 10652 19216 10654 19236
rect 10598 18692 10654 18728
rect 10598 18672 10600 18692
rect 10600 18672 10652 18692
rect 10652 18672 10654 18692
rect 9494 13504 9550 13560
rect 8482 8472 8538 8528
rect 8390 8336 8446 8392
rect 9218 7540 9274 7576
rect 9218 7520 9220 7540
rect 9220 7520 9272 7540
rect 9272 7520 9274 7540
rect 9494 11092 9496 11112
rect 9496 11092 9548 11112
rect 9548 11092 9550 11112
rect 9494 11056 9550 11092
rect 10598 17720 10654 17776
rect 10506 17448 10562 17504
rect 10046 12824 10102 12880
rect 9678 10376 9734 10432
rect 9678 10260 9734 10296
rect 9678 10240 9680 10260
rect 9680 10240 9732 10260
rect 9732 10240 9734 10260
rect 9678 9868 9680 9888
rect 9680 9868 9732 9888
rect 9732 9868 9734 9888
rect 9678 9832 9734 9868
rect 10322 15272 10378 15328
rect 10230 14728 10286 14784
rect 10506 15020 10562 15056
rect 10506 15000 10508 15020
rect 10508 15000 10560 15020
rect 10560 15000 10562 15020
rect 10414 13776 10470 13832
rect 10598 14476 10654 14512
rect 10598 14456 10600 14476
rect 10600 14456 10652 14476
rect 10652 14456 10654 14476
rect 11150 18828 11206 18864
rect 11150 18808 11152 18828
rect 11152 18808 11204 18828
rect 11204 18808 11206 18828
rect 10782 13232 10838 13288
rect 11058 14764 11060 14784
rect 11060 14764 11112 14784
rect 11112 14764 11114 14784
rect 11058 14728 11114 14764
rect 11150 12708 11206 12744
rect 11150 12688 11152 12708
rect 11152 12688 11204 12708
rect 11204 12688 11206 12708
rect 11886 19372 11942 19408
rect 11886 19352 11888 19372
rect 11888 19352 11940 19372
rect 11940 19352 11942 19372
rect 11610 16516 11666 16552
rect 11610 16496 11612 16516
rect 11612 16496 11664 16516
rect 11664 16496 11666 16516
rect 11518 14220 11520 14240
rect 11520 14220 11572 14240
rect 11572 14220 11574 14240
rect 11518 14184 11574 14220
rect 11334 14048 11390 14104
rect 10230 11092 10232 11112
rect 10232 11092 10284 11112
rect 10284 11092 10286 11112
rect 10230 11056 10286 11092
rect 10598 10376 10654 10432
rect 10414 10124 10470 10160
rect 10414 10104 10416 10124
rect 10416 10104 10468 10124
rect 10468 10104 10470 10124
rect 10966 11464 11022 11520
rect 11242 11056 11298 11112
rect 11426 11228 11428 11248
rect 11428 11228 11480 11248
rect 11480 11228 11482 11248
rect 11426 11192 11482 11228
rect 11702 12588 11704 12608
rect 11704 12588 11756 12608
rect 11756 12588 11758 12608
rect 11702 12552 11758 12588
rect 12070 21956 12126 21992
rect 12070 21936 12072 21956
rect 12072 21936 12124 21956
rect 12124 21936 12126 21956
rect 12622 26988 12678 27024
rect 12622 26968 12624 26988
rect 12624 26968 12676 26988
rect 12676 26968 12678 26988
rect 12622 24792 12678 24848
rect 12714 19624 12770 19680
rect 11978 15972 12034 16008
rect 11978 15952 11980 15972
rect 11980 15952 12032 15972
rect 12032 15952 12034 15972
rect 11886 15544 11942 15600
rect 11978 14048 12034 14104
rect 11886 11328 11942 11384
rect 12162 14184 12218 14240
rect 12162 12688 12218 12744
rect 12346 12588 12348 12608
rect 12348 12588 12400 12608
rect 12400 12588 12402 12608
rect 12346 12552 12402 12588
rect 12622 16360 12678 16416
rect 12530 13932 12586 13968
rect 12530 13912 12532 13932
rect 12532 13912 12584 13932
rect 12584 13912 12586 13932
rect 13266 24792 13322 24848
rect 12898 18944 12954 19000
rect 12346 11600 12402 11656
rect 13358 21392 13414 21448
rect 13358 20576 13414 20632
rect 13266 19252 13268 19272
rect 13268 19252 13320 19272
rect 13320 19252 13322 19272
rect 13266 19216 13322 19252
rect 13082 16632 13138 16688
rect 13358 17992 13414 18048
rect 14002 17856 14058 17912
rect 14646 21936 14702 21992
rect 14462 21564 14464 21584
rect 14464 21564 14516 21584
rect 14516 21564 14518 21584
rect 14462 21528 14518 21564
rect 14186 20984 14242 21040
rect 14462 20440 14518 20496
rect 14830 20440 14886 20496
rect 13358 8880 13414 8936
rect 13634 11192 13690 11248
rect 14186 15408 14242 15464
rect 13910 11056 13966 11112
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 16302 23024 16358 23080
rect 15842 20984 15898 21040
rect 14922 17620 14924 17640
rect 14924 17620 14976 17640
rect 14976 17620 14978 17640
rect 14922 17584 14978 17620
rect 14278 12280 14334 12336
rect 13910 9832 13966 9888
rect 14738 11464 14794 11520
rect 14738 11056 14794 11112
rect 15198 14340 15254 14376
rect 15198 14320 15200 14340
rect 15200 14320 15252 14340
rect 15252 14320 15254 14340
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 17130 21936 17186 21992
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 17314 23060 17316 23080
rect 17316 23060 17368 23080
rect 17368 23060 17370 23080
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 17314 23024 17370 23060
rect 17038 19780 17094 19816
rect 17038 19760 17040 19780
rect 17040 19760 17092 19780
rect 17092 19760 17094 19780
rect 16394 19624 16450 19680
rect 17314 19488 17370 19544
rect 17682 20460 17738 20496
rect 17682 20440 17684 20460
rect 17684 20440 17736 20460
rect 17736 20440 17738 20460
rect 16670 15408 16726 15464
rect 17038 17720 17094 17776
rect 16946 16496 17002 16552
rect 18142 21392 18198 21448
rect 18326 20712 18382 20768
rect 17130 12180 17132 12200
rect 17132 12180 17184 12200
rect 17184 12180 17186 12200
rect 17130 12144 17186 12180
rect 17038 10240 17094 10296
rect 18326 18672 18382 18728
rect 18326 16088 18382 16144
rect 18418 14728 18474 14784
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19246 22344 19302 22400
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37186 38120 37242 38176
rect 21086 18264 21142 18320
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19522 10668 19578 10704
rect 19522 10648 19524 10668
rect 19524 10648 19576 10668
rect 19576 10648 19578 10668
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 21822 13776 21878 13832
rect 22006 13776 22062 13832
rect 23478 13776 23534 13832
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 38198 36760 38254 36816
rect 38198 34720 38254 34776
rect 38198 33380 38254 33416
rect 38198 33360 38200 33380
rect 38200 33360 38252 33380
rect 38252 33360 38254 33380
rect 38290 31320 38346 31376
rect 38290 29960 38346 30016
rect 38198 28600 38254 28656
rect 38198 26560 38254 26616
rect 38290 25236 38292 25256
rect 38292 25236 38344 25256
rect 38344 25236 38346 25256
rect 38290 25200 38346 25236
rect 38290 23160 38346 23216
rect 38290 21800 38346 21856
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 38290 19796 38292 19816
rect 38292 19796 38344 19816
rect 38344 19796 38346 19816
rect 38290 19760 38346 19796
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 38290 18400 38346 18456
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 38198 17060 38254 17096
rect 38198 17040 38200 17060
rect 38200 17040 38252 17060
rect 38252 17040 38254 17060
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 38290 15000 38346 15056
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 38198 13676 38200 13696
rect 38200 13676 38252 13696
rect 38252 13676 38254 13696
rect 38198 13640 38254 13676
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 3974 1400 4030 1456
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38290 11600 38346 11656
rect 38198 10240 38254 10296
rect 38198 8880 38254 8936
rect 38290 6840 38346 6896
rect 38198 5516 38200 5536
rect 38200 5516 38252 5536
rect 38252 5516 38254 5536
rect 38198 5480 38254 5516
rect 38290 3476 38292 3496
rect 38292 3476 38344 3496
rect 38344 3476 38346 3496
rect 38290 3440 38346 3476
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38198 2080 38254 2136
rect 37278 40 37334 96
<< metal3 >>
rect 200 39538 800 39568
rect 2773 39538 2839 39541
rect 200 39536 2839 39538
rect 200 39480 2778 39536
rect 2834 39480 2839 39536
rect 200 39478 2839 39480
rect 200 39448 800 39478
rect 2773 39475 2839 39478
rect 37181 38178 37247 38181
rect 39200 38178 39800 38208
rect 37181 38176 39800 38178
rect 37181 38120 37186 38176
rect 37242 38120 39800 38176
rect 37181 38118 39800 38120
rect 37181 38115 37247 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 2957 37498 3023 37501
rect 200 37496 3023 37498
rect 200 37440 2962 37496
rect 3018 37440 3023 37496
rect 200 37438 3023 37440
rect 200 37408 800 37438
rect 2957 37435 3023 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 38193 36818 38259 36821
rect 39200 36818 39800 36848
rect 38193 36816 39800 36818
rect 38193 36760 38198 36816
rect 38254 36760 39800 36816
rect 38193 36758 39800 36760
rect 38193 36755 38259 36758
rect 39200 36728 39800 36758
rect 4245 36682 4311 36685
rect 5206 36682 5212 36684
rect 4245 36680 5212 36682
rect 4245 36624 4250 36680
rect 4306 36624 5212 36680
rect 4245 36622 5212 36624
rect 4245 36619 4311 36622
rect 5206 36620 5212 36622
rect 5276 36620 5282 36684
rect 7189 36548 7255 36549
rect 7189 36544 7236 36548
rect 7300 36546 7306 36548
rect 7189 36488 7194 36544
rect 7189 36484 7236 36488
rect 7300 36486 7346 36546
rect 7300 36484 7306 36486
rect 7189 36483 7255 36484
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1577 36138 1643 36141
rect 200 36136 1643 36138
rect 200 36080 1582 36136
rect 1638 36080 1643 36136
rect 200 36078 1643 36080
rect 200 36048 800 36078
rect 1577 36075 1643 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 38193 34778 38259 34781
rect 39200 34778 39800 34808
rect 38193 34776 39800 34778
rect 38193 34720 38198 34776
rect 38254 34720 39800 34776
rect 38193 34718 39800 34720
rect 38193 34715 38259 34718
rect 39200 34688 39800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1669 34098 1735 34101
rect 200 34096 1735 34098
rect 200 34040 1674 34096
rect 1730 34040 1735 34096
rect 200 34038 1735 34040
rect 200 34008 800 34038
rect 1669 34035 1735 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32768
rect 1577 32738 1643 32741
rect 200 32736 1643 32738
rect 200 32680 1582 32736
rect 1638 32680 1643 32736
rect 200 32678 1643 32680
rect 200 32648 800 32678
rect 1577 32675 1643 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 38285 31378 38351 31381
rect 39200 31378 39800 31408
rect 38285 31376 39800 31378
rect 38285 31320 38290 31376
rect 38346 31320 39800 31376
rect 38285 31318 39800 31320
rect 38285 31315 38351 31318
rect 39200 31288 39800 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1577 30698 1643 30701
rect 200 30696 1643 30698
rect 200 30640 1582 30696
rect 1638 30640 1643 30696
rect 200 30638 1643 30640
rect 200 30608 800 30638
rect 1577 30635 1643 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38285 30018 38351 30021
rect 39200 30018 39800 30048
rect 38285 30016 39800 30018
rect 38285 29960 38290 30016
rect 38346 29960 39800 30016
rect 38285 29958 39800 29960
rect 38285 29955 38351 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1669 29338 1735 29341
rect 200 29336 1735 29338
rect 200 29280 1674 29336
rect 1730 29280 1735 29336
rect 200 29278 1735 29280
rect 200 29248 800 29278
rect 1669 29275 1735 29278
rect 5073 29066 5139 29069
rect 9438 29066 9444 29068
rect 5073 29064 9444 29066
rect 5073 29008 5078 29064
rect 5134 29008 9444 29064
rect 5073 29006 9444 29008
rect 5073 29003 5139 29006
rect 9438 29004 9444 29006
rect 9508 29004 9514 29068
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 38193 28658 38259 28661
rect 39200 28658 39800 28688
rect 38193 28656 39800 28658
rect 38193 28600 38198 28656
rect 38254 28600 39800 28656
rect 38193 28598 39800 28600
rect 38193 28595 38259 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 200 27978 800 28008
rect 1577 27978 1643 27981
rect 200 27976 1643 27978
rect 200 27920 1582 27976
rect 1638 27920 1643 27976
rect 200 27918 1643 27920
rect 200 27888 800 27918
rect 1577 27915 1643 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 6494 26964 6500 27028
rect 6564 27026 6570 27028
rect 12617 27026 12683 27029
rect 6564 27024 12683 27026
rect 6564 26968 12622 27024
rect 12678 26968 12683 27024
rect 6564 26966 12683 26968
rect 6564 26964 6570 26966
rect 12617 26963 12683 26966
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 38193 26618 38259 26621
rect 39200 26618 39800 26648
rect 38193 26616 39800 26618
rect 38193 26560 38198 26616
rect 38254 26560 39800 26616
rect 38193 26558 39800 26560
rect 38193 26555 38259 26558
rect 39200 26528 39800 26558
rect 1853 26348 1919 26349
rect 1853 26344 1900 26348
rect 1964 26346 1970 26348
rect 4061 26346 4127 26349
rect 6126 26346 6132 26348
rect 1853 26288 1858 26344
rect 1853 26284 1900 26288
rect 1964 26286 2010 26346
rect 4061 26344 6132 26346
rect 4061 26288 4066 26344
rect 4122 26288 6132 26344
rect 4061 26286 6132 26288
rect 1964 26284 1970 26286
rect 1853 26283 1919 26284
rect 4061 26283 4127 26286
rect 6126 26284 6132 26286
rect 6196 26284 6202 26348
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25938 800 25968
rect 1577 25938 1643 25941
rect 200 25936 1643 25938
rect 200 25880 1582 25936
rect 1638 25880 1643 25936
rect 200 25878 1643 25880
rect 200 25848 800 25878
rect 1577 25875 1643 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 38285 25258 38351 25261
rect 39200 25258 39800 25288
rect 38285 25256 39800 25258
rect 38285 25200 38290 25256
rect 38346 25200 39800 25256
rect 38285 25198 39800 25200
rect 38285 25195 38351 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 8150 24924 8156 24988
rect 8220 24986 8226 24988
rect 11145 24986 11211 24989
rect 8220 24984 11211 24986
rect 8220 24928 11150 24984
rect 11206 24928 11211 24984
rect 8220 24926 11211 24928
rect 8220 24924 8226 24926
rect 11145 24923 11211 24926
rect 5717 24850 5783 24853
rect 7230 24850 7236 24852
rect 5717 24848 7236 24850
rect 5717 24792 5722 24848
rect 5778 24792 7236 24848
rect 5717 24790 7236 24792
rect 5717 24787 5783 24790
rect 7230 24788 7236 24790
rect 7300 24788 7306 24852
rect 10317 24850 10383 24853
rect 12617 24850 12683 24853
rect 13261 24850 13327 24853
rect 10317 24848 13327 24850
rect 10317 24792 10322 24848
rect 10378 24792 12622 24848
rect 12678 24792 13266 24848
rect 13322 24792 13327 24848
rect 10317 24790 13327 24792
rect 10317 24787 10383 24790
rect 12617 24787 12683 24790
rect 13261 24787 13327 24790
rect 200 24578 800 24608
rect 1669 24578 1735 24581
rect 200 24576 1735 24578
rect 200 24520 1674 24576
rect 1730 24520 1735 24576
rect 200 24518 1735 24520
rect 200 24488 800 24518
rect 1669 24515 1735 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4337 23762 4403 23765
rect 8753 23762 8819 23765
rect 4337 23760 8819 23762
rect 4337 23704 4342 23760
rect 4398 23704 8758 23760
rect 8814 23704 8819 23760
rect 4337 23702 8819 23704
rect 4337 23699 4403 23702
rect 8753 23699 8819 23702
rect 3049 23626 3115 23629
rect 7966 23626 7972 23628
rect 3049 23624 7972 23626
rect 3049 23568 3054 23624
rect 3110 23568 7972 23624
rect 3049 23566 7972 23568
rect 3049 23563 3115 23566
rect 7966 23564 7972 23566
rect 8036 23564 8042 23628
rect 3325 23492 3391 23493
rect 3325 23488 3372 23492
rect 3436 23490 3442 23492
rect 5901 23490 5967 23493
rect 3325 23432 3330 23488
rect 3325 23428 3372 23432
rect 3436 23430 3482 23490
rect 4662 23488 5967 23490
rect 4662 23432 5906 23488
rect 5962 23432 5967 23488
rect 4662 23430 5967 23432
rect 3436 23428 3442 23430
rect 3325 23427 3391 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 3182 23156 3188 23220
rect 3252 23218 3258 23220
rect 4662 23218 4722 23430
rect 5901 23427 5967 23430
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 5257 23354 5323 23357
rect 5257 23352 5458 23354
rect 5257 23296 5262 23352
rect 5318 23296 5458 23352
rect 5257 23294 5458 23296
rect 5257 23291 5323 23294
rect 3252 23158 4722 23218
rect 3252 23156 3258 23158
rect 200 22538 800 22568
rect 1577 22538 1643 22541
rect 200 22536 1643 22538
rect 200 22480 1582 22536
rect 1638 22480 1643 22536
rect 200 22478 1643 22480
rect 200 22448 800 22478
rect 1577 22475 1643 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 5398 22133 5458 23294
rect 38285 23218 38351 23221
rect 39200 23218 39800 23248
rect 38285 23216 39800 23218
rect 38285 23160 38290 23216
rect 38346 23160 39800 23216
rect 38285 23158 39800 23160
rect 38285 23155 38351 23158
rect 39200 23128 39800 23158
rect 9949 23082 10015 23085
rect 16297 23082 16363 23085
rect 17309 23082 17375 23085
rect 9949 23080 17375 23082
rect 9949 23024 9954 23080
rect 10010 23024 16302 23080
rect 16358 23024 17314 23080
rect 17370 23024 17375 23080
rect 9949 23022 17375 23024
rect 9949 23019 10015 23022
rect 16297 23019 16363 23022
rect 17309 23019 17375 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 8937 22810 9003 22813
rect 9581 22810 9647 22813
rect 8937 22808 9647 22810
rect 8937 22752 8942 22808
rect 8998 22752 9586 22808
rect 9642 22752 9647 22808
rect 8937 22750 9647 22752
rect 8937 22747 9003 22750
rect 9581 22747 9647 22750
rect 5574 22612 5580 22676
rect 5644 22674 5650 22676
rect 9581 22674 9647 22677
rect 5644 22672 9647 22674
rect 5644 22616 9586 22672
rect 9642 22616 9647 22672
rect 5644 22614 9647 22616
rect 5644 22612 5650 22614
rect 9581 22611 9647 22614
rect 9765 22402 9831 22405
rect 19241 22402 19307 22405
rect 9765 22400 19307 22402
rect 9765 22344 9770 22400
rect 9826 22344 19246 22400
rect 19302 22344 19307 22400
rect 9765 22342 19307 22344
rect 9765 22339 9831 22342
rect 19241 22339 19307 22342
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 5809 22266 5875 22269
rect 8201 22266 8267 22269
rect 5809 22264 8267 22266
rect 5809 22208 5814 22264
rect 5870 22208 8206 22264
rect 8262 22208 8267 22264
rect 5809 22206 8267 22208
rect 5809 22203 5875 22206
rect 8201 22203 8267 22206
rect 5398 22128 5507 22133
rect 5398 22072 5446 22128
rect 5502 22072 5507 22128
rect 5398 22070 5507 22072
rect 5441 22067 5507 22070
rect 7925 22130 7991 22133
rect 9305 22130 9371 22133
rect 7925 22128 9371 22130
rect 7925 22072 7930 22128
rect 7986 22072 9310 22128
rect 9366 22072 9371 22128
rect 7925 22070 9371 22072
rect 7925 22067 7991 22070
rect 9305 22067 9371 22070
rect 12065 21994 12131 21997
rect 14641 21994 14707 21997
rect 17125 21994 17191 21997
rect 12065 21992 17191 21994
rect 12065 21936 12070 21992
rect 12126 21936 14646 21992
rect 14702 21936 17130 21992
rect 17186 21936 17191 21992
rect 12065 21934 17191 21936
rect 12065 21931 12131 21934
rect 14641 21931 14707 21934
rect 17125 21931 17191 21934
rect 38285 21858 38351 21861
rect 39200 21858 39800 21888
rect 38285 21856 39800 21858
rect 38285 21800 38290 21856
rect 38346 21800 39800 21856
rect 38285 21798 39800 21800
rect 38285 21795 38351 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 10133 21586 10199 21589
rect 14457 21586 14523 21589
rect 10133 21584 14523 21586
rect 10133 21528 10138 21584
rect 10194 21528 14462 21584
rect 14518 21528 14523 21584
rect 10133 21526 14523 21528
rect 10133 21523 10199 21526
rect 14457 21523 14523 21526
rect 13353 21450 13419 21453
rect 18137 21450 18203 21453
rect 13353 21448 18203 21450
rect 13353 21392 13358 21448
rect 13414 21392 18142 21448
rect 18198 21392 18203 21448
rect 13353 21390 18203 21392
rect 13353 21387 13419 21390
rect 18137 21387 18203 21390
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1669 21178 1735 21181
rect 5349 21180 5415 21181
rect 5349 21178 5396 21180
rect 200 21176 1735 21178
rect 200 21120 1674 21176
rect 1730 21120 1735 21176
rect 200 21118 1735 21120
rect 5304 21176 5396 21178
rect 5304 21120 5354 21176
rect 5304 21118 5396 21120
rect 200 21088 800 21118
rect 1669 21115 1735 21118
rect 5349 21116 5396 21118
rect 5460 21116 5466 21180
rect 5349 21115 5415 21116
rect 14181 21042 14247 21045
rect 15837 21042 15903 21045
rect 14181 21040 15903 21042
rect 14181 20984 14186 21040
rect 14242 20984 15842 21040
rect 15898 20984 15903 21040
rect 14181 20982 15903 20984
rect 14181 20979 14247 20982
rect 15837 20979 15903 20982
rect 3785 20770 3851 20773
rect 6678 20770 6684 20772
rect 3785 20768 6684 20770
rect 3785 20712 3790 20768
rect 3846 20712 6684 20768
rect 3785 20710 6684 20712
rect 3785 20707 3851 20710
rect 6678 20708 6684 20710
rect 6748 20708 6754 20772
rect 10225 20770 10291 20773
rect 18321 20770 18387 20773
rect 10225 20768 18387 20770
rect 10225 20712 10230 20768
rect 10286 20712 18326 20768
rect 18382 20712 18387 20768
rect 10225 20710 18387 20712
rect 10225 20707 10291 20710
rect 18321 20707 18387 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 6913 20634 6979 20637
rect 13353 20634 13419 20637
rect 6913 20632 13419 20634
rect 6913 20576 6918 20632
rect 6974 20576 13358 20632
rect 13414 20576 13419 20632
rect 6913 20574 13419 20576
rect 6913 20571 6979 20574
rect 13353 20571 13419 20574
rect 9857 20498 9923 20501
rect 14457 20498 14523 20501
rect 9857 20496 14523 20498
rect 9857 20440 9862 20496
rect 9918 20440 14462 20496
rect 14518 20440 14523 20496
rect 9857 20438 14523 20440
rect 9857 20435 9923 20438
rect 14457 20435 14523 20438
rect 14825 20498 14891 20501
rect 17677 20498 17743 20501
rect 14825 20496 17743 20498
rect 14825 20440 14830 20496
rect 14886 20440 17682 20496
rect 17738 20440 17743 20496
rect 14825 20438 17743 20440
rect 14825 20435 14891 20438
rect 17677 20435 17743 20438
rect 7281 20362 7347 20365
rect 9581 20362 9647 20365
rect 7281 20360 9647 20362
rect 7281 20304 7286 20360
rect 7342 20304 9586 20360
rect 9642 20304 9647 20360
rect 7281 20302 9647 20304
rect 7281 20299 7347 20302
rect 9581 20299 9647 20302
rect 8017 20226 8083 20229
rect 8753 20226 8819 20229
rect 8017 20224 8819 20226
rect 8017 20168 8022 20224
rect 8078 20168 8758 20224
rect 8814 20168 8819 20224
rect 8017 20166 8819 20168
rect 8017 20163 8083 20166
rect 8753 20163 8819 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 200 19818 800 19848
rect 2773 19818 2839 19821
rect 200 19816 2839 19818
rect 200 19760 2778 19816
rect 2834 19760 2839 19816
rect 200 19758 2839 19760
rect 200 19728 800 19758
rect 2773 19755 2839 19758
rect 9949 19818 10015 19821
rect 17033 19818 17099 19821
rect 9949 19816 17099 19818
rect 9949 19760 9954 19816
rect 10010 19760 17038 19816
rect 17094 19760 17099 19816
rect 9949 19758 17099 19760
rect 9949 19755 10015 19758
rect 17033 19755 17099 19758
rect 38285 19818 38351 19821
rect 39200 19818 39800 19848
rect 38285 19816 39800 19818
rect 38285 19760 38290 19816
rect 38346 19760 39800 19816
rect 38285 19758 39800 19760
rect 38285 19755 38351 19758
rect 39200 19728 39800 19758
rect 9213 19682 9279 19685
rect 12709 19682 12775 19685
rect 9213 19680 12775 19682
rect 9213 19624 9218 19680
rect 9274 19624 12714 19680
rect 12770 19624 12775 19680
rect 9213 19622 12775 19624
rect 9213 19619 9279 19622
rect 12709 19619 12775 19622
rect 15878 19620 15884 19684
rect 15948 19682 15954 19684
rect 16389 19682 16455 19685
rect 15948 19680 16455 19682
rect 15948 19624 16394 19680
rect 16450 19624 16455 19680
rect 15948 19622 16455 19624
rect 15948 19620 15954 19622
rect 16389 19619 16455 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 3693 19546 3759 19549
rect 17309 19546 17375 19549
rect 3693 19544 17375 19546
rect 3693 19488 3698 19544
rect 3754 19488 17314 19544
rect 17370 19488 17375 19544
rect 3693 19486 17375 19488
rect 3693 19483 3759 19486
rect 17309 19483 17375 19486
rect 9029 19410 9095 19413
rect 9489 19410 9555 19413
rect 9029 19408 9555 19410
rect 9029 19352 9034 19408
rect 9090 19352 9494 19408
rect 9550 19352 9555 19408
rect 9029 19350 9555 19352
rect 9029 19347 9095 19350
rect 9489 19347 9555 19350
rect 11881 19410 11947 19413
rect 12014 19410 12020 19412
rect 11881 19408 12020 19410
rect 11881 19352 11886 19408
rect 11942 19352 12020 19408
rect 11881 19350 12020 19352
rect 11881 19347 11947 19350
rect 12014 19348 12020 19350
rect 12084 19348 12090 19412
rect 7649 19272 7715 19277
rect 7649 19216 7654 19272
rect 7710 19216 7715 19272
rect 7649 19211 7715 19216
rect 8661 19274 8727 19277
rect 9581 19274 9647 19277
rect 8661 19272 9647 19274
rect 8661 19216 8666 19272
rect 8722 19216 9586 19272
rect 9642 19216 9647 19272
rect 8661 19214 9647 19216
rect 8661 19211 8727 19214
rect 9581 19211 9647 19214
rect 10593 19274 10659 19277
rect 13261 19274 13327 19277
rect 10593 19272 13327 19274
rect 10593 19216 10598 19272
rect 10654 19216 13266 19272
rect 13322 19216 13327 19272
rect 10593 19214 13327 19216
rect 10593 19211 10659 19214
rect 13261 19211 13327 19214
rect 7652 19138 7712 19211
rect 9581 19138 9647 19141
rect 7652 19136 9647 19138
rect 7652 19080 9586 19136
rect 9642 19080 9647 19136
rect 7652 19078 9647 19080
rect 9581 19075 9647 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 5165 19002 5231 19005
rect 5533 19002 5599 19005
rect 12893 19002 12959 19005
rect 5165 19000 12959 19002
rect 5165 18944 5170 19000
rect 5226 18944 5538 19000
rect 5594 18944 12898 19000
rect 12954 18944 12959 19000
rect 5165 18942 12959 18944
rect 5165 18939 5231 18942
rect 5533 18939 5599 18942
rect 12893 18939 12959 18942
rect 7649 18866 7715 18869
rect 8201 18866 8267 18869
rect 11145 18866 11211 18869
rect 7649 18864 11211 18866
rect 7649 18808 7654 18864
rect 7710 18808 8206 18864
rect 8262 18808 11150 18864
rect 11206 18808 11211 18864
rect 7649 18806 11211 18808
rect 7649 18803 7715 18806
rect 8201 18803 8267 18806
rect 11145 18803 11211 18806
rect 3049 18730 3115 18733
rect 9489 18732 9555 18733
rect 3182 18730 3188 18732
rect 3049 18728 3188 18730
rect 3049 18672 3054 18728
rect 3110 18672 3188 18728
rect 3049 18670 3188 18672
rect 3049 18667 3115 18670
rect 3182 18668 3188 18670
rect 3252 18668 3258 18732
rect 9438 18730 9444 18732
rect 9398 18670 9444 18730
rect 9508 18728 9555 18732
rect 9550 18672 9555 18728
rect 9438 18668 9444 18670
rect 9508 18668 9555 18672
rect 9489 18667 9555 18668
rect 10133 18730 10199 18733
rect 10593 18730 10659 18733
rect 18321 18730 18387 18733
rect 10133 18728 18387 18730
rect 10133 18672 10138 18728
rect 10194 18672 10598 18728
rect 10654 18672 18326 18728
rect 18382 18672 18387 18728
rect 10133 18670 18387 18672
rect 10133 18667 10199 18670
rect 10593 18667 10659 18670
rect 18321 18667 18387 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 38285 18458 38351 18461
rect 39200 18458 39800 18488
rect 38285 18456 39800 18458
rect 38285 18400 38290 18456
rect 38346 18400 39800 18456
rect 38285 18398 39800 18400
rect 38285 18395 38351 18398
rect 39200 18368 39800 18398
rect 8109 18322 8175 18325
rect 21081 18322 21147 18325
rect 8109 18320 21147 18322
rect 8109 18264 8114 18320
rect 8170 18264 21086 18320
rect 21142 18264 21147 18320
rect 8109 18262 21147 18264
rect 8109 18259 8175 18262
rect 21081 18259 21147 18262
rect 1945 18186 2011 18189
rect 8150 18186 8156 18188
rect 1945 18184 8156 18186
rect 1945 18128 1950 18184
rect 2006 18128 8156 18184
rect 1945 18126 8156 18128
rect 1945 18123 2011 18126
rect 8150 18124 8156 18126
rect 8220 18124 8226 18188
rect 6085 18050 6151 18053
rect 8109 18050 8175 18053
rect 6085 18048 8175 18050
rect 6085 17992 6090 18048
rect 6146 17992 8114 18048
rect 8170 17992 8175 18048
rect 6085 17990 8175 17992
rect 6085 17987 6151 17990
rect 8109 17987 8175 17990
rect 13353 18050 13419 18053
rect 13486 18050 13492 18052
rect 13353 18048 13492 18050
rect 13353 17992 13358 18048
rect 13414 17992 13492 18048
rect 13353 17990 13492 17992
rect 13353 17987 13419 17990
rect 13486 17988 13492 17990
rect 13556 17988 13562 18052
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 13854 17852 13860 17916
rect 13924 17914 13930 17916
rect 13997 17914 14063 17917
rect 13924 17912 14063 17914
rect 13924 17856 14002 17912
rect 14058 17856 14063 17912
rect 13924 17854 14063 17856
rect 13924 17852 13930 17854
rect 13997 17851 14063 17854
rect 13 17778 79 17781
rect 200 17778 800 17808
rect 13 17776 800 17778
rect 13 17720 18 17776
rect 74 17720 800 17776
rect 13 17718 800 17720
rect 13 17715 79 17718
rect 200 17688 800 17718
rect 10593 17778 10659 17781
rect 17033 17778 17099 17781
rect 10593 17776 17099 17778
rect 10593 17720 10598 17776
rect 10654 17720 17038 17776
rect 17094 17720 17099 17776
rect 10593 17718 17099 17720
rect 10593 17715 10659 17718
rect 17033 17715 17099 17718
rect 5349 17642 5415 17645
rect 6361 17642 6427 17645
rect 6494 17642 6500 17644
rect 5349 17640 6500 17642
rect 5349 17584 5354 17640
rect 5410 17584 6366 17640
rect 6422 17584 6500 17640
rect 5349 17582 6500 17584
rect 5349 17579 5415 17582
rect 6361 17579 6427 17582
rect 6494 17580 6500 17582
rect 6564 17580 6570 17644
rect 8150 17580 8156 17644
rect 8220 17642 8226 17644
rect 8937 17642 9003 17645
rect 8220 17640 9003 17642
rect 8220 17584 8942 17640
rect 8998 17584 9003 17640
rect 8220 17582 9003 17584
rect 8220 17580 8226 17582
rect 8937 17579 9003 17582
rect 14917 17642 14983 17645
rect 15142 17642 15148 17644
rect 14917 17640 15148 17642
rect 14917 17584 14922 17640
rect 14978 17584 15148 17640
rect 14917 17582 15148 17584
rect 14917 17579 14983 17582
rect 15142 17580 15148 17582
rect 15212 17580 15218 17644
rect 3918 17444 3924 17508
rect 3988 17506 3994 17508
rect 4613 17506 4679 17509
rect 3988 17504 4679 17506
rect 3988 17448 4618 17504
rect 4674 17448 4679 17504
rect 3988 17446 4679 17448
rect 3988 17444 3994 17446
rect 4613 17443 4679 17446
rect 7005 17506 7071 17509
rect 10501 17506 10567 17509
rect 7005 17504 10567 17506
rect 7005 17448 7010 17504
rect 7066 17448 10506 17504
rect 10562 17448 10567 17504
rect 7005 17446 10567 17448
rect 7005 17443 7071 17446
rect 10501 17443 10567 17446
rect 4616 17370 4676 17443
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 9213 17370 9279 17373
rect 4616 17368 9279 17370
rect 4616 17312 9218 17368
rect 9274 17312 9279 17368
rect 4616 17310 9279 17312
rect 9213 17307 9279 17310
rect 38193 17098 38259 17101
rect 39200 17098 39800 17128
rect 38193 17096 39800 17098
rect 38193 17040 38198 17096
rect 38254 17040 39800 17096
rect 38193 17038 39800 17040
rect 38193 17035 38259 17038
rect 39200 17008 39800 17038
rect 4981 16964 5047 16965
rect 4981 16962 5028 16964
rect 4936 16960 5028 16962
rect 4936 16904 4986 16960
rect 4936 16902 5028 16904
rect 4981 16900 5028 16902
rect 5092 16900 5098 16964
rect 4981 16899 5047 16900
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 5349 16692 5415 16693
rect 13077 16692 13143 16693
rect 5349 16688 5396 16692
rect 5460 16690 5466 16692
rect 5349 16632 5354 16688
rect 5349 16628 5396 16632
rect 5460 16630 5506 16690
rect 13077 16688 13124 16692
rect 13188 16690 13194 16692
rect 13077 16632 13082 16688
rect 5460 16628 5466 16630
rect 13077 16628 13124 16632
rect 13188 16630 13234 16690
rect 13188 16628 13194 16630
rect 5349 16627 5415 16628
rect 13077 16627 13143 16628
rect 11605 16554 11671 16557
rect 16941 16554 17007 16557
rect 11605 16552 17007 16554
rect 11605 16496 11610 16552
rect 11666 16496 16946 16552
rect 17002 16496 17007 16552
rect 11605 16494 17007 16496
rect 11605 16491 11671 16494
rect 16941 16491 17007 16494
rect 200 16418 800 16448
rect 1577 16418 1643 16421
rect 12617 16420 12683 16421
rect 200 16416 1643 16418
rect 200 16360 1582 16416
rect 1638 16360 1643 16416
rect 200 16358 1643 16360
rect 200 16328 800 16358
rect 1577 16355 1643 16358
rect 12566 16356 12572 16420
rect 12636 16418 12683 16420
rect 12636 16416 12728 16418
rect 12678 16360 12728 16416
rect 12636 16358 12728 16360
rect 12636 16356 12683 16358
rect 12617 16355 12683 16356
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 2037 16282 2103 16285
rect 8569 16282 8635 16285
rect 2037 16280 8635 16282
rect 2037 16224 2042 16280
rect 2098 16224 8574 16280
rect 8630 16224 8635 16280
rect 2037 16222 8635 16224
rect 2037 16219 2103 16222
rect 8569 16219 8635 16222
rect 4705 16146 4771 16149
rect 4889 16146 4955 16149
rect 8109 16146 8175 16149
rect 4705 16144 8175 16146
rect 4705 16088 4710 16144
rect 4766 16088 4894 16144
rect 4950 16088 8114 16144
rect 8170 16088 8175 16144
rect 4705 16086 8175 16088
rect 4705 16083 4771 16086
rect 4889 16083 4955 16086
rect 8109 16083 8175 16086
rect 9673 16146 9739 16149
rect 18321 16146 18387 16149
rect 9673 16144 18387 16146
rect 9673 16088 9678 16144
rect 9734 16088 18326 16144
rect 18382 16088 18387 16144
rect 9673 16086 18387 16088
rect 9673 16083 9739 16086
rect 18321 16083 18387 16086
rect 6545 16010 6611 16013
rect 9857 16010 9923 16013
rect 11973 16010 12039 16013
rect 6545 16008 12039 16010
rect 6545 15952 6550 16008
rect 6606 15952 9862 16008
rect 9918 15952 11978 16008
rect 12034 15952 12039 16008
rect 6545 15950 12039 15952
rect 6545 15947 6611 15950
rect 9857 15947 9923 15950
rect 11973 15947 12039 15950
rect 6913 15874 6979 15877
rect 9397 15874 9463 15877
rect 6913 15872 9463 15874
rect 6913 15816 6918 15872
rect 6974 15816 9402 15872
rect 9458 15816 9463 15872
rect 6913 15814 9463 15816
rect 6913 15811 6979 15814
rect 9397 15811 9463 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 4889 15602 4955 15605
rect 11881 15602 11947 15605
rect 4889 15600 11947 15602
rect 4889 15544 4894 15600
rect 4950 15544 11886 15600
rect 11942 15544 11947 15600
rect 4889 15542 11947 15544
rect 4889 15539 4955 15542
rect 11881 15539 11947 15542
rect 7281 15466 7347 15469
rect 8477 15466 8543 15469
rect 7281 15464 8543 15466
rect 7281 15408 7286 15464
rect 7342 15408 8482 15464
rect 8538 15408 8543 15464
rect 7281 15406 8543 15408
rect 7281 15403 7347 15406
rect 8477 15403 8543 15406
rect 14181 15466 14247 15469
rect 16665 15466 16731 15469
rect 14181 15464 16731 15466
rect 14181 15408 14186 15464
rect 14242 15408 16670 15464
rect 16726 15408 16731 15464
rect 14181 15406 16731 15408
rect 14181 15403 14247 15406
rect 16665 15403 16731 15406
rect 5257 15330 5323 15333
rect 10317 15330 10383 15333
rect 5257 15328 10383 15330
rect 5257 15272 5262 15328
rect 5318 15272 10322 15328
rect 10378 15272 10383 15328
rect 5257 15270 10383 15272
rect 5257 15267 5323 15270
rect 10317 15267 10383 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 7925 15196 7991 15197
rect 7925 15192 7972 15196
rect 8036 15194 8042 15196
rect 7925 15136 7930 15192
rect 7925 15132 7972 15136
rect 8036 15134 8082 15194
rect 8036 15132 8042 15134
rect 7925 15131 7991 15132
rect 9029 15058 9095 15061
rect 10501 15058 10567 15061
rect 9029 15056 10567 15058
rect 9029 15000 9034 15056
rect 9090 15000 10506 15056
rect 10562 15000 10567 15056
rect 9029 14998 10567 15000
rect 9029 14995 9095 14998
rect 10501 14995 10567 14998
rect 38285 15058 38351 15061
rect 39200 15058 39800 15088
rect 38285 15056 39800 15058
rect 38285 15000 38290 15056
rect 38346 15000 39800 15056
rect 38285 14998 39800 15000
rect 38285 14995 38351 14998
rect 39200 14968 39800 14998
rect 6361 14786 6427 14789
rect 10225 14786 10291 14789
rect 6361 14784 10291 14786
rect 6361 14728 6366 14784
rect 6422 14728 10230 14784
rect 10286 14728 10291 14784
rect 6361 14726 10291 14728
rect 6361 14723 6427 14726
rect 10225 14723 10291 14726
rect 11053 14786 11119 14789
rect 18413 14786 18479 14789
rect 11053 14784 18479 14786
rect 11053 14728 11058 14784
rect 11114 14728 18418 14784
rect 18474 14728 18479 14784
rect 11053 14726 18479 14728
rect 11053 14723 11119 14726
rect 18413 14723 18479 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 2773 14514 2839 14517
rect 3417 14514 3483 14517
rect 2773 14512 3483 14514
rect 2773 14456 2778 14512
rect 2834 14456 3422 14512
rect 3478 14456 3483 14512
rect 2773 14454 3483 14456
rect 2773 14451 2839 14454
rect 3417 14451 3483 14454
rect 4613 14514 4679 14517
rect 10593 14514 10659 14517
rect 4613 14512 10659 14514
rect 4613 14456 4618 14512
rect 4674 14456 10598 14512
rect 10654 14456 10659 14512
rect 4613 14454 10659 14456
rect 4613 14451 4679 14454
rect 10593 14451 10659 14454
rect 200 14378 800 14408
rect 3693 14378 3759 14381
rect 200 14376 3759 14378
rect 200 14320 3698 14376
rect 3754 14320 3759 14376
rect 200 14318 3759 14320
rect 200 14288 800 14318
rect 3693 14315 3759 14318
rect 15193 14378 15259 14381
rect 15878 14378 15884 14380
rect 15193 14376 15884 14378
rect 15193 14320 15198 14376
rect 15254 14320 15884 14376
rect 15193 14318 15884 14320
rect 15193 14315 15259 14318
rect 15878 14316 15884 14318
rect 15948 14316 15954 14380
rect 11513 14242 11579 14245
rect 12157 14242 12223 14245
rect 11513 14240 12223 14242
rect 11513 14184 11518 14240
rect 11574 14184 12162 14240
rect 12218 14184 12223 14240
rect 11513 14182 12223 14184
rect 11513 14179 11579 14182
rect 12157 14179 12223 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 11329 14106 11395 14109
rect 11973 14106 12039 14109
rect 11329 14104 12039 14106
rect 11329 14048 11334 14104
rect 11390 14048 11978 14104
rect 12034 14048 12039 14104
rect 11329 14046 12039 14048
rect 11329 14043 11395 14046
rect 11973 14043 12039 14046
rect 8385 13970 8451 13973
rect 12525 13970 12591 13973
rect 8385 13968 12591 13970
rect 8385 13912 8390 13968
rect 8446 13912 12530 13968
rect 12586 13912 12591 13968
rect 8385 13910 12591 13912
rect 8385 13907 8451 13910
rect 12525 13907 12591 13910
rect 10409 13834 10475 13837
rect 10542 13834 10548 13836
rect 10409 13832 10548 13834
rect 10409 13776 10414 13832
rect 10470 13776 10548 13832
rect 10409 13774 10548 13776
rect 10409 13771 10475 13774
rect 10542 13772 10548 13774
rect 10612 13772 10618 13836
rect 21817 13834 21883 13837
rect 22001 13834 22067 13837
rect 23473 13834 23539 13837
rect 21817 13832 23539 13834
rect 21817 13776 21822 13832
rect 21878 13776 22006 13832
rect 22062 13776 23478 13832
rect 23534 13776 23539 13832
rect 21817 13774 23539 13776
rect 21817 13771 21883 13774
rect 22001 13771 22067 13774
rect 23473 13771 23539 13774
rect 6126 13636 6132 13700
rect 6196 13698 6202 13700
rect 6913 13698 6979 13701
rect 6196 13696 6979 13698
rect 6196 13640 6918 13696
rect 6974 13640 6979 13696
rect 6196 13638 6979 13640
rect 6196 13636 6202 13638
rect 6913 13635 6979 13638
rect 38193 13698 38259 13701
rect 39200 13698 39800 13728
rect 38193 13696 39800 13698
rect 38193 13640 38198 13696
rect 38254 13640 39800 13696
rect 38193 13638 39800 13640
rect 38193 13635 38259 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 3785 13562 3851 13565
rect 3918 13562 3924 13564
rect 3785 13560 3924 13562
rect 3785 13504 3790 13560
rect 3846 13504 3924 13560
rect 3785 13502 3924 13504
rect 3785 13499 3851 13502
rect 3918 13500 3924 13502
rect 3988 13500 3994 13564
rect 5758 13500 5764 13564
rect 5828 13562 5834 13564
rect 9489 13562 9555 13565
rect 5828 13560 9555 13562
rect 5828 13504 9494 13560
rect 9550 13504 9555 13560
rect 5828 13502 9555 13504
rect 5828 13500 5834 13502
rect 9489 13499 9555 13502
rect 8477 13290 8543 13293
rect 10777 13290 10843 13293
rect 8477 13288 10843 13290
rect 8477 13232 8482 13288
rect 8538 13232 10782 13288
rect 10838 13232 10843 13288
rect 8477 13230 10843 13232
rect 8477 13227 8543 13230
rect 10777 13227 10843 13230
rect 19570 13088 19886 13089
rect 200 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4061 13018 4127 13021
rect 200 13016 4127 13018
rect 200 12960 4066 13016
rect 4122 12960 4127 13016
rect 200 12958 4127 12960
rect 200 12928 800 12958
rect 4061 12955 4127 12958
rect 10041 12884 10107 12885
rect 9990 12882 9996 12884
rect 9950 12822 9996 12882
rect 10060 12880 10107 12884
rect 10102 12824 10107 12880
rect 9990 12820 9996 12822
rect 10060 12820 10107 12824
rect 10041 12819 10107 12820
rect 5574 12684 5580 12748
rect 5644 12746 5650 12748
rect 6085 12746 6151 12749
rect 5644 12744 6151 12746
rect 5644 12688 6090 12744
rect 6146 12688 6151 12744
rect 5644 12686 6151 12688
rect 5644 12684 5650 12686
rect 6085 12683 6151 12686
rect 11145 12746 11211 12749
rect 12157 12746 12223 12749
rect 11145 12744 12223 12746
rect 11145 12688 11150 12744
rect 11206 12688 12162 12744
rect 12218 12688 12223 12744
rect 11145 12686 12223 12688
rect 11145 12683 11211 12686
rect 12157 12683 12223 12686
rect 3918 12548 3924 12612
rect 3988 12610 3994 12612
rect 4061 12610 4127 12613
rect 3988 12608 4127 12610
rect 3988 12552 4066 12608
rect 4122 12552 4127 12608
rect 3988 12550 4127 12552
rect 3988 12548 3994 12550
rect 4061 12547 4127 12550
rect 11697 12610 11763 12613
rect 12341 12610 12407 12613
rect 11697 12608 12407 12610
rect 11697 12552 11702 12608
rect 11758 12552 12346 12608
rect 12402 12552 12407 12608
rect 11697 12550 12407 12552
rect 11697 12547 11763 12550
rect 12341 12547 12407 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 5390 12276 5396 12340
rect 5460 12338 5466 12340
rect 14273 12338 14339 12341
rect 5460 12336 14339 12338
rect 5460 12280 14278 12336
rect 14334 12280 14339 12336
rect 5460 12278 14339 12280
rect 5460 12276 5466 12278
rect 14273 12275 14339 12278
rect 15142 12140 15148 12204
rect 15212 12202 15218 12204
rect 17125 12202 17191 12205
rect 15212 12200 17191 12202
rect 15212 12144 17130 12200
rect 17186 12144 17191 12200
rect 15212 12142 17191 12144
rect 15212 12140 15218 12142
rect 17125 12139 17191 12142
rect 4245 12066 4311 12069
rect 4838 12066 4844 12068
rect 4245 12064 4844 12066
rect 4245 12008 4250 12064
rect 4306 12008 4844 12064
rect 4245 12006 4844 12008
rect 4245 12003 4311 12006
rect 4838 12004 4844 12006
rect 4908 12004 4914 12068
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 2313 11794 2379 11797
rect 6821 11794 6887 11797
rect 2313 11792 6887 11794
rect 2313 11736 2318 11792
rect 2374 11736 6826 11792
rect 6882 11736 6887 11792
rect 2313 11734 6887 11736
rect 2313 11731 2379 11734
rect 6821 11731 6887 11734
rect 7465 11794 7531 11797
rect 8477 11794 8543 11797
rect 7465 11792 8543 11794
rect 7465 11736 7470 11792
rect 7526 11736 8482 11792
rect 8538 11736 8543 11792
rect 7465 11734 8543 11736
rect 7465 11731 7531 11734
rect 8477 11731 8543 11734
rect 1894 11596 1900 11660
rect 1964 11658 1970 11660
rect 12341 11658 12407 11661
rect 1964 11656 12407 11658
rect 1964 11600 12346 11656
rect 12402 11600 12407 11656
rect 1964 11598 12407 11600
rect 1964 11596 1970 11598
rect 12341 11595 12407 11598
rect 38285 11658 38351 11661
rect 39200 11658 39800 11688
rect 38285 11656 39800 11658
rect 38285 11600 38290 11656
rect 38346 11600 39800 11656
rect 38285 11598 39800 11600
rect 38285 11595 38351 11598
rect 39200 11568 39800 11598
rect 5022 11460 5028 11524
rect 5092 11522 5098 11524
rect 5441 11522 5507 11525
rect 5092 11520 5507 11522
rect 5092 11464 5446 11520
rect 5502 11464 5507 11520
rect 5092 11462 5507 11464
rect 5092 11460 5098 11462
rect 5441 11459 5507 11462
rect 7833 11522 7899 11525
rect 8385 11522 8451 11525
rect 7833 11520 8451 11522
rect 7833 11464 7838 11520
rect 7894 11464 8390 11520
rect 8446 11464 8451 11520
rect 7833 11462 8451 11464
rect 7833 11459 7899 11462
rect 8385 11459 8451 11462
rect 10961 11522 11027 11525
rect 14733 11522 14799 11525
rect 10961 11520 14799 11522
rect 10961 11464 10966 11520
rect 11022 11464 14738 11520
rect 14794 11464 14799 11520
rect 10961 11462 14799 11464
rect 10961 11459 11027 11462
rect 14733 11459 14799 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 4705 11386 4771 11389
rect 11881 11386 11947 11389
rect 4705 11384 11947 11386
rect 4705 11328 4710 11384
rect 4766 11328 11886 11384
rect 11942 11328 11947 11384
rect 4705 11326 11947 11328
rect 4705 11323 4771 11326
rect 11881 11323 11947 11326
rect 2681 11250 2747 11253
rect 3366 11250 3372 11252
rect 2681 11248 3372 11250
rect 2681 11192 2686 11248
rect 2742 11192 3372 11248
rect 2681 11190 3372 11192
rect 2681 11187 2747 11190
rect 3366 11188 3372 11190
rect 3436 11188 3442 11252
rect 5993 11250 6059 11253
rect 8569 11250 8635 11253
rect 5993 11248 8635 11250
rect 5993 11192 5998 11248
rect 6054 11192 8574 11248
rect 8630 11192 8635 11248
rect 5993 11190 8635 11192
rect 5993 11187 6059 11190
rect 8569 11187 8635 11190
rect 11421 11250 11487 11253
rect 13629 11250 13695 11253
rect 11421 11248 13695 11250
rect 11421 11192 11426 11248
rect 11482 11192 13634 11248
rect 13690 11192 13695 11248
rect 11421 11190 13695 11192
rect 11421 11187 11487 11190
rect 13629 11187 13695 11190
rect 7833 11114 7899 11117
rect 8150 11114 8156 11116
rect 7833 11112 8156 11114
rect 7833 11056 7838 11112
rect 7894 11056 8156 11112
rect 7833 11054 8156 11056
rect 7833 11051 7899 11054
rect 8150 11052 8156 11054
rect 8220 11052 8226 11116
rect 9489 11112 9555 11117
rect 9489 11056 9494 11112
rect 9550 11056 9555 11112
rect 9489 11051 9555 11056
rect 10225 11114 10291 11117
rect 11237 11114 11303 11117
rect 13905 11116 13971 11117
rect 10225 11112 11303 11114
rect 10225 11056 10230 11112
rect 10286 11056 11242 11112
rect 11298 11056 11303 11112
rect 10225 11054 11303 11056
rect 10225 11051 10291 11054
rect 11237 11051 11303 11054
rect 13854 11052 13860 11116
rect 13924 11114 13971 11116
rect 14733 11114 14799 11117
rect 15142 11114 15148 11116
rect 13924 11112 14016 11114
rect 13966 11056 14016 11112
rect 13924 11054 14016 11056
rect 14733 11112 15148 11114
rect 14733 11056 14738 11112
rect 14794 11056 15148 11112
rect 14733 11054 15148 11056
rect 13924 11052 13971 11054
rect 13905 11051 13971 11052
rect 14733 11051 14799 11054
rect 15142 11052 15148 11054
rect 15212 11052 15218 11116
rect 200 10978 800 11008
rect 1945 10978 2011 10981
rect 5574 10978 5580 10980
rect 200 10918 1410 10978
rect 200 10888 800 10918
rect 1350 10570 1410 10918
rect 1945 10976 5580 10978
rect 1945 10920 1950 10976
rect 2006 10920 5580 10976
rect 1945 10918 5580 10920
rect 1945 10915 2011 10918
rect 5574 10916 5580 10918
rect 5644 10916 5650 10980
rect 9492 10978 9552 11051
rect 6364 10918 9552 10978
rect 3969 10844 4035 10845
rect 3918 10780 3924 10844
rect 3988 10842 4035 10844
rect 6364 10842 6424 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 6637 10844 6703 10845
rect 6637 10842 6684 10844
rect 3988 10840 6424 10842
rect 4030 10784 6424 10840
rect 3988 10782 6424 10784
rect 6592 10840 6684 10842
rect 6592 10784 6642 10840
rect 6592 10782 6684 10784
rect 3988 10780 4035 10782
rect 3969 10779 4035 10780
rect 6637 10780 6684 10782
rect 6748 10780 6754 10844
rect 6637 10779 6703 10780
rect 3918 10644 3924 10708
rect 3988 10706 3994 10708
rect 4838 10706 4844 10708
rect 3988 10646 4844 10706
rect 3988 10644 3994 10646
rect 4838 10644 4844 10646
rect 4908 10706 4914 10708
rect 19517 10706 19583 10709
rect 4908 10704 19583 10706
rect 4908 10648 19522 10704
rect 19578 10648 19583 10704
rect 4908 10646 19583 10648
rect 4908 10644 4914 10646
rect 19517 10643 19583 10646
rect 2865 10570 2931 10573
rect 1350 10568 2931 10570
rect 1350 10512 2870 10568
rect 2926 10512 2931 10568
rect 1350 10510 2931 10512
rect 2865 10507 2931 10510
rect 9673 10434 9739 10437
rect 10593 10434 10659 10437
rect 9673 10432 10659 10434
rect 9673 10376 9678 10432
rect 9734 10376 10598 10432
rect 10654 10376 10659 10432
rect 9673 10374 10659 10376
rect 9673 10371 9739 10374
rect 10593 10371 10659 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 5625 10298 5691 10301
rect 8109 10298 8175 10301
rect 5625 10296 8175 10298
rect 5625 10240 5630 10296
rect 5686 10240 8114 10296
rect 8170 10240 8175 10296
rect 5625 10238 8175 10240
rect 5625 10235 5691 10238
rect 8109 10235 8175 10238
rect 9673 10298 9739 10301
rect 17033 10298 17099 10301
rect 9673 10296 17099 10298
rect 9673 10240 9678 10296
rect 9734 10240 17038 10296
rect 17094 10240 17099 10296
rect 9673 10238 17099 10240
rect 9673 10235 9739 10238
rect 17033 10235 17099 10238
rect 38193 10298 38259 10301
rect 39200 10298 39800 10328
rect 38193 10296 39800 10298
rect 38193 10240 38198 10296
rect 38254 10240 39800 10296
rect 38193 10238 39800 10240
rect 38193 10235 38259 10238
rect 39200 10208 39800 10238
rect 8937 10162 9003 10165
rect 10409 10162 10475 10165
rect 8937 10160 10475 10162
rect 8937 10104 8942 10160
rect 8998 10104 10414 10160
rect 10470 10104 10475 10160
rect 8937 10102 10475 10104
rect 8937 10099 9003 10102
rect 10409 10099 10475 10102
rect 9673 9890 9739 9893
rect 13905 9890 13971 9893
rect 9673 9888 13971 9890
rect 9673 9832 9678 9888
rect 9734 9832 13910 9888
rect 13966 9832 13971 9888
rect 9673 9830 13971 9832
rect 9673 9827 9739 9830
rect 13905 9827 13971 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9648
rect 3233 9618 3299 9621
rect 200 9616 3299 9618
rect 200 9560 3238 9616
rect 3294 9560 3299 9616
rect 200 9558 3299 9560
rect 200 9528 800 9558
rect 3233 9555 3299 9558
rect 7097 9618 7163 9621
rect 8109 9618 8175 9621
rect 7097 9616 8175 9618
rect 7097 9560 7102 9616
rect 7158 9560 8114 9616
rect 8170 9560 8175 9616
rect 7097 9558 8175 9560
rect 7097 9555 7163 9558
rect 8109 9555 8175 9558
rect 1761 9482 1827 9485
rect 5758 9482 5764 9484
rect 1761 9480 5764 9482
rect 1761 9424 1766 9480
rect 1822 9424 5764 9480
rect 1761 9422 5764 9424
rect 1761 9419 1827 9422
rect 5758 9420 5764 9422
rect 5828 9420 5834 9484
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 5533 9074 5599 9077
rect 6361 9074 6427 9077
rect 5533 9072 6427 9074
rect 5533 9016 5538 9072
rect 5594 9016 6366 9072
rect 6422 9016 6427 9072
rect 5533 9014 6427 9016
rect 5533 9011 5599 9014
rect 6361 9011 6427 9014
rect 13353 8938 13419 8941
rect 13486 8938 13492 8940
rect 13353 8936 13492 8938
rect 13353 8880 13358 8936
rect 13414 8880 13492 8936
rect 13353 8878 13492 8880
rect 13353 8875 13419 8878
rect 13486 8876 13492 8878
rect 13556 8876 13562 8940
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 1945 8666 2011 8669
rect 8109 8666 8175 8669
rect 1945 8664 8175 8666
rect 1945 8608 1950 8664
rect 2006 8608 8114 8664
rect 8170 8608 8175 8664
rect 1945 8606 8175 8608
rect 1945 8603 2011 8606
rect 8109 8603 8175 8606
rect 5625 8530 5691 8533
rect 8477 8530 8543 8533
rect 5625 8528 8543 8530
rect 5625 8472 5630 8528
rect 5686 8472 8482 8528
rect 8538 8472 8543 8528
rect 5625 8470 8543 8472
rect 5625 8467 5691 8470
rect 8477 8467 8543 8470
rect 7465 8394 7531 8397
rect 8385 8394 8451 8397
rect 7465 8392 8451 8394
rect 7465 8336 7470 8392
rect 7526 8336 8390 8392
rect 8446 8336 8451 8392
rect 7465 8334 8451 8336
rect 7465 8331 7531 8334
rect 8385 8331 8451 8334
rect 200 8258 800 8288
rect 1577 8258 1643 8261
rect 200 8256 1643 8258
rect 200 8200 1582 8256
rect 1638 8200 1643 8256
rect 200 8198 1643 8200
rect 200 8168 800 8198
rect 1577 8195 1643 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 3417 8122 3483 8125
rect 3918 8122 3924 8124
rect 3417 8120 3924 8122
rect 3417 8064 3422 8120
rect 3478 8064 3924 8120
rect 3417 8062 3924 8064
rect 3417 8059 3483 8062
rect 3918 8060 3924 8062
rect 3988 8060 3994 8124
rect 4429 7850 4495 7853
rect 13118 7850 13124 7852
rect 4429 7848 13124 7850
rect 4429 7792 4434 7848
rect 4490 7792 13124 7848
rect 4429 7790 13124 7792
rect 4429 7787 4495 7790
rect 13118 7788 13124 7790
rect 13188 7788 13194 7852
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 9213 7578 9279 7581
rect 12014 7578 12020 7580
rect 9213 7576 12020 7578
rect 9213 7520 9218 7576
rect 9274 7520 12020 7576
rect 9213 7518 12020 7520
rect 9213 7515 9279 7518
rect 12014 7516 12020 7518
rect 12084 7516 12090 7580
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 2681 6898 2747 6901
rect 10542 6898 10548 6900
rect 2681 6896 10548 6898
rect 2681 6840 2686 6896
rect 2742 6840 10548 6896
rect 2681 6838 10548 6840
rect 2681 6835 2747 6838
rect 10542 6836 10548 6838
rect 10612 6836 10618 6900
rect 38285 6898 38351 6901
rect 39200 6898 39800 6928
rect 38285 6896 39800 6898
rect 38285 6840 38290 6896
rect 38346 6840 39800 6896
rect 38285 6838 39800 6840
rect 38285 6835 38351 6838
rect 39200 6808 39800 6838
rect 3325 6762 3391 6765
rect 12566 6762 12572 6764
rect 3325 6760 12572 6762
rect 3325 6704 3330 6760
rect 3386 6704 12572 6760
rect 3325 6702 12572 6704
rect 3325 6699 3391 6702
rect 12566 6700 12572 6702
rect 12636 6700 12642 6764
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 200 6218 800 6248
rect 2773 6218 2839 6221
rect 200 6216 2839 6218
rect 200 6160 2778 6216
rect 2834 6160 2839 6216
rect 200 6158 2839 6160
rect 200 6128 800 6158
rect 2773 6155 2839 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1669 4858 1735 4861
rect 200 4856 1735 4858
rect 200 4800 1674 4856
rect 1730 4800 1735 4856
rect 200 4798 1735 4800
rect 200 4768 800 4798
rect 1669 4795 1735 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 3509 4042 3575 4045
rect 9990 4042 9996 4044
rect 3509 4040 9996 4042
rect 3509 3984 3514 4040
rect 3570 3984 9996 4040
rect 3509 3982 9996 3984
rect 3509 3979 3575 3982
rect 9990 3980 9996 3982
rect 10060 3980 10066 4044
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 38285 3498 38351 3501
rect 39200 3498 39800 3528
rect 38285 3496 39800 3498
rect 38285 3440 38290 3496
rect 38346 3440 39800 3496
rect 38285 3438 39800 3440
rect 38285 3435 38351 3438
rect 39200 3408 39800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 200 2818 800 2848
rect 3509 2818 3575 2821
rect 200 2816 3575 2818
rect 200 2760 3514 2816
rect 3570 2760 3575 2816
rect 200 2758 3575 2760
rect 200 2728 800 2758
rect 3509 2755 3575 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 38193 2138 38259 2141
rect 39200 2138 39800 2168
rect 38193 2136 39800 2138
rect 38193 2080 38198 2136
rect 38254 2080 39800 2136
rect 38193 2078 39800 2080
rect 38193 2075 38259 2078
rect 39200 2048 39800 2078
rect 200 1458 800 1488
rect 3969 1458 4035 1461
rect 200 1456 4035 1458
rect 200 1400 3974 1456
rect 4030 1400 4035 1456
rect 200 1398 4035 1400
rect 200 1368 800 1398
rect 3969 1395 4035 1398
rect 37273 98 37339 101
rect 39200 98 39800 128
rect 37273 96 39800 98
rect 37273 40 37278 96
rect 37334 40 39800 96
rect 37273 38 39800 40
rect 37273 35 37339 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 5212 36620 5276 36684
rect 7236 36544 7300 36548
rect 7236 36488 7250 36544
rect 7250 36488 7300 36544
rect 7236 36484 7300 36488
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 9444 29004 9508 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 6500 26964 6564 27028
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 1900 26344 1964 26348
rect 1900 26288 1914 26344
rect 1914 26288 1964 26344
rect 1900 26284 1964 26288
rect 6132 26284 6196 26348
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 8156 24924 8220 24988
rect 7236 24788 7300 24852
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 7972 23564 8036 23628
rect 3372 23488 3436 23492
rect 3372 23432 3386 23488
rect 3386 23432 3436 23488
rect 3372 23428 3436 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 3188 23156 3252 23220
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 5580 22612 5644 22676
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 5396 21176 5460 21180
rect 5396 21120 5410 21176
rect 5410 21120 5460 21176
rect 5396 21116 5460 21120
rect 6684 20708 6748 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 15884 19620 15948 19684
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 12020 19348 12084 19412
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 3188 18668 3252 18732
rect 9444 18728 9508 18732
rect 9444 18672 9494 18728
rect 9494 18672 9508 18728
rect 9444 18668 9508 18672
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 8156 18124 8220 18188
rect 13492 17988 13556 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 13860 17852 13924 17916
rect 6500 17580 6564 17644
rect 8156 17580 8220 17644
rect 15148 17580 15212 17644
rect 3924 17444 3988 17508
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 5028 16960 5092 16964
rect 5028 16904 5042 16960
rect 5042 16904 5092 16960
rect 5028 16900 5092 16904
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 5396 16688 5460 16692
rect 5396 16632 5410 16688
rect 5410 16632 5460 16688
rect 5396 16628 5460 16632
rect 13124 16688 13188 16692
rect 13124 16632 13138 16688
rect 13138 16632 13188 16688
rect 13124 16628 13188 16632
rect 12572 16416 12636 16420
rect 12572 16360 12622 16416
rect 12622 16360 12636 16416
rect 12572 16356 12636 16360
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 7972 15192 8036 15196
rect 7972 15136 7986 15192
rect 7986 15136 8036 15192
rect 7972 15132 8036 15136
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 15884 14316 15948 14380
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 10548 13772 10612 13836
rect 6132 13636 6196 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 3924 13500 3988 13564
rect 5764 13500 5828 13564
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 9996 12880 10060 12884
rect 9996 12824 10046 12880
rect 10046 12824 10060 12880
rect 9996 12820 10060 12824
rect 5580 12684 5644 12748
rect 3924 12548 3988 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 5396 12276 5460 12340
rect 15148 12140 15212 12204
rect 4844 12004 4908 12068
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 1900 11596 1964 11660
rect 5028 11460 5092 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 3372 11188 3436 11252
rect 8156 11052 8220 11116
rect 13860 11112 13924 11116
rect 13860 11056 13910 11112
rect 13910 11056 13924 11112
rect 13860 11052 13924 11056
rect 15148 11052 15212 11116
rect 5580 10916 5644 10980
rect 3924 10840 3988 10844
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 3924 10784 3974 10840
rect 3974 10784 3988 10840
rect 3924 10780 3988 10784
rect 6684 10840 6748 10844
rect 6684 10784 6698 10840
rect 6698 10784 6748 10840
rect 6684 10780 6748 10784
rect 3924 10644 3988 10708
rect 4844 10644 4908 10708
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 5764 9420 5828 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 13492 8876 13556 8940
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 3924 8060 3988 8124
rect 13124 7788 13188 7852
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 12020 7516 12084 7580
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 10548 6836 10612 6900
rect 12572 6700 12636 6764
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 9996 3980 10060 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 5211 36684 5277 36685
rect 5211 36620 5212 36684
rect 5276 36620 5277 36684
rect 5211 36619 5277 36620
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 5214 31770 5274 36619
rect 7235 36548 7301 36549
rect 7235 36484 7236 36548
rect 7300 36484 7301 36548
rect 7235 36483 7301 36484
rect 5214 31710 5458 31770
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 1899 26348 1965 26349
rect 1899 26284 1900 26348
rect 1964 26284 1965 26348
rect 1899 26283 1965 26284
rect 1902 11661 1962 26283
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 3371 23492 3437 23493
rect 3371 23428 3372 23492
rect 3436 23428 3437 23492
rect 3371 23427 3437 23428
rect 3187 23220 3253 23221
rect 3187 23156 3188 23220
rect 3252 23156 3253 23220
rect 3187 23155 3253 23156
rect 3190 18733 3250 23155
rect 3187 18732 3253 18733
rect 3187 18668 3188 18732
rect 3252 18668 3253 18732
rect 3187 18667 3253 18668
rect 1899 11660 1965 11661
rect 1899 11596 1900 11660
rect 1964 11596 1965 11660
rect 1899 11595 1965 11596
rect 3374 11253 3434 23427
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 5398 22810 5458 31710
rect 6499 27028 6565 27029
rect 6499 26964 6500 27028
rect 6564 26964 6565 27028
rect 6499 26963 6565 26964
rect 6131 26348 6197 26349
rect 6131 26284 6132 26348
rect 6196 26284 6197 26348
rect 6131 26283 6197 26284
rect 5398 22750 5642 22810
rect 5398 21181 5458 22750
rect 5582 22677 5642 22750
rect 5579 22676 5645 22677
rect 5579 22612 5580 22676
rect 5644 22612 5645 22676
rect 5579 22611 5645 22612
rect 5395 21180 5461 21181
rect 5395 21116 5396 21180
rect 5460 21116 5461 21180
rect 5395 21115 5461 21116
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 3923 17508 3989 17509
rect 3923 17444 3924 17508
rect 3988 17444 3989 17508
rect 3923 17443 3989 17444
rect 3926 13565 3986 17443
rect 4208 16896 4528 17920
rect 5027 16964 5093 16965
rect 5027 16900 5028 16964
rect 5092 16900 5093 16964
rect 5027 16899 5093 16900
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 3923 13564 3989 13565
rect 3923 13500 3924 13564
rect 3988 13500 3989 13564
rect 3923 13499 3989 13500
rect 3923 12612 3989 12613
rect 3923 12548 3924 12612
rect 3988 12548 3989 12612
rect 3923 12547 3989 12548
rect 3371 11252 3437 11253
rect 3371 11188 3372 11252
rect 3436 11188 3437 11252
rect 3371 11187 3437 11188
rect 3926 10845 3986 12547
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4843 12068 4909 12069
rect 4843 12004 4844 12068
rect 4908 12004 4909 12068
rect 4843 12003 4909 12004
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 3923 10844 3989 10845
rect 3923 10780 3924 10844
rect 3988 10780 3989 10844
rect 3923 10779 3989 10780
rect 3923 10708 3989 10709
rect 3923 10644 3924 10708
rect 3988 10644 3989 10708
rect 3923 10643 3989 10644
rect 3926 8125 3986 10643
rect 4208 10368 4528 11392
rect 4846 10709 4906 12003
rect 5030 11525 5090 16899
rect 5395 16692 5461 16693
rect 5395 16628 5396 16692
rect 5460 16628 5461 16692
rect 5395 16627 5461 16628
rect 5398 12341 5458 16627
rect 6134 13701 6194 26283
rect 6502 17645 6562 26963
rect 7238 24853 7298 36483
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 9443 29068 9509 29069
rect 9443 29004 9444 29068
rect 9508 29004 9509 29068
rect 9443 29003 9509 29004
rect 8155 24988 8221 24989
rect 8155 24924 8156 24988
rect 8220 24924 8221 24988
rect 8155 24923 8221 24924
rect 7235 24852 7301 24853
rect 7235 24788 7236 24852
rect 7300 24788 7301 24852
rect 7235 24787 7301 24788
rect 7971 23628 8037 23629
rect 7971 23564 7972 23628
rect 8036 23564 8037 23628
rect 7971 23563 8037 23564
rect 6683 20772 6749 20773
rect 6683 20708 6684 20772
rect 6748 20708 6749 20772
rect 6683 20707 6749 20708
rect 6499 17644 6565 17645
rect 6499 17580 6500 17644
rect 6564 17580 6565 17644
rect 6499 17579 6565 17580
rect 6131 13700 6197 13701
rect 6131 13636 6132 13700
rect 6196 13636 6197 13700
rect 6131 13635 6197 13636
rect 5763 13564 5829 13565
rect 5763 13500 5764 13564
rect 5828 13500 5829 13564
rect 5763 13499 5829 13500
rect 5579 12748 5645 12749
rect 5579 12684 5580 12748
rect 5644 12684 5645 12748
rect 5579 12683 5645 12684
rect 5395 12340 5461 12341
rect 5395 12276 5396 12340
rect 5460 12276 5461 12340
rect 5395 12275 5461 12276
rect 5027 11524 5093 11525
rect 5027 11460 5028 11524
rect 5092 11460 5093 11524
rect 5027 11459 5093 11460
rect 5582 10981 5642 12683
rect 5579 10980 5645 10981
rect 5579 10916 5580 10980
rect 5644 10916 5645 10980
rect 5579 10915 5645 10916
rect 4843 10708 4909 10709
rect 4843 10644 4844 10708
rect 4908 10644 4909 10708
rect 4843 10643 4909 10644
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 5766 9485 5826 13499
rect 6686 10845 6746 20707
rect 7974 15197 8034 23563
rect 8158 18189 8218 24923
rect 9446 18733 9506 29003
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 15883 19684 15949 19685
rect 15883 19620 15884 19684
rect 15948 19620 15949 19684
rect 15883 19619 15949 19620
rect 12019 19412 12085 19413
rect 12019 19348 12020 19412
rect 12084 19348 12085 19412
rect 12019 19347 12085 19348
rect 9443 18732 9509 18733
rect 9443 18668 9444 18732
rect 9508 18668 9509 18732
rect 9443 18667 9509 18668
rect 8155 18188 8221 18189
rect 8155 18124 8156 18188
rect 8220 18124 8221 18188
rect 8155 18123 8221 18124
rect 8155 17644 8221 17645
rect 8155 17580 8156 17644
rect 8220 17580 8221 17644
rect 8155 17579 8221 17580
rect 7971 15196 8037 15197
rect 7971 15132 7972 15196
rect 8036 15132 8037 15196
rect 7971 15131 8037 15132
rect 8158 11117 8218 17579
rect 10547 13836 10613 13837
rect 10547 13772 10548 13836
rect 10612 13772 10613 13836
rect 10547 13771 10613 13772
rect 9995 12884 10061 12885
rect 9995 12820 9996 12884
rect 10060 12820 10061 12884
rect 9995 12819 10061 12820
rect 8155 11116 8221 11117
rect 8155 11052 8156 11116
rect 8220 11052 8221 11116
rect 8155 11051 8221 11052
rect 6683 10844 6749 10845
rect 6683 10780 6684 10844
rect 6748 10780 6749 10844
rect 6683 10779 6749 10780
rect 5763 9484 5829 9485
rect 5763 9420 5764 9484
rect 5828 9420 5829 9484
rect 5763 9419 5829 9420
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 3923 8124 3989 8125
rect 3923 8060 3924 8124
rect 3988 8060 3989 8124
rect 3923 8059 3989 8060
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 9998 4045 10058 12819
rect 10550 6901 10610 13771
rect 12022 7581 12082 19347
rect 13491 18052 13557 18053
rect 13491 17988 13492 18052
rect 13556 17988 13557 18052
rect 13491 17987 13557 17988
rect 13123 16692 13189 16693
rect 13123 16628 13124 16692
rect 13188 16628 13189 16692
rect 13123 16627 13189 16628
rect 12571 16420 12637 16421
rect 12571 16356 12572 16420
rect 12636 16356 12637 16420
rect 12571 16355 12637 16356
rect 12019 7580 12085 7581
rect 12019 7516 12020 7580
rect 12084 7516 12085 7580
rect 12019 7515 12085 7516
rect 10547 6900 10613 6901
rect 10547 6836 10548 6900
rect 10612 6836 10613 6900
rect 10547 6835 10613 6836
rect 12574 6765 12634 16355
rect 13126 7853 13186 16627
rect 13494 8941 13554 17987
rect 13859 17916 13925 17917
rect 13859 17852 13860 17916
rect 13924 17852 13925 17916
rect 13859 17851 13925 17852
rect 13862 11117 13922 17851
rect 15147 17644 15213 17645
rect 15147 17580 15148 17644
rect 15212 17580 15213 17644
rect 15147 17579 15213 17580
rect 15150 12205 15210 17579
rect 15886 14381 15946 19619
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 15883 14380 15949 14381
rect 15883 14316 15884 14380
rect 15948 14316 15949 14380
rect 15883 14315 15949 14316
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 15147 12204 15213 12205
rect 15147 12140 15148 12204
rect 15212 12140 15213 12204
rect 15147 12139 15213 12140
rect 15150 11117 15210 12139
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 13859 11116 13925 11117
rect 13859 11052 13860 11116
rect 13924 11052 13925 11116
rect 13859 11051 13925 11052
rect 15147 11116 15213 11117
rect 15147 11052 15148 11116
rect 15212 11052 15213 11116
rect 15147 11051 15213 11052
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 13491 8940 13557 8941
rect 13491 8876 13492 8940
rect 13556 8876 13557 8940
rect 13491 8875 13557 8876
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 13123 7852 13189 7853
rect 13123 7788 13124 7852
rect 13188 7788 13189 7852
rect 13123 7787 13189 7788
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 12571 6764 12637 6765
rect 12571 6700 12572 6764
rect 12636 6700 12637 6764
rect 12571 6699 12637 6700
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 9995 4044 10061 4045
rect 9995 3980 9996 4044
rect 10060 3980 10061 4044
rect 9995 3979 10061 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20
timestamp 1667941163
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62
timestamp 1667941163
transform 1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70
timestamp 1667941163
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76
timestamp 1667941163
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1667941163
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1667941163
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1667941163
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_154
timestamp 1667941163
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1667941163
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_174
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_186 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1667941163
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_210
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_238
timestamp 1667941163
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 1667941163
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_294
timestamp 1667941163
transform 1 0 28152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1667941163
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_322
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1667941163
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_342
timestamp 1667941163
transform 1 0 32568 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 1667941163
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1667941163
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 1667941163
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_399
timestamp 1667941163
transform 1 0 37812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1667941163
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1667941163
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_29
timestamp 1667941163
transform 1 0 3772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_41
timestamp 1667941163
transform 1 0 4876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1667941163
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_89
timestamp 1667941163
transform 1 0 9292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1667941163
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1667941163
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1667941163
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_34
timestamp 1667941163
transform 1 0 4232 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_46
timestamp 1667941163
transform 1 0 5336 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_58
timestamp 1667941163
transform 1 0 6440 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_70
timestamp 1667941163
transform 1 0 7544 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_9
timestamp 1667941163
transform 1 0 1932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_17
timestamp 1667941163
transform 1 0 2668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_21
timestamp 1667941163
transform 1 0 3036 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_28
timestamp 1667941163
transform 1 0 3680 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_40
timestamp 1667941163
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1667941163
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_89
timestamp 1667941163
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_95
timestamp 1667941163
transform 1 0 9844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1667941163
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_8
timestamp 1667941163
transform 1 0 1840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22
timestamp 1667941163
transform 1 0 3128 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1667941163
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp 1667941163
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_93
timestamp 1667941163
transform 1 0 9660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_105
timestamp 1667941163
transform 1 0 10764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_117
timestamp 1667941163
transform 1 0 11868 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_129
timestamp 1667941163
transform 1 0 12972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1667941163
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_171
timestamp 1667941163
transform 1 0 16836 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_175
timestamp 1667941163
transform 1 0 17204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1667941163
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_20
timestamp 1667941163
transform 1 0 2944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1667941163
transform 1 0 4508 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1667941163
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_75
timestamp 1667941163
transform 1 0 8004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_87
timestamp 1667941163
transform 1 0 9108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_99
timestamp 1667941163
transform 1 0 10212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_174
timestamp 1667941163
transform 1 0 17112 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_186
timestamp 1667941163
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_198
timestamp 1667941163
transform 1 0 19320 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_206
timestamp 1667941163
transform 1 0 20056 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_210
timestamp 1667941163
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1667941163
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_268
timestamp 1667941163
transform 1 0 25760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_286
timestamp 1667941163
transform 1 0 27416 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_298
timestamp 1667941163
transform 1 0 28520 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_310
timestamp 1667941163
transform 1 0 29624 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_322
timestamp 1667941163
transform 1 0 30728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1667941163
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_398
timestamp 1667941163
transform 1 0 37720 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1667941163
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_8
timestamp 1667941163
transform 1 0 1840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_19
timestamp 1667941163
transform 1 0 2852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_38
timestamp 1667941163
transform 1 0 4600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1667941163
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1667941163
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_64
timestamp 1667941163
transform 1 0 6992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_68
timestamp 1667941163
transform 1 0 7360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_75
timestamp 1667941163
transform 1 0 8004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1667941163
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1667941163
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_98
timestamp 1667941163
transform 1 0 10120 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_110
timestamp 1667941163
transform 1 0 11224 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_122
timestamp 1667941163
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1667941163
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_159
timestamp 1667941163
transform 1 0 15732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_171
timestamp 1667941163
transform 1 0 16836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_183
timestamp 1667941163
transform 1 0 17940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_348
timestamp 1667941163
transform 1 0 33120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1667941163
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_385
timestamp 1667941163
transform 1 0 36524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_391
timestamp 1667941163
transform 1 0 37076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_399
timestamp 1667941163
transform 1 0 37812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_8
timestamp 1667941163
transform 1 0 1840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1667941163
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_26
timestamp 1667941163
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_30
timestamp 1667941163
transform 1 0 3864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1667941163
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1667941163
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1667941163
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_62
timestamp 1667941163
transform 1 0 6808 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_74
timestamp 1667941163
transform 1 0 7912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1667941163
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_85
timestamp 1667941163
transform 1 0 8924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_97
timestamp 1667941163
transform 1 0 10028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1667941163
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_289
timestamp 1667941163
transform 1 0 27692 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_295
timestamp 1667941163
transform 1 0 28244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_307
timestamp 1667941163
transform 1 0 29348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_319
timestamp 1667941163
transform 1 0 30452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_331
timestamp 1667941163
transform 1 0 31556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1667941163
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_19
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1667941163
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_47
timestamp 1667941163
transform 1 0 5428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_54
timestamp 1667941163
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_61
timestamp 1667941163
transform 1 0 6716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_73
timestamp 1667941163
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1667941163
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_96
timestamp 1667941163
transform 1 0 9936 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_108
timestamp 1667941163
transform 1 0 11040 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_120
timestamp 1667941163
transform 1 0 12144 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1667941163
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_146
timestamp 1667941163
transform 1 0 14536 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_158
timestamp 1667941163
transform 1 0 15640 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_170
timestamp 1667941163
transform 1 0 16744 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_182
timestamp 1667941163
transform 1 0 17848 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1667941163
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_217
timestamp 1667941163
transform 1 0 21068 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_314
timestamp 1667941163
transform 1 0 29992 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_323
timestamp 1667941163
transform 1 0 30820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_335
timestamp 1667941163
transform 1 0 31924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_347
timestamp 1667941163
transform 1 0 33028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1667941163
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_372
timestamp 1667941163
transform 1 0 35328 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_384
timestamp 1667941163
transform 1 0 36432 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_396
timestamp 1667941163
transform 1 0 37536 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_404
timestamp 1667941163
transform 1 0 38272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1667941163
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1667941163
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1667941163
transform 1 0 3864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_62
timestamp 1667941163
transform 1 0 6808 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_74
timestamp 1667941163
transform 1 0 7912 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_86
timestamp 1667941163
transform 1 0 9016 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_90
timestamp 1667941163
transform 1 0 9384 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_102
timestamp 1667941163
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_253
timestamp 1667941163
transform 1 0 24380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_257
timestamp 1667941163
transform 1 0 24748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1667941163
transform 1 0 25852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1667941163
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_357
timestamp 1667941163
transform 1 0 33948 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_363
timestamp 1667941163
transform 1 0 34500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_375
timestamp 1667941163
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 1667941163
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_401
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_38
timestamp 1667941163
transform 1 0 4600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_42
timestamp 1667941163
transform 1 0 4968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_63
timestamp 1667941163
transform 1 0 6900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_70
timestamp 1667941163
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_78
timestamp 1667941163
transform 1 0 8280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_96
timestamp 1667941163
transform 1 0 9936 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_108
timestamp 1667941163
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_115
timestamp 1667941163
transform 1 0 11684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_127
timestamp 1667941163
transform 1 0 12788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_371
timestamp 1667941163
transform 1 0 35236 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_375
timestamp 1667941163
transform 1 0 35604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_387
timestamp 1667941163
transform 1 0 36708 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_399
timestamp 1667941163
transform 1 0 37812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_26
timestamp 1667941163
transform 1 0 3496 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1667941163
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_76
timestamp 1667941163
transform 1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_80
timestamp 1667941163
transform 1 0 8464 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_84
timestamp 1667941163
transform 1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_91
timestamp 1667941163
transform 1 0 9476 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_99
timestamp 1667941163
transform 1 0 10212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_103
timestamp 1667941163
transform 1 0 10580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_118
timestamp 1667941163
transform 1 0 11960 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_124
timestamp 1667941163
transform 1 0 12512 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_128
timestamp 1667941163
transform 1 0 12880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_140
timestamp 1667941163
transform 1 0 13984 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_146
timestamp 1667941163
transform 1 0 14536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_150
timestamp 1667941163
transform 1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_157
timestamp 1667941163
transform 1 0 15548 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1667941163
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_174
timestamp 1667941163
transform 1 0 17112 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_186
timestamp 1667941163
transform 1 0 18216 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_198
timestamp 1667941163
transform 1 0 19320 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_210
timestamp 1667941163
transform 1 0 20424 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1667941163
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_34
timestamp 1667941163
transform 1 0 4232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_45
timestamp 1667941163
transform 1 0 5244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_49
timestamp 1667941163
transform 1 0 5612 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_70
timestamp 1667941163
transform 1 0 7544 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_78
timestamp 1667941163
transform 1 0 8280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_96
timestamp 1667941163
transform 1 0 9936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_103
timestamp 1667941163
transform 1 0 10580 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_113
timestamp 1667941163
transform 1 0 11500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1667941163
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_124
timestamp 1667941163
transform 1 0 12512 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_128
timestamp 1667941163
transform 1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1667941163
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1667941163
transform 1 0 14628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1667941163
transform 1 0 15272 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_161
timestamp 1667941163
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_168
timestamp 1667941163
transform 1 0 16560 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_180
timestamp 1667941163
transform 1 0 17664 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1667941163
transform 1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1667941163
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_264
timestamp 1667941163
transform 1 0 25392 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_276
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_288
timestamp 1667941163
transform 1 0 27600 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_300
timestamp 1667941163
transform 1 0 28704 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_326
timestamp 1667941163
transform 1 0 31096 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_338
timestamp 1667941163
transform 1 0 32200 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_350
timestamp 1667941163
transform 1 0 33304 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1667941163
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_9
timestamp 1667941163
transform 1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_36
timestamp 1667941163
transform 1 0 4416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_43
timestamp 1667941163
transform 1 0 5060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1667941163
transform 1 0 6808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_124
timestamp 1667941163
transform 1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1667941163
transform 1 0 13156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_138
timestamp 1667941163
transform 1 0 13800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1667941163
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_152
timestamp 1667941163
transform 1 0 15088 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_159
timestamp 1667941163
transform 1 0 15732 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_174
timestamp 1667941163
transform 1 0 17112 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_183
timestamp 1667941163
transform 1 0 17940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_195
timestamp 1667941163
transform 1 0 19044 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_207
timestamp 1667941163
transform 1 0 20148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1667941163
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_366
timestamp 1667941163
transform 1 0 34776 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_378
timestamp 1667941163
transform 1 0 35880 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1667941163
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_34
timestamp 1667941163
transform 1 0 4232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1667941163
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_91
timestamp 1667941163
transform 1 0 9476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_98
timestamp 1667941163
transform 1 0 10120 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_105
timestamp 1667941163
transform 1 0 10764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_112
timestamp 1667941163
transform 1 0 11408 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_119
timestamp 1667941163
transform 1 0 12052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_126
timestamp 1667941163
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_147
timestamp 1667941163
transform 1 0 14628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_151
timestamp 1667941163
transform 1 0 14996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_160
timestamp 1667941163
transform 1 0 15824 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_167
timestamp 1667941163
transform 1 0 16468 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_178
timestamp 1667941163
transform 1 0 17480 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_185
timestamp 1667941163
transform 1 0 18124 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1667941163
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_370
timestamp 1667941163
transform 1 0 35144 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_382
timestamp 1667941163
transform 1 0 36248 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_394
timestamp 1667941163
transform 1 0 37352 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1667941163
transform 1 0 38456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_26
timestamp 1667941163
transform 1 0 3496 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1667941163
transform 1 0 6808 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_70
timestamp 1667941163
transform 1 0 7544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_91
timestamp 1667941163
transform 1 0 9476 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_95
timestamp 1667941163
transform 1 0 9844 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1667941163
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1667941163
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1667941163
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_121
timestamp 1667941163
transform 1 0 12236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_128
timestamp 1667941163
transform 1 0 12880 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_144
timestamp 1667941163
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_151
timestamp 1667941163
transform 1 0 14996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_155
timestamp 1667941163
transform 1 0 15364 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1667941163
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1667941163
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_185
timestamp 1667941163
transform 1 0 18124 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_194
timestamp 1667941163
transform 1 0 18952 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 1667941163
transform 1 0 19780 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_210
timestamp 1667941163
transform 1 0 20424 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_313
timestamp 1667941163
transform 1 0 29900 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1667941163
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1667941163
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_54
timestamp 1667941163
transform 1 0 6072 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1667941163
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_108
timestamp 1667941163
transform 1 0 11040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_114
timestamp 1667941163
transform 1 0 11592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1667941163
transform 1 0 11960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1667941163
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1667941163
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_147
timestamp 1667941163
transform 1 0 14628 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_158
timestamp 1667941163
transform 1 0 15640 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1667941163
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1667941163
transform 1 0 16836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1667941163
transform 1 0 17480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1667941163
transform 1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1667941163
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_204
timestamp 1667941163
transform 1 0 19872 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_211
timestamp 1667941163
transform 1 0 20516 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_223
timestamp 1667941163
transform 1 0 21620 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_235
timestamp 1667941163
transform 1 0 22724 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1667941163
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1667941163
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_33
timestamp 1667941163
transform 1 0 4140 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_43
timestamp 1667941163
transform 1 0 5060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_64
timestamp 1667941163
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_88
timestamp 1667941163
transform 1 0 9200 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_100
timestamp 1667941163
transform 1 0 10304 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1667941163
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1667941163
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_130
timestamp 1667941163
transform 1 0 13064 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1667941163
transform 1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_146
timestamp 1667941163
transform 1 0 14536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_150
timestamp 1667941163
transform 1 0 14904 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1667941163
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 1667941163
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1667941163
transform 1 0 17572 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_186
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_204
timestamp 1667941163
transform 1 0 19872 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_211
timestamp 1667941163
transform 1 0 20516 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_215
timestamp 1667941163
transform 1 0 20884 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1667941163
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_231
timestamp 1667941163
transform 1 0 22356 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_238
timestamp 1667941163
transform 1 0 23000 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_245
timestamp 1667941163
transform 1 0 23644 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_257
timestamp 1667941163
transform 1 0 24748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1667941163
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1667941163
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_285
timestamp 1667941163
transform 1 0 27324 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_289
timestamp 1667941163
transform 1 0 27692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_301
timestamp 1667941163
transform 1 0 28796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_313
timestamp 1667941163
transform 1 0 29900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_325
timestamp 1667941163
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1667941163
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_357
timestamp 1667941163
transform 1 0 33948 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_362
timestamp 1667941163
transform 1 0 34408 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_374
timestamp 1667941163
transform 1 0 35512 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_386
timestamp 1667941163
transform 1 0 36616 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_401
timestamp 1667941163
transform 1 0 37996 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1667941163
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1667941163
transform 1 0 6072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_58
timestamp 1667941163
transform 1 0 6440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1667941163
transform 1 0 10948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1667941163
transform 1 0 12052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_131
timestamp 1667941163
transform 1 0 13156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_146
timestamp 1667941163
transform 1 0 14536 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1667941163
transform 1 0 15640 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1667941163
transform 1 0 16744 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_182
timestamp 1667941163
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_203
timestamp 1667941163
transform 1 0 19780 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_217
timestamp 1667941163
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1667941163
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_228
timestamp 1667941163
transform 1 0 22080 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_232
timestamp 1667941163
transform 1 0 22448 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1667941163
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1667941163
transform 1 0 6808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_120
timestamp 1667941163
transform 1 0 12144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_132
timestamp 1667941163
transform 1 0 13248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_140
timestamp 1667941163
transform 1 0 13984 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1667941163
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1667941163
transform 1 0 14996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1667941163
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1667941163
transform 1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_207
timestamp 1667941163
transform 1 0 20148 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1667941163
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1667941163
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_251
timestamp 1667941163
transform 1 0 24196 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_263
timestamp 1667941163
transform 1 0 25300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1667941163
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_309
timestamp 1667941163
transform 1 0 29532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_313
timestamp 1667941163
transform 1 0 29900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_325
timestamp 1667941163
transform 1 0 31004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1667941163
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_35
timestamp 1667941163
transform 1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_39
timestamp 1667941163
transform 1 0 4692 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_43
timestamp 1667941163
transform 1 0 5060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_68
timestamp 1667941163
transform 1 0 7360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_75
timestamp 1667941163
transform 1 0 8004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1667941163
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_119
timestamp 1667941163
transform 1 0 12052 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_127
timestamp 1667941163
transform 1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_154
timestamp 1667941163
transform 1 0 15272 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_162
timestamp 1667941163
transform 1 0 16008 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_171
timestamp 1667941163
transform 1 0 16836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_179
timestamp 1667941163
transform 1 0 17572 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1667941163
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1667941163
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_212
timestamp 1667941163
transform 1 0 20608 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1667941163
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_226
timestamp 1667941163
transform 1 0 21896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_239
timestamp 1667941163
transform 1 0 23092 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1667941163
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_317
timestamp 1667941163
transform 1 0 30268 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_323
timestamp 1667941163
transform 1 0 30820 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_335
timestamp 1667941163
transform 1 0 31924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_347
timestamp 1667941163
transform 1 0 33028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_359
timestamp 1667941163
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_28
timestamp 1667941163
transform 1 0 3680 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1667941163
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1667941163
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1667941163
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1667941163
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_124
timestamp 1667941163
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_128
timestamp 1667941163
transform 1 0 12880 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1667941163
transform 1 0 13248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1667941163
transform 1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1667941163
transform 1 0 15548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1667941163
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_174
timestamp 1667941163
transform 1 0 17112 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1667941163
transform 1 0 18032 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_191
timestamp 1667941163
transform 1 0 18676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_197
timestamp 1667941163
transform 1 0 19228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_206
timestamp 1667941163
transform 1 0 20056 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_244
timestamp 1667941163
transform 1 0 23552 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_251
timestamp 1667941163
transform 1 0 24196 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_263
timestamp 1667941163
transform 1 0 25300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1667941163
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_370
timestamp 1667941163
transform 1 0 35144 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_382
timestamp 1667941163
transform 1 0 36248 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1667941163
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1667941163
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_72
timestamp 1667941163
transform 1 0 7728 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_78
timestamp 1667941163
transform 1 0 8280 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_107
timestamp 1667941163
transform 1 0 10948 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_124
timestamp 1667941163
transform 1 0 12512 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_152
timestamp 1667941163
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_159
timestamp 1667941163
transform 1 0 15732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_171
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1667941163
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_202
timestamp 1667941163
transform 1 0 19688 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_214
timestamp 1667941163
transform 1 0 20792 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_218
timestamp 1667941163
transform 1 0 21160 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_222
timestamp 1667941163
transform 1 0 21528 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_226
timestamp 1667941163
transform 1 0 21896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_235
timestamp 1667941163
transform 1 0 22724 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_242
timestamp 1667941163
transform 1 0 23368 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1667941163
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_258
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_351
timestamp 1667941163
transform 1 0 33396 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_355
timestamp 1667941163
transform 1 0 33764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_9
timestamp 1667941163
transform 1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_16
timestamp 1667941163
transform 1 0 2576 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_23
timestamp 1667941163
transform 1 0 3220 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1667941163
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_80
timestamp 1667941163
transform 1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1667941163
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_124
timestamp 1667941163
transform 1 0 12512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_136
timestamp 1667941163
transform 1 0 13616 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_144
timestamp 1667941163
transform 1 0 14352 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1667941163
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1667941163
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_177
timestamp 1667941163
transform 1 0 17388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1667941163
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_194
timestamp 1667941163
transform 1 0 18952 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_203
timestamp 1667941163
transform 1 0 19780 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1667941163
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_234
timestamp 1667941163
transform 1 0 22632 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1667941163
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_251
timestamp 1667941163
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_258
timestamp 1667941163
transform 1 0 24840 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_270
timestamp 1667941163
transform 1 0 25944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_308
timestamp 1667941163
transform 1 0 29440 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_320
timestamp 1667941163
transform 1 0 30544 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1667941163
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1667941163
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1667941163
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_68
timestamp 1667941163
transform 1 0 7360 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_107
timestamp 1667941163
transform 1 0 10948 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1667941163
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_128
timestamp 1667941163
transform 1 0 12880 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1667941163
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_147
timestamp 1667941163
transform 1 0 14628 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_160
timestamp 1667941163
transform 1 0 15824 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_168
timestamp 1667941163
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_173
timestamp 1667941163
transform 1 0 17020 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_186
timestamp 1667941163
transform 1 0 18216 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_190
timestamp 1667941163
transform 1 0 18584 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_211
timestamp 1667941163
transform 1 0 20516 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_226
timestamp 1667941163
transform 1 0 21896 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_243
timestamp 1667941163
transform 1 0 23460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_258
timestamp 1667941163
transform 1 0 24840 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_270
timestamp 1667941163
transform 1 0 25944 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_282
timestamp 1667941163
transform 1 0 27048 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_294
timestamp 1667941163
transform 1 0 28152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1667941163
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_17
timestamp 1667941163
transform 1 0 2668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_42
timestamp 1667941163
transform 1 0 4968 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_50
timestamp 1667941163
transform 1 0 5704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_64
timestamp 1667941163
transform 1 0 6992 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_68
timestamp 1667941163
transform 1 0 7360 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_90
timestamp 1667941163
transform 1 0 9384 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_96
timestamp 1667941163
transform 1 0 9936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1667941163
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_147
timestamp 1667941163
transform 1 0 14628 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_173
timestamp 1667941163
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_177
timestamp 1667941163
transform 1 0 17388 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_189
timestamp 1667941163
transform 1 0 18492 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_197
timestamp 1667941163
transform 1 0 19228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_206
timestamp 1667941163
transform 1 0 20056 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1667941163
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_235
timestamp 1667941163
transform 1 0 22724 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_242
timestamp 1667941163
transform 1 0 23368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_256
timestamp 1667941163
transform 1 0 24656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_263
timestamp 1667941163
transform 1 0 25300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1667941163
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1667941163
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1667941163
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_56
timestamp 1667941163
transform 1 0 6256 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1667941163
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_107
timestamp 1667941163
transform 1 0 10948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_131
timestamp 1667941163
transform 1 0 13156 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1667941163
transform 1 0 14720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_161
timestamp 1667941163
transform 1 0 15916 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_168
timestamp 1667941163
transform 1 0 16560 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1667941163
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_213
timestamp 1667941163
transform 1 0 20700 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1667941163
transform 1 0 21252 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_223
timestamp 1667941163
transform 1 0 21620 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_229
timestamp 1667941163
transform 1 0 22172 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_238
timestamp 1667941163
transform 1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_263
timestamp 1667941163
transform 1 0 25300 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_270
timestamp 1667941163
transform 1 0 25944 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_282
timestamp 1667941163
transform 1 0 27048 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_294
timestamp 1667941163
transform 1 0 28152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1667941163
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_370
timestamp 1667941163
transform 1 0 35144 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_382
timestamp 1667941163
transform 1 0 36248 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_394
timestamp 1667941163
transform 1 0 37352 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1667941163
transform 1 0 38456 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_34
timestamp 1667941163
transform 1 0 4232 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_42
timestamp 1667941163
transform 1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_47
timestamp 1667941163
transform 1 0 5428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_64
timestamp 1667941163
transform 1 0 6992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_88
timestamp 1667941163
transform 1 0 9200 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_94
timestamp 1667941163
transform 1 0 9752 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_104
timestamp 1667941163
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_135
timestamp 1667941163
transform 1 0 13524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_147
timestamp 1667941163
transform 1 0 14628 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_155
timestamp 1667941163
transform 1 0 15364 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1667941163
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1667941163
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_190
timestamp 1667941163
transform 1 0 18584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_202
timestamp 1667941163
transform 1 0 19688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1667941163
transform 1 0 20332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1667941163
transform 1 0 20700 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_230
timestamp 1667941163
transform 1 0 22264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_245
timestamp 1667941163
transform 1 0 23644 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_255
timestamp 1667941163
transform 1 0 24564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_268
timestamp 1667941163
transform 1 0 25760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1667941163
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_298
timestamp 1667941163
transform 1 0 28520 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_310
timestamp 1667941163
transform 1 0 29624 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_322
timestamp 1667941163
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1667941163
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_358
timestamp 1667941163
transform 1 0 34040 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_370
timestamp 1667941163
transform 1 0 35144 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_382
timestamp 1667941163
transform 1 0 36248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1667941163
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 1667941163
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_34
timestamp 1667941163
transform 1 0 4232 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1667941163
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1667941163
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1667941163
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_107
timestamp 1667941163
transform 1 0 10948 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_120
timestamp 1667941163
transform 1 0 12144 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_128
timestamp 1667941163
transform 1 0 12880 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_151
timestamp 1667941163
transform 1 0 14996 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_164
timestamp 1667941163
transform 1 0 16192 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_168
timestamp 1667941163
transform 1 0 16560 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_172
timestamp 1667941163
transform 1 0 16928 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1667941163
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_191
timestamp 1667941163
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_206
timestamp 1667941163
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_219
timestamp 1667941163
transform 1 0 21252 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_235
timestamp 1667941163
transform 1 0 22724 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_247
timestamp 1667941163
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1667941163
transform 1 0 24840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_272
timestamp 1667941163
transform 1 0 26128 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_284
timestamp 1667941163
transform 1 0 27232 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_296
timestamp 1667941163
transform 1 0 28336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_314
timestamp 1667941163
transform 1 0 29992 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_326
timestamp 1667941163
transform 1 0 31096 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_338
timestamp 1667941163
transform 1 0 32200 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_350
timestamp 1667941163
transform 1 0 33304 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1667941163
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_26
timestamp 1667941163
transform 1 0 3496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_30
timestamp 1667941163
transform 1 0 3864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_80
timestamp 1667941163
transform 1 0 8464 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_104
timestamp 1667941163
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1667941163
transform 1 0 12420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_136
timestamp 1667941163
transform 1 0 13616 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1667941163
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1667941163
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_179
timestamp 1667941163
transform 1 0 17572 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_194
timestamp 1667941163
transform 1 0 18952 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_208
timestamp 1667941163
transform 1 0 20240 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_235
timestamp 1667941163
transform 1 0 22724 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_243
timestamp 1667941163
transform 1 0 23460 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_253
timestamp 1667941163
transform 1 0 24380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_260
timestamp 1667941163
transform 1 0 25024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_267
timestamp 1667941163
transform 1 0 25668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1667941163
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_357
timestamp 1667941163
transform 1 0 33948 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_362
timestamp 1667941163
transform 1 0 34408 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_374
timestamp 1667941163
transform 1 0 35512 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 1667941163
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1667941163
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_36
timestamp 1667941163
transform 1 0 4416 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1667941163
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_68
timestamp 1667941163
transform 1 0 7360 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_107
timestamp 1667941163
transform 1 0 10948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_113
timestamp 1667941163
transform 1 0 11500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_122
timestamp 1667941163
transform 1 0 12328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1667941163
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_150
timestamp 1667941163
transform 1 0 14904 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_163
timestamp 1667941163
transform 1 0 16100 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_176
timestamp 1667941163
transform 1 0 17296 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1667941163
transform 1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_207
timestamp 1667941163
transform 1 0 20148 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_216
timestamp 1667941163
transform 1 0 20976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_223
timestamp 1667941163
transform 1 0 21620 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_230
timestamp 1667941163
transform 1 0 22264 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_237
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1667941163
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1667941163
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1667941163
transform 1 0 26036 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_278
timestamp 1667941163
transform 1 0 26680 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_290
timestamp 1667941163
transform 1 0 27784 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1667941163
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_327
timestamp 1667941163
transform 1 0 31188 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_339
timestamp 1667941163
transform 1 0 32292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_351
timestamp 1667941163
transform 1 0 33396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_405
timestamp 1667941163
transform 1 0 38364 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_16
timestamp 1667941163
transform 1 0 2576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_23
timestamp 1667941163
transform 1 0 3220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1667941163
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_66
timestamp 1667941163
transform 1 0 7176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_91
timestamp 1667941163
transform 1 0 9476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1667941163
transform 1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1667941163
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1667941163
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_175
timestamp 1667941163
transform 1 0 17204 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1667941163
transform 1 0 18032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_196
timestamp 1667941163
transform 1 0 19136 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_210
timestamp 1667941163
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_230
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_238
timestamp 1667941163
transform 1 0 23000 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_247
timestamp 1667941163
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_259
timestamp 1667941163
transform 1 0 24932 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_266
timestamp 1667941163
transform 1 0 25576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_33
timestamp 1667941163
transform 1 0 4140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_37
timestamp 1667941163
transform 1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_44
timestamp 1667941163
transform 1 0 5152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_71
timestamp 1667941163
transform 1 0 7636 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_107
timestamp 1667941163
transform 1 0 10948 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_115
timestamp 1667941163
transform 1 0 11684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_125
timestamp 1667941163
transform 1 0 12604 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1667941163
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1667941163
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1667941163
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1667941163
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1667941163
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_203
timestamp 1667941163
transform 1 0 19780 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_210
timestamp 1667941163
transform 1 0 20424 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_217
timestamp 1667941163
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1667941163
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_231
timestamp 1667941163
transform 1 0 22356 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_239
timestamp 1667941163
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1667941163
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_258
timestamp 1667941163
transform 1 0 24840 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1667941163
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_9
timestamp 1667941163
transform 1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_13
timestamp 1667941163
transform 1 0 2300 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_37
timestamp 1667941163
transform 1 0 4508 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_43
timestamp 1667941163
transform 1 0 5060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_47
timestamp 1667941163
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1667941163
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_65
timestamp 1667941163
transform 1 0 7084 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_92
timestamp 1667941163
transform 1 0 9568 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_96
timestamp 1667941163
transform 1 0 9936 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_100
timestamp 1667941163
transform 1 0 10304 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_123
timestamp 1667941163
transform 1 0 12420 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_131
timestamp 1667941163
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_136
timestamp 1667941163
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_143
timestamp 1667941163
transform 1 0 14260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_150
timestamp 1667941163
transform 1 0 14904 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_162
timestamp 1667941163
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1667941163
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_177
timestamp 1667941163
transform 1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_189
timestamp 1667941163
transform 1 0 18492 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_196
timestamp 1667941163
transform 1 0 19136 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_203
timestamp 1667941163
transform 1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_210
timestamp 1667941163
transform 1 0 20424 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_218
timestamp 1667941163
transform 1 0 21160 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1667941163
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_239
timestamp 1667941163
transform 1 0 23092 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_246
timestamp 1667941163
transform 1 0 23736 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_253
timestamp 1667941163
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_265
timestamp 1667941163
transform 1 0 25484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1667941163
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1667941163
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_35
timestamp 1667941163
transform 1 0 4324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_39
timestamp 1667941163
transform 1 0 4692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_64
timestamp 1667941163
transform 1 0 6992 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_75
timestamp 1667941163
transform 1 0 8004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_107
timestamp 1667941163
transform 1 0 10948 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_115
timestamp 1667941163
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_125
timestamp 1667941163
transform 1 0 12604 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_151
timestamp 1667941163
transform 1 0 14996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_163
timestamp 1667941163
transform 1 0 16100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_169
timestamp 1667941163
transform 1 0 16652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_179
timestamp 1667941163
transform 1 0 17572 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_185
timestamp 1667941163
transform 1 0 18124 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1667941163
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_215
timestamp 1667941163
transform 1 0 20884 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_228
timestamp 1667941163
transform 1 0 22080 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_234
timestamp 1667941163
transform 1 0 22632 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1667941163
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_339
timestamp 1667941163
transform 1 0 32292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_351
timestamp 1667941163
transform 1 0 33396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_28
timestamp 1667941163
transform 1 0 3680 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_68
timestamp 1667941163
transform 1 0 7360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_92
timestamp 1667941163
transform 1 0 9568 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_96
timestamp 1667941163
transform 1 0 9936 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_100
timestamp 1667941163
transform 1 0 10304 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 1667941163
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_122
timestamp 1667941163
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_129
timestamp 1667941163
transform 1 0 12972 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_136
timestamp 1667941163
transform 1 0 13616 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_157
timestamp 1667941163
transform 1 0 15548 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_179
timestamp 1667941163
transform 1 0 17572 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_188
timestamp 1667941163
transform 1 0 18400 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_201
timestamp 1667941163
transform 1 0 19596 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_208
timestamp 1667941163
transform 1 0 20240 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_216
timestamp 1667941163
transform 1 0 20976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1667941163
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_230
timestamp 1667941163
transform 1 0 22264 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_239
timestamp 1667941163
transform 1 0 23092 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_251
timestamp 1667941163
transform 1 0 24196 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_263
timestamp 1667941163
transform 1 0 25300 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1667941163
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_310
timestamp 1667941163
transform 1 0 29624 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_318
timestamp 1667941163
transform 1 0 30360 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_323
timestamp 1667941163
transform 1 0 30820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_34
timestamp 1667941163
transform 1 0 4232 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_58
timestamp 1667941163
transform 1 0 6440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_107
timestamp 1667941163
transform 1 0 10948 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1667941163
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1667941163
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_152
timestamp 1667941163
transform 1 0 15088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1667941163
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_171
timestamp 1667941163
transform 1 0 16836 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_181
timestamp 1667941163
transform 1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_202
timestamp 1667941163
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_217
timestamp 1667941163
transform 1 0 21068 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_228
timestamp 1667941163
transform 1 0 22080 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_240
timestamp 1667941163
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_32
timestamp 1667941163
transform 1 0 4048 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_43
timestamp 1667941163
transform 1 0 5060 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_47
timestamp 1667941163
transform 1 0 5428 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1667941163
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_68
timestamp 1667941163
transform 1 0 7360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_92
timestamp 1667941163
transform 1 0 9568 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_100
timestamp 1667941163
transform 1 0 10304 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_123
timestamp 1667941163
transform 1 0 12420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1667941163
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_145
timestamp 1667941163
transform 1 0 14444 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_153
timestamp 1667941163
transform 1 0 15180 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1667941163
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_180
timestamp 1667941163
transform 1 0 17664 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_192
timestamp 1667941163
transform 1 0 18768 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_199
timestamp 1667941163
transform 1 0 19412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_215
timestamp 1667941163
transform 1 0 20884 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1667941163
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_34
timestamp 1667941163
transform 1 0 4232 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_52
timestamp 1667941163
transform 1 0 5888 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1667941163
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_96
timestamp 1667941163
transform 1 0 9936 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_112
timestamp 1667941163
transform 1 0 11408 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_116
timestamp 1667941163
transform 1 0 11776 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_125
timestamp 1667941163
transform 1 0 12604 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_155
timestamp 1667941163
transform 1 0 15364 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_161
timestamp 1667941163
transform 1 0 15916 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1667941163
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_175
timestamp 1667941163
transform 1 0 17204 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_179
timestamp 1667941163
transform 1 0 17572 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_185
timestamp 1667941163
transform 1 0 18124 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_207
timestamp 1667941163
transform 1 0 20148 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_214
timestamp 1667941163
transform 1 0 20792 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_226
timestamp 1667941163
transform 1 0 21896 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_238
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_8
timestamp 1667941163
transform 1 0 1840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_12
timestamp 1667941163
transform 1 0 2208 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_16
timestamp 1667941163
transform 1 0 2576 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_23
timestamp 1667941163
transform 1 0 3220 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_30
timestamp 1667941163
transform 1 0 3864 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_37
timestamp 1667941163
transform 1 0 4508 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_44
timestamp 1667941163
transform 1 0 5152 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_50
timestamp 1667941163
transform 1 0 5704 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1667941163
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_74
timestamp 1667941163
transform 1 0 7912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_86
timestamp 1667941163
transform 1 0 9016 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_92
timestamp 1667941163
transform 1 0 9568 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_101
timestamp 1667941163
transform 1 0 10396 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_126
timestamp 1667941163
transform 1 0 12696 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_135
timestamp 1667941163
transform 1 0 13524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1667941163
transform 1 0 14168 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1667941163
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_179
timestamp 1667941163
transform 1 0 17572 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1667941163
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_212
timestamp 1667941163
transform 1 0 20608 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_358
timestamp 1667941163
transform 1 0 34040 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_370
timestamp 1667941163
transform 1 0 35144 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_382
timestamp 1667941163
transform 1 0 36248 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1667941163
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_401
timestamp 1667941163
transform 1 0 37996 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_12
timestamp 1667941163
transform 1 0 2208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_19
timestamp 1667941163
transform 1 0 2852 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1667941163
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_39
timestamp 1667941163
transform 1 0 4692 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_45
timestamp 1667941163
transform 1 0 5244 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_54
timestamp 1667941163
transform 1 0 6072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_67
timestamp 1667941163
transform 1 0 7268 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1667941163
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_92
timestamp 1667941163
transform 1 0 9568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1667941163
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1667941163
transform 1 0 10856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_118
timestamp 1667941163
transform 1 0 11960 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_126
timestamp 1667941163
transform 1 0 12696 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_131
timestamp 1667941163
transform 1 0 13156 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1667941163
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_155
timestamp 1667941163
transform 1 0 15364 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_163
timestamp 1667941163
transform 1 0 16100 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_167
timestamp 1667941163
transform 1 0 16468 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1667941163
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_186
timestamp 1667941163
transform 1 0 18216 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_190
timestamp 1667941163
transform 1 0 18584 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_202
timestamp 1667941163
transform 1 0 19688 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_218
timestamp 1667941163
transform 1 0 21160 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_230
timestamp 1667941163
transform 1 0 22264 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_242
timestamp 1667941163
transform 1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1667941163
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_369
timestamp 1667941163
transform 1 0 35052 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_373
timestamp 1667941163
transform 1 0 35420 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_385
timestamp 1667941163
transform 1 0 36524 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_397
timestamp 1667941163
transform 1 0 37628 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_13
timestamp 1667941163
transform 1 0 2300 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_17
timestamp 1667941163
transform 1 0 2668 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_29
timestamp 1667941163
transform 1 0 3772 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_33
timestamp 1667941163
transform 1 0 4140 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_42
timestamp 1667941163
transform 1 0 4968 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_50
timestamp 1667941163
transform 1 0 5704 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1667941163
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_63
timestamp 1667941163
transform 1 0 6900 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_70
timestamp 1667941163
transform 1 0 7544 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_82
timestamp 1667941163
transform 1 0 8648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_89
timestamp 1667941163
transform 1 0 9292 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_96
timestamp 1667941163
transform 1 0 9936 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_103
timestamp 1667941163
transform 1 0 10580 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_123
timestamp 1667941163
transform 1 0 12420 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_136
timestamp 1667941163
transform 1 0 13616 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_150
timestamp 1667941163
transform 1 0 14904 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_156
timestamp 1667941163
transform 1 0 15456 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_165
timestamp 1667941163
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_185
timestamp 1667941163
transform 1 0 18124 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1667941163
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_214
timestamp 1667941163
transform 1 0 20792 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1667941163
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_7
timestamp 1667941163
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1667941163
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_18
timestamp 1667941163
transform 1 0 2760 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1667941163
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_40
timestamp 1667941163
transform 1 0 4784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_47
timestamp 1667941163
transform 1 0 5428 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_54
timestamp 1667941163
transform 1 0 6072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_61
timestamp 1667941163
transform 1 0 6716 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_68
timestamp 1667941163
transform 1 0 7360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_75
timestamp 1667941163
transform 1 0 8004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1667941163
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_91
timestamp 1667941163
transform 1 0 9476 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_98
timestamp 1667941163
transform 1 0 10120 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_105
timestamp 1667941163
transform 1 0 10764 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_113
timestamp 1667941163
transform 1 0 11500 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_118
timestamp 1667941163
transform 1 0 11960 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_125
timestamp 1667941163
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_146
timestamp 1667941163
transform 1 0 14536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_150
timestamp 1667941163
transform 1 0 14904 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_159
timestamp 1667941163
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_171
timestamp 1667941163
transform 1 0 16836 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_180
timestamp 1667941163
transform 1 0 17664 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1667941163
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_201
timestamp 1667941163
transform 1 0 19596 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_205
timestamp 1667941163
transform 1 0 19964 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_212
timestamp 1667941163
transform 1 0 20608 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_224
timestamp 1667941163
transform 1 0 21712 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_236
timestamp 1667941163
transform 1 0 22816 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1667941163
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_373
timestamp 1667941163
transform 1 0 35420 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_378
timestamp 1667941163
transform 1 0 35880 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_390
timestamp 1667941163
transform 1 0 36984 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_8
timestamp 1667941163
transform 1 0 1840 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_17
timestamp 1667941163
transform 1 0 2668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_24
timestamp 1667941163
transform 1 0 3312 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_31
timestamp 1667941163
transform 1 0 3956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_38
timestamp 1667941163
transform 1 0 4600 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_47
timestamp 1667941163
transform 1 0 5428 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1667941163
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_63
timestamp 1667941163
transform 1 0 6900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_67
timestamp 1667941163
transform 1 0 7268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_79
timestamp 1667941163
transform 1 0 8372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_88
timestamp 1667941163
transform 1 0 9200 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_100
timestamp 1667941163
transform 1 0 10304 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_106
timestamp 1667941163
transform 1 0 10856 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_118
timestamp 1667941163
transform 1 0 11960 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_132
timestamp 1667941163
transform 1 0 13248 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_138
timestamp 1667941163
transform 1 0 13800 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_142
timestamp 1667941163
transform 1 0 14168 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_155
timestamp 1667941163
transform 1 0 15364 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_159
timestamp 1667941163
transform 1 0 15732 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1667941163
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_179
timestamp 1667941163
transform 1 0 17572 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_183
timestamp 1667941163
transform 1 0 17940 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_192
timestamp 1667941163
transform 1 0 18768 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_198
timestamp 1667941163
transform 1 0 19320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_202
timestamp 1667941163
transform 1 0 19688 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_209
timestamp 1667941163
transform 1 0 20332 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1667941163
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_312
timestamp 1667941163
transform 1 0 29808 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_324
timestamp 1667941163
transform 1 0 30912 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_14
timestamp 1667941163
transform 1 0 2392 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1667941163
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_38
timestamp 1667941163
transform 1 0 4600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_45
timestamp 1667941163
transform 1 0 5244 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_51
timestamp 1667941163
transform 1 0 5796 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_60
timestamp 1667941163
transform 1 0 6624 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_68
timestamp 1667941163
transform 1 0 7360 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_78
timestamp 1667941163
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_90
timestamp 1667941163
transform 1 0 9384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_105
timestamp 1667941163
transform 1 0 10764 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_110
timestamp 1667941163
transform 1 0 11224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_117
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_124
timestamp 1667941163
transform 1 0 12512 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_131
timestamp 1667941163
transform 1 0 13156 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_147
timestamp 1667941163
transform 1 0 14628 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_155
timestamp 1667941163
transform 1 0 15364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_160
timestamp 1667941163
transform 1 0 15824 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_167
timestamp 1667941163
transform 1 0 16468 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_174
timestamp 1667941163
transform 1 0 17112 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_181
timestamp 1667941163
transform 1 0 17756 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1667941163
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_202
timestamp 1667941163
transform 1 0 19688 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_214
timestamp 1667941163
transform 1 0 20792 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_226
timestamp 1667941163
transform 1 0 21896 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_238
timestamp 1667941163
transform 1 0 23000 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1667941163
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_383
timestamp 1667941163
transform 1 0 36340 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_395
timestamp 1667941163
transform 1 0 37444 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_8
timestamp 1667941163
transform 1 0 1840 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_12
timestamp 1667941163
transform 1 0 2208 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_16
timestamp 1667941163
transform 1 0 2576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_23
timestamp 1667941163
transform 1 0 3220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_30
timestamp 1667941163
transform 1 0 3864 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_37
timestamp 1667941163
transform 1 0 4508 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_44
timestamp 1667941163
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_71
timestamp 1667941163
transform 1 0 7636 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_78
timestamp 1667941163
transform 1 0 8280 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_85
timestamp 1667941163
transform 1 0 8924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_97
timestamp 1667941163
transform 1 0 10028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1667941163
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_118
timestamp 1667941163
transform 1 0 11960 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_124
timestamp 1667941163
transform 1 0 12512 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_128
timestamp 1667941163
transform 1 0 12880 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_132
timestamp 1667941163
transform 1 0 13248 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_136
timestamp 1667941163
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_143
timestamp 1667941163
transform 1 0 14260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1667941163
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_159
timestamp 1667941163
transform 1 0 15732 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_179
timestamp 1667941163
transform 1 0 17572 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_185
timestamp 1667941163
transform 1 0 18124 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1667941163
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_196
timestamp 1667941163
transform 1 0 19136 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_208
timestamp 1667941163
transform 1 0 20240 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1667941163
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_314
timestamp 1667941163
transform 1 0 29992 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_326
timestamp 1667941163
transform 1 0 31096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1667941163
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_8
timestamp 1667941163
transform 1 0 1840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1667941163
transform 1 0 3128 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_34
timestamp 1667941163
transform 1 0 4232 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_49
timestamp 1667941163
transform 1 0 5612 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_55
timestamp 1667941163
transform 1 0 6164 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_62
timestamp 1667941163
transform 1 0 6808 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_69
timestamp 1667941163
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1667941163
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_90
timestamp 1667941163
transform 1 0 9384 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_102
timestamp 1667941163
transform 1 0 10488 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_114
timestamp 1667941163
transform 1 0 11592 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_126
timestamp 1667941163
transform 1 0 12696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_162
timestamp 1667941163
transform 1 0 16008 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1667941163
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_181
timestamp 1667941163
transform 1 0 17756 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1667941163
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_12
timestamp 1667941163
transform 1 0 2208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_19
timestamp 1667941163
transform 1 0 2852 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_25
timestamp 1667941163
transform 1 0 3404 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_29
timestamp 1667941163
transform 1 0 3772 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_36
timestamp 1667941163
transform 1 0 4416 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_48
timestamp 1667941163
transform 1 0 5520 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_64
timestamp 1667941163
transform 1 0 6992 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_76
timestamp 1667941163
transform 1 0 8096 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_88
timestamp 1667941163
transform 1 0 9200 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_100
timestamp 1667941163
transform 1 0 10304 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_157
timestamp 1667941163
transform 1 0 15548 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_163
timestamp 1667941163
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_174
timestamp 1667941163
transform 1 0 17112 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_186
timestamp 1667941163
transform 1 0 18216 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_198
timestamp 1667941163
transform 1 0 19320 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_210
timestamp 1667941163
transform 1 0 20424 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_356
timestamp 1667941163
transform 1 0 33856 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_368
timestamp 1667941163
transform 1 0 34960 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_380
timestamp 1667941163
transform 1 0 36064 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_17
timestamp 1667941163
transform 1 0 2668 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_25
timestamp 1667941163
transform 1 0 3404 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_34
timestamp 1667941163
transform 1 0 4232 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_46
timestamp 1667941163
transform 1 0 5336 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_58
timestamp 1667941163
transform 1 0 6440 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_70
timestamp 1667941163
transform 1 0 7544 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1667941163
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_168
timestamp 1667941163
transform 1 0 16560 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_180
timestamp 1667941163
transform 1 0 17664 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1667941163
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_204
timestamp 1667941163
transform 1 0 19872 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_216
timestamp 1667941163
transform 1 0 20976 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_228
timestamp 1667941163
transform 1 0 22080 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_240
timestamp 1667941163
transform 1 0 23184 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_349
timestamp 1667941163
transform 1 0 33212 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_353
timestamp 1667941163
transform 1 0 33580 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1667941163
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_12
timestamp 1667941163
transform 1 0 2208 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_19
timestamp 1667941163
transform 1 0 2852 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_31
timestamp 1667941163
transform 1 0 3956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_38
timestamp 1667941163
transform 1 0 4600 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1667941163
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_9
timestamp 1667941163
transform 1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1667941163
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_46
timestamp 1667941163
transform 1 0 5336 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_60
timestamp 1667941163
transform 1 0 6624 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_72
timestamp 1667941163
transform 1 0 7728 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_117
timestamp 1667941163
transform 1 0 11868 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_169
timestamp 1667941163
transform 1 0 16652 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_176
timestamp 1667941163
transform 1 0 17296 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_188
timestamp 1667941163
transform 1 0 18400 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_258
timestamp 1667941163
transform 1 0 24840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_262
timestamp 1667941163
transform 1 0 25208 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_266
timestamp 1667941163
transform 1 0 25576 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_278
timestamp 1667941163
transform 1 0 26680 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_290
timestamp 1667941163
transform 1 0 27784 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_302
timestamp 1667941163
transform 1 0 28888 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_317
timestamp 1667941163
transform 1 0 30268 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_11
timestamp 1667941163
transform 1 0 2116 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_18
timestamp 1667941163
transform 1 0 2760 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_30
timestamp 1667941163
transform 1 0 3864 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_42
timestamp 1667941163
transform 1 0 4968 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1667941163
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_62
timestamp 1667941163
transform 1 0 6808 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_74
timestamp 1667941163
transform 1 0 7912 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_86
timestamp 1667941163
transform 1 0 9016 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_98
timestamp 1667941163
transform 1 0 10120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_118
timestamp 1667941163
transform 1 0 11960 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_130
timestamp 1667941163
transform 1 0 13064 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_142
timestamp 1667941163
transform 1 0 14168 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_154
timestamp 1667941163
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_213
timestamp 1667941163
transform 1 0 20700 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_286
timestamp 1667941163
transform 1 0 27416 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_298
timestamp 1667941163
transform 1 0 28520 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_307
timestamp 1667941163
transform 1 0 29348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_319
timestamp 1667941163
transform 1 0 30452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_331
timestamp 1667941163
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_353
timestamp 1667941163
transform 1 0 33580 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_365
timestamp 1667941163
transform 1 0 34684 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_377
timestamp 1667941163
transform 1 0 35788 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 1667941163
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_401
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_8
timestamp 1667941163
transform 1 0 1840 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1667941163
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_34
timestamp 1667941163
transform 1 0 4232 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_46
timestamp 1667941163
transform 1 0 5336 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_57
timestamp 1667941163
transform 1 0 6348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_69
timestamp 1667941163
transform 1 0 7452 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_75
timestamp 1667941163
transform 1 0 8004 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_79
timestamp 1667941163
transform 1 0 8372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_370
timestamp 1667941163
transform 1 0 35144 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_382
timestamp 1667941163
transform 1 0 36248 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_394
timestamp 1667941163
transform 1 0 37352 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1667941163
transform 1 0 38456 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_174
timestamp 1667941163
transform 1 0 17112 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_186
timestamp 1667941163
transform 1 0 18216 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_198
timestamp 1667941163
transform 1 0 19320 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_210
timestamp 1667941163
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1667941163
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_242
timestamp 1667941163
transform 1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1667941163
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_48
timestamp 1667941163
transform 1 0 5520 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_358
timestamp 1667941163
transform 1 0 34040 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_370
timestamp 1667941163
transform 1 0 35144 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_382
timestamp 1667941163
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1667941163
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_8
timestamp 1667941163
transform 1 0 1840 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1667941163
transform 1 0 2944 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_141
timestamp 1667941163
transform 1 0 14076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_145
timestamp 1667941163
transform 1 0 14444 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_157
timestamp 1667941163
transform 1 0 15548 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1667941163
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_201
timestamp 1667941163
transform 1 0 19596 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_206
timestamp 1667941163
transform 1 0 20056 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_218
timestamp 1667941163
transform 1 0 21160 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_308
timestamp 1667941163
transform 1 0 29440 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_320
timestamp 1667941163
transform 1 0 30544 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1667941163
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1667941163
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_103
timestamp 1667941163
transform 1 0 10580 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_115
timestamp 1667941163
transform 1 0 11684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_127
timestamp 1667941163
transform 1 0 12788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_318
timestamp 1667941163
transform 1 0 30360 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_330
timestamp 1667941163
transform 1 0 31464 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_342
timestamp 1667941163
transform 1 0 32568 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_354
timestamp 1667941163
transform 1 0 33672 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1667941163
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1667941163
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1667941163
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1667941163
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1667941163
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_64
timestamp 1667941163
transform 1 0 6992 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_76
timestamp 1667941163
transform 1 0 8096 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_88
timestamp 1667941163
transform 1 0 9200 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_100
timestamp 1667941163
transform 1 0 10304 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_152
timestamp 1667941163
transform 1 0 15088 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_159
timestamp 1667941163
transform 1 0 15732 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_214
timestamp 1667941163
transform 1 0 20792 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1667941163
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_233
timestamp 1667941163
transform 1 0 22540 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_265
timestamp 1667941163
transform 1 0 25484 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_269
timestamp 1667941163
transform 1 0 25852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1667941163
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_345
timestamp 1667941163
transform 1 0 32844 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_350
timestamp 1667941163
transform 1 0 33304 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_362
timestamp 1667941163
transform 1 0 34408 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_374
timestamp 1667941163
transform 1 0 35512 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_386
timestamp 1667941163
transform 1 0 36616 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_57
timestamp 1667941163
transform 1 0 6348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_61
timestamp 1667941163
transform 1 0 6716 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_73
timestamp 1667941163
transform 1 0 7820 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_81
timestamp 1667941163
transform 1 0 8556 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_174
timestamp 1667941163
transform 1 0 17112 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_181
timestamp 1667941163
transform 1 0 17756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_193
timestamp 1667941163
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_47
timestamp 1667941163
transform 1 0 5428 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1667941163
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_174
timestamp 1667941163
transform 1 0 17112 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_186
timestamp 1667941163
transform 1 0 18216 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_198
timestamp 1667941163
transform 1 0 19320 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_210
timestamp 1667941163
transform 1 0 20424 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1667941163
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_401
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_20
timestamp 1667941163
transform 1 0 2944 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_393
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_21
timestamp 1667941163
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_33
timestamp 1667941163
transform 1 0 4140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_45
timestamp 1667941163
transform 1 0 5244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1667941163
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_400
timestamp 1667941163
transform 1 0 37904 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_406
timestamp 1667941163
transform 1 0 38456 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_16
timestamp 1667941163
transform 1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_43
timestamp 1667941163
transform 1 0 5060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_49
timestamp 1667941163
transform 1 0 5612 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1667941163
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_65
timestamp 1667941163
transform 1 0 7084 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_69
timestamp 1667941163
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1667941163
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_104
timestamp 1667941163
transform 1 0 10672 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_118
timestamp 1667941163
transform 1 0 11960 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1667941163
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_149
timestamp 1667941163
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_203
timestamp 1667941163
transform 1 0 19780 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_211
timestamp 1667941163
transform 1 0 20516 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_216
timestamp 1667941163
transform 1 0 20976 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_233
timestamp 1667941163
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1667941163
transform 1 0 26220 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1667941163
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_286
timestamp 1667941163
transform 1 0 27416 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_298
timestamp 1667941163
transform 1 0 28520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1667941163
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_342
timestamp 1667941163
transform 1 0 32568 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_356
timestamp 1667941163
transform 1 0 33856 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_382
timestamp 1667941163
transform 1 0 36248 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_386
timestamp 1667941163
transform 1 0 36616 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0416_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform -1 0 5428 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform -1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform -1 0 17664 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform -1 0 18952 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform -1 0 7360 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform -1 0 8648 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform -1 0 11960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform -1 0 13616 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 6992 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform -1 0 6716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform -1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform -1 0 21252 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 23920 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform -1 0 23092 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 23460 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 16836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 20700 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 20056 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform -1 0 16560 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 17480 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 10028 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 14444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform -1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform -1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 12972 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform -1 0 11224 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 13524 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform -1 0 8648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform -1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform -1 0 7176 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1667941163
transform 1 0 10304 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1667941163
transform 1 0 11592 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0454_
timestamp 1667941163
transform -1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1667941163
transform -1 0 8648 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform -1 0 13248 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform -1 0 14352 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 12328 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform -1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform -1 0 21252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 19596 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform -1 0 20516 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform -1 0 20516 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform -1 0 22356 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 23368 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform -1 0 4232 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 7728 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform -1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform -1 0 14628 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 4416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform -1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform -1 0 5428 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform -1 0 5152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform -1 0 7360 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform -1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0480_
timestamp 1667941163
transform 1 0 24380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1667941163
transform 1 0 23736 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 8004 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 9108 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0486_
timestamp 1667941163
transform -1 0 8924 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1667941163
transform 1 0 9752 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0488_
timestamp 1667941163
transform 1 0 7176 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1667941163
transform 1 0 6532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform -1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 7268 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1667941163
transform -1 0 6072 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0493_
timestamp 1667941163
transform -1 0 6072 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1667941163
transform -1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0495_
timestamp 1667941163
transform -1 0 14536 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform -1 0 4600 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 5152 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1667941163
transform 1 0 4324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0499_
timestamp 1667941163
transform 1 0 3036 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0500_
timestamp 1667941163
transform 1 0 4968 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0501_
timestamp 1667941163
transform 1 0 4232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 23920 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform -1 0 21712 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1667941163
transform 1 0 23276 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0505_
timestamp 1667941163
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1667941163
transform -1 0 23000 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 23460 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform -1 0 4232 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0510_
timestamp 1667941163
transform -1 0 12880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0511_
timestamp 1667941163
transform -1 0 13248 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0512_
timestamp 1667941163
transform -1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1667941163
transform 1 0 17848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 17296 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform -1 0 4416 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform -1 0 16376 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1667941163
transform -1 0 17572 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 16192 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1667941163
transform -1 0 14168 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0521_
timestamp 1667941163
transform 1 0 14628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0522_
timestamp 1667941163
transform -1 0 13248 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform -1 0 21528 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform -1 0 20424 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform -1 0 21712 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0526_
timestamp 1667941163
transform 1 0 22080 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 17112 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0530_
timestamp 1667941163
transform -1 0 21528 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1667941163
transform 1 0 23092 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform -1 0 19688 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 13340 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 18124 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0535_
timestamp 1667941163
transform -1 0 17756 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform -1 0 20240 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1667941163
transform 1 0 20056 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform -1 0 18952 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0539_
timestamp 1667941163
transform -1 0 19136 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0540_
timestamp 1667941163
transform 1 0 19504 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 17296 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 23736 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 21344 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0544_
timestamp 1667941163
transform 1 0 21252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform -1 0 18768 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1667941163
transform 1 0 18584 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform -1 0 19780 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1667941163
transform 1 0 23276 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1667941163
transform 1 0 17112 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1667941163
transform -1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 13064 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform -1 0 12512 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1667941163
transform 1 0 16100 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0558_
timestamp 1667941163
transform -1 0 15824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 3956 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 19136 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 20516 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1667941163
transform -1 0 18400 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0564_
timestamp 1667941163
transform -1 0 6992 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 14996 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1667941163
transform -1 0 17020 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform -1 0 18676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 10672 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1667941163
transform 1 0 14260 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0571_
timestamp 1667941163
transform -1 0 13800 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 13892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform -1 0 13524 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0575_
timestamp 1667941163
transform -1 0 17112 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1667941163
transform 1 0 20332 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 15364 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 13432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1667941163
transform 1 0 14720 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform -1 0 13616 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1667941163
transform -1 0 15180 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 13984 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0584_
timestamp 1667941163
transform 1 0 15456 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1667941163
transform -1 0 13800 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 17204 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1667941163
transform 1 0 17664 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0589_
timestamp 1667941163
transform 1 0 17204 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0590_
timestamp 1667941163
transform -1 0 19780 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1667941163
transform 1 0 19596 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform -1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0593_
timestamp 1667941163
transform 1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1667941163
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1667941163
transform -1 0 6072 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 1667941163
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1667941163
transform -1 0 15732 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 14720 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1667941163
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1667941163
transform -1 0 6992 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 23368 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1667941163
transform 1 0 25760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0607_
timestamp 1667941163
transform 1 0 25208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1667941163
transform -1 0 24380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0609_
timestamp 1667941163
transform 1 0 25300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0611_
timestamp 1667941163
transform -1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1667941163
transform 1 0 24748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform -1 0 26312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform -1 0 25668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1667941163
transform -1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0616_
timestamp 1667941163
transform 1 0 26404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1667941163
transform 1 0 25668 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 26128 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0620_
timestamp 1667941163
transform 1 0 25668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1667941163
transform 1 0 25024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 21988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1667941163
transform -1 0 20976 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0625_
timestamp 1667941163
transform 1 0 20792 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1667941163
transform 1 0 15456 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1667941163
transform -1 0 13800 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 19780 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1667941163
transform -1 0 22264 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform -1 0 3220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1667941163
transform -1 0 19780 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0634_
timestamp 1667941163
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1667941163
transform -1 0 2576 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 21160 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0638_
timestamp 1667941163
transform 1 0 21252 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1667941163
transform -1 0 20884 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 9292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1667941163
transform 1 0 10948 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1667941163
transform -1 0 9936 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1667941163
transform -1 0 11960 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1667941163
transform -1 0 14260 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 15456 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0647_
timestamp 1667941163
transform -1 0 16100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1667941163
transform 1 0 15732 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 4784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1667941163
transform 1 0 10488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1667941163
transform -1 0 10212 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1667941163
transform 1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1667941163
transform -1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 1667941163
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform -1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1667941163
transform -1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0661_
timestamp 1667941163
transform 1 0 13064 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1667941163
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1667941163
transform 1 0 15456 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0665_
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1667941163
transform 1 0 15272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 10580 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform -1 0 11960 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1667941163
transform -1 0 1932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0670_
timestamp 1667941163
transform -1 0 8004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1667941163
transform -1 0 12144 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1667941163
transform -1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform -1 0 16376 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0674_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0675_
timestamp 1667941163
transform -1 0 15824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 2300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 9016 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1667941163
transform -1 0 8648 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0679_
timestamp 1667941163
transform -1 0 10212 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1667941163
transform -1 0 6808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1667941163
transform -1 0 11408 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 9200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0683_
timestamp 1667941163
transform 1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1667941163
transform -1 0 3220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 14352 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 16100 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1667941163
transform 1 0 18216 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1667941163
transform 1 0 17480 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1667941163
transform -1 0 13800 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0690_
timestamp 1667941163
transform -1 0 14812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 19412 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0692_
timestamp 1667941163
transform -1 0 19964 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0693_
timestamp 1667941163
transform -1 0 20608 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 14168 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform -1 0 14996 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0696_
timestamp 1667941163
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1667941163
transform -1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0699_
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1667941163
transform -1 0 12880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1667941163
transform -1 0 16468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0702_
timestamp 1667941163
transform -1 0 16376 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 10488 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 17112 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 16652 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 1667941163
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1667941163
transform -1 0 14628 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0708_
timestamp 1667941163
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1667941163
transform -1 0 8004 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform -1 0 30820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform -1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform -1 0 27416 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform -1 0 10120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform -1 0 33856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 6440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform -1 0 28244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 18584 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform -1 0 25484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform -1 0 8372 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform -1 0 8648 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform -1 0 10120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 16376 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 6716 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform -1 0 20056 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform -1 0 31188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform -1 0 34040 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform -1 0 12236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform -1 0 33764 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 29348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform -1 0 29992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 29532 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform -1 0 32292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform -1 0 35144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 29716 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 9200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 29992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform -1 0 34776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 19596 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 14260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 17020 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform -1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform -1 0 23368 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform -1 0 33304 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 17204 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform -1 0 11960 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform -1 0 34224 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform -1 0 30636 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform -1 0 35328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform -1 0 30820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 35604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 7176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 27416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform -1 0 20792 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 33304 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 29624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 25116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform -1 0 34500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform -1 0 4232 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform -1 0 25576 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 1840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 36800 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 6532 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform -1 0 6348 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform -1 0 9936 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform -1 0 34408 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform -1 0 13156 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform -1 0 29440 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 4324 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform -1 0 30820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 20792 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 6624 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 7268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform -1 0 9200 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 14168 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform -1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform -1 0 29348 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 16836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform -1 0 30360 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 24564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform -1 0 24748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform -1 0 3956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 10304 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0804_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37536 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 9108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0806_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 9660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0807_
timestamp 1667941163
transform -1 0 2852 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform -1 0 2484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform -1 0 3496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform -1 0 2392 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 7820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform -1 0 6808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0818_
timestamp 1667941163
transform -1 0 2668 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform -1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform -1 0 2576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform -1 0 5152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 2944 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 6532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform -1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0829_
timestamp 1667941163
transform -1 0 2852 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform -1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform -1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform -1 0 4692 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform -1 0 2576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform -1 0 6072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0840_
timestamp 1667941163
transform -1 0 2760 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 4140 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 4600 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform -1 0 4232 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 1932 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform -1 0 1840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 3496 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform -1 0 3496 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 4876 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 2576 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1667941163
transform 1 0 2392 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0851_
timestamp 1667941163
transform -1 0 8004 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 4232 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 2392 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 4600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform -1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1667941163
transform 1 0 2668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0862_
timestamp 1667941163
transform -1 0 8004 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1667941163
transform 1 0 3956 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1667941163
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1667941163
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1667941163
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1667941163
transform 1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1667941163
transform -1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1667941163
transform 1 0 3956 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0873_
timestamp 1667941163
transform -1 0 8004 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1667941163
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1667941163
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1667941163
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1667941163
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1667941163
transform 1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1667941163
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1667941163
transform 1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1667941163
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1667941163
transform 1 0 3128 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1667941163
transform 1 0 2944 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1667941163
transform 1 0 2760 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1667941163
transform 1 0 6348 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1667941163
transform 1 0 4968 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1667941163
transform 1 0 5060 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1667941163
transform 1 0 5704 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0890_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11316 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0891_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5520 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 1656 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0893_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 3496 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1667941163
transform -1 0 3496 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0895_
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0896_
timestamp 1667941163
transform -1 0 9476 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0897_
timestamp 1667941163
transform 1 0 5244 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0898_
timestamp 1667941163
transform 1 0 4600 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0899_
timestamp 1667941163
transform 1 0 2024 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform -1 0 3496 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0901_
timestamp 1667941163
transform -1 0 5980 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1667941163
transform 1 0 5060 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0903_
timestamp 1667941163
transform 1 0 1564 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0904_
timestamp 1667941163
transform -1 0 3496 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0905_
timestamp 1667941163
transform -1 0 7728 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 1564 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0907_
timestamp 1667941163
transform -1 0 4508 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 2208 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0909_
timestamp 1667941163
transform -1 0 4232 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0910_
timestamp 1667941163
transform 1 0 1564 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0911_
timestamp 1667941163
transform 1 0 4140 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 4048 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0913_
timestamp 1667941163
transform 1 0 2852 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 1656 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0915_
timestamp 1667941163
transform -1 0 8464 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0916_
timestamp 1667941163
transform 1 0 1656 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0917_
timestamp 1667941163
transform -1 0 3680 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform -1 0 6072 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0919_
timestamp 1667941163
transform 1 0 3956 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1667941163
transform -1 0 5796 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0921_
timestamp 1667941163
transform 1 0 4784 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 1656 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0923_
timestamp 1667941163
transform -1 0 3680 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform -1 0 3404 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0925_
timestamp 1667941163
transform -1 0 5704 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0926_
timestamp 1667941163
transform -1 0 3496 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0927_
timestamp 1667941163
transform -1 0 6716 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 1656 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0929_
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 8832 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0931_
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0932_
timestamp 1667941163
transform -1 0 6992 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0933_
timestamp 1667941163
transform -1 0 9476 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0934_
timestamp 1667941163
transform -1 0 9200 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 9016 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0936_
timestamp 1667941163
transform -1 0 6072 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform -1 0 8648 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform -1 0 6072 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform -1 0 8648 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 7360 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1667941163
transform 1 0 4600 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0942_
timestamp 1667941163
transform -1 0 8648 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1667941163
transform -1 0 10948 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0944_
timestamp 1667941163
transform -1 0 7360 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0945_
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0946_
timestamp 1667941163
transform -1 0 10948 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 1656 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform -1 0 8648 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1667941163
transform -1 0 7544 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform -1 0 10948 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1667941163
transform 1 0 11684 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 9108 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0954_
timestamp 1667941163
transform 1 0 4232 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0955_
timestamp 1667941163
transform -1 0 6072 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1667941163
transform -1 0 10672 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1667941163
transform -1 0 9568 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0959_
timestamp 1667941163
transform -1 0 8096 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0960_
timestamp 1667941163
transform 1 0 6532 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0961_
timestamp 1667941163
transform -1 0 8372 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0962_
timestamp 1667941163
transform -1 0 10948 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0963_
timestamp 1667941163
transform -1 0 10948 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0964_
timestamp 1667941163
transform 1 0 9108 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0965_
timestamp 1667941163
transform -1 0 9568 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform -1 0 33580 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform -1 0 37628 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 15456 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 2852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform -1 0 22908 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform -1 0 35604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform -1 0 33120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform -1 0 36340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 6440 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 7176 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform -1 0 17756 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform -1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform -1 0 35144 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform -1 0 34040 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform -1 0 35144 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform -1 0 35420 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform -1 0 27416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 11684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform -1 0 35144 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 5704 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1667941163
transform -1 0 37720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 3956 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1667941163
transform -1 0 25760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform -1 0 34408 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 6716 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 14076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform -1 0 17112 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform -1 0 20424 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform -1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 4508 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1667941163
transform -1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform -1 0 34040 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1042_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15364 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1043_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1043__100 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1044_
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1045_
timestamp 1667941163
transform 1 0 18124 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1046_
timestamp 1667941163
transform -1 0 18676 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1047_
timestamp 1667941163
transform 1 0 10672 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1048_
timestamp 1667941163
transform -1 0 16836 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1049_
timestamp 1667941163
transform 1 0 12512 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1049__101
timestamp 1667941163
transform -1 0 12512 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1050_
timestamp 1667941163
transform 1 0 12972 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 14720 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1052_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1053_
timestamp 1667941163
transform 1 0 14444 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1054_
timestamp 1667941163
transform -1 0 15272 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1055__102
timestamp 1667941163
transform 1 0 21160 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1055_
timestamp 1667941163
transform -1 0 21160 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1056_
timestamp 1667941163
transform 1 0 17480 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1057_
timestamp 1667941163
transform -1 0 15364 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1058_
timestamp 1667941163
transform -1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1059_
timestamp 1667941163
transform 1 0 17388 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1060_
timestamp 1667941163
transform 1 0 11684 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1061_
timestamp 1667941163
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1061__103
timestamp 1667941163
transform -1 0 5060 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1062_
timestamp 1667941163
transform 1 0 10488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1063_
timestamp 1667941163
transform 1 0 11316 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1064_
timestamp 1667941163
transform 1 0 12420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1065_
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1066_
timestamp 1667941163
transform -1 0 12512 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1067_
timestamp 1667941163
transform 1 0 16100 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1067__104
timestamp 1667941163
transform -1 0 15732 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1068_
timestamp 1667941163
transform 1 0 13892 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1069_
timestamp 1667941163
transform -1 0 12512 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1070_
timestamp 1667941163
transform -1 0 16744 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1071_
timestamp 1667941163
transform 1 0 11592 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1072_
timestamp 1667941163
transform 1 0 15364 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1073_
timestamp 1667941163
transform 1 0 14996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1073__105
timestamp 1667941163
transform 1 0 14996 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1074_
timestamp 1667941163
transform 1 0 12880 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1075_
timestamp 1667941163
transform 1 0 14444 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 14904 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1077_
timestamp 1667941163
transform 1 0 11316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1078_
timestamp 1667941163
transform 1 0 10396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1079_
timestamp 1667941163
transform 1 0 10304 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1079__106
timestamp 1667941163
transform 1 0 10304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1080_
timestamp 1667941163
transform 1 0 11316 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1081_
timestamp 1667941163
transform 1 0 11684 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1082_
timestamp 1667941163
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1083_
timestamp 1667941163
transform 1 0 10028 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1084_
timestamp 1667941163
transform -1 0 15364 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1085__107
timestamp 1667941163
transform 1 0 15456 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1085_
timestamp 1667941163
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1086_
timestamp 1667941163
transform 1 0 11684 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1087_
timestamp 1667941163
transform 1 0 11868 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1088_
timestamp 1667941163
transform -1 0 17572 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1089_
timestamp 1667941163
transform 1 0 11224 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1090_
timestamp 1667941163
transform -1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1091__108
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1091_
timestamp 1667941163
transform -1 0 22080 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1092_
timestamp 1667941163
transform -1 0 18952 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1093_
timestamp 1667941163
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1094_
timestamp 1667941163
transform -1 0 22080 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1095_
timestamp 1667941163
transform 1 0 10488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform -1 0 16100 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1097__109
timestamp 1667941163
transform 1 0 22632 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1097_
timestamp 1667941163
transform -1 0 21528 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1098_
timestamp 1667941163
transform -1 0 20240 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1099_
timestamp 1667941163
transform -1 0 16376 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1100_
timestamp 1667941163
transform -1 0 21528 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1101_
timestamp 1667941163
transform -1 0 20148 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1102_
timestamp 1667941163
transform 1 0 24932 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1103__110
timestamp 1667941163
transform 1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1103_
timestamp 1667941163
transform -1 0 25300 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1104_
timestamp 1667941163
transform -1 0 24932 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1105_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1106_
timestamp 1667941163
transform -1 0 24564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1107_
timestamp 1667941163
transform 1 0 23644 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1108_
timestamp 1667941163
transform 1 0 23276 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1109_
timestamp 1667941163
transform -1 0 22724 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1109__111
timestamp 1667941163
transform 1 0 22632 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1110_
timestamp 1667941163
transform -1 0 23828 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1111_
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1112_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1113_
timestamp 1667941163
transform -1 0 23828 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1114_
timestamp 1667941163
transform 1 0 16468 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1115__112
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1116_
timestamp 1667941163
transform -1 0 13432 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1117_
timestamp 1667941163
transform 1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1118_
timestamp 1667941163
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1119_
timestamp 1667941163
transform 1 0 11868 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1120_
timestamp 1667941163
transform 1 0 19320 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1121_
timestamp 1667941163
transform -1 0 18952 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1121__113
timestamp 1667941163
transform -1 0 18952 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1122_
timestamp 1667941163
transform 1 0 17112 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1123_
timestamp 1667941163
transform 1 0 18124 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1124_
timestamp 1667941163
transform 1 0 17664 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1125_
timestamp 1667941163
transform -1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1126_
timestamp 1667941163
transform 1 0 16744 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1127_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1127__114
timestamp 1667941163
transform -1 0 12972 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1128_
timestamp 1667941163
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1129_
timestamp 1667941163
transform 1 0 15088 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1130_
timestamp 1667941163
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1131_
timestamp 1667941163
transform -1 0 14352 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 15364 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1133_
timestamp 1667941163
transform -1 0 17572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1133__115
timestamp 1667941163
transform -1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1134_
timestamp 1667941163
transform -1 0 16100 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 13616 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1136_
timestamp 1667941163
transform -1 0 16376 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1137_
timestamp 1667941163
transform 1 0 11868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform -1 0 13800 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1139_
timestamp 1667941163
transform 1 0 18952 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1139__116
timestamp 1667941163
transform -1 0 18032 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1140_
timestamp 1667941163
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform -1 0 13616 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1142_
timestamp 1667941163
transform 1 0 17848 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1143_
timestamp 1667941163
transform -1 0 20148 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform -1 0 13800 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1145__117
timestamp 1667941163
transform 1 0 16192 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1145_
timestamp 1667941163
transform 1 0 16100 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1146_
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform -1 0 13616 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1148_
timestamp 1667941163
transform 1 0 14996 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1149_
timestamp 1667941163
transform -1 0 18768 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1150_
timestamp 1667941163
transform -1 0 18308 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1151_
timestamp 1667941163
transform -1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1151__118
timestamp 1667941163
transform 1 0 21620 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1152_
timestamp 1667941163
transform -1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform -1 0 18216 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1154_
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1155_
timestamp 1667941163
transform -1 0 20792 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1157__119
timestamp 1667941163
transform 1 0 20148 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1157_
timestamp 1667941163
transform -1 0 18952 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1158_
timestamp 1667941163
transform 1 0 18032 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1159_
timestamp 1667941163
transform 1 0 18768 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1160_
timestamp 1667941163
transform 1 0 18400 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1161_
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 20700 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1163_
timestamp 1667941163
transform 1 0 19964 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1163__120
timestamp 1667941163
transform -1 0 18952 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1164_
timestamp 1667941163
transform -1 0 21528 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 21068 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1166_
timestamp 1667941163
transform 1 0 19320 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1167_
timestamp 1667941163
transform -1 0 20424 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 16008 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1169__121
timestamp 1667941163
transform -1 0 12328 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1169_
timestamp 1667941163
transform 1 0 15272 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1170_
timestamp 1667941163
transform -1 0 18032 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1171_
timestamp 1667941163
transform -1 0 17664 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1172_
timestamp 1667941163
transform 1 0 14536 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1173_
timestamp 1667941163
transform 1 0 11684 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1174_
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1174__122
timestamp 1667941163
transform 1 0 17940 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 13892 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1176_
timestamp 1667941163
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1177_
timestamp 1667941163
transform 1 0 12972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1178__123
timestamp 1667941163
transform 1 0 23920 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1178_
timestamp 1667941163
transform -1 0 22908 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1179_
timestamp 1667941163
transform -1 0 22724 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1180_
timestamp 1667941163
transform 1 0 22264 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1181_
timestamp 1667941163
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1182_
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1182__124
timestamp 1667941163
transform -1 0 2852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 3036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1184_
timestamp 1667941163
transform 1 0 4232 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform -1 0 9016 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1186_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16376 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1186__125
timestamp 1667941163
transform -1 0 16376 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1187_
timestamp 1667941163
transform 1 0 6440 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1188_
timestamp 1667941163
transform 1 0 10028 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1189_
timestamp 1667941163
transform 1 0 7636 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1190__126
timestamp 1667941163
transform 1 0 5888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1190_
timestamp 1667941163
transform 1 0 5888 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform -1 0 8372 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1192_
timestamp 1667941163
transform -1 0 7636 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform -1 0 8280 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1194_
timestamp 1667941163
transform -1 0 23552 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1194__127
timestamp 1667941163
transform -1 0 23368 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1195_
timestamp 1667941163
transform -1 0 23000 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 22632 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1197_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1198__128
timestamp 1667941163
transform -1 0 11224 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1198_
timestamp 1667941163
transform 1 0 11868 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1199_
timestamp 1667941163
transform 1 0 11868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1200_
timestamp 1667941163
transform 1 0 12512 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 11684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 14996 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1202__129
timestamp 1667941163
transform -1 0 14536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform 1 0 5336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1204_
timestamp 1667941163
transform 1 0 9844 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1205_
timestamp 1667941163
transform 1 0 7912 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1206__130
timestamp 1667941163
transform -1 0 22448 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1206_
timestamp 1667941163
transform 1 0 22816 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1207_
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1208_
timestamp 1667941163
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 19872 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1210__131
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1210_
timestamp 1667941163
transform 1 0 14260 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1211_
timestamp 1667941163
transform -1 0 14996 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1212_
timestamp 1667941163
transform 1 0 11316 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 15640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1214__132
timestamp 1667941163
transform -1 0 14628 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1215_
timestamp 1667941163
transform 1 0 9108 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1216_
timestamp 1667941163
transform 1 0 14260 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1217_
timestamp 1667941163
transform 1 0 6164 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1218__133
timestamp 1667941163
transform -1 0 12604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1218_
timestamp 1667941163
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1219_
timestamp 1667941163
transform -1 0 18768 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1220_
timestamp 1667941163
transform -1 0 14812 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1221_
timestamp 1667941163
transform -1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1222__134
timestamp 1667941163
transform 1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1222_
timestamp 1667941163
transform -1 0 17112 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1223_
timestamp 1667941163
transform -1 0 18768 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1224_
timestamp 1667941163
transform -1 0 17572 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1225_
timestamp 1667941163
transform -1 0 18860 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1226_
timestamp 1667941163
transform 1 0 22724 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1226__135
timestamp 1667941163
transform 1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1227_
timestamp 1667941163
transform 1 0 19044 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1228_
timestamp 1667941163
transform 1 0 20424 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1229_
timestamp 1667941163
transform -1 0 20516 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1230__136
timestamp 1667941163
transform -1 0 5888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1230_
timestamp 1667941163
transform 1 0 6532 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1231_
timestamp 1667941163
transform -1 0 14904 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1232_
timestamp 1667941163
transform -1 0 7912 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1233_
timestamp 1667941163
transform -1 0 10304 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1234_
timestamp 1667941163
transform 1 0 18768 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1234__137
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1235_
timestamp 1667941163
transform 1 0 18124 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1236_
timestamp 1667941163
transform 1 0 18492 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1237_
timestamp 1667941163
transform 1 0 9108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1667941163
transform -1 0 3496 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1667941163
transform -1 0 4416 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1667941163
transform -1 0 9660 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1667941163
transform 1 0 7820 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1667941163
transform -1 0 3496 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1667941163
transform -1 0 3496 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1667941163
transform 1 0 6808 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1667941163
transform -1 0 10948 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform -1 0 1840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 38088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 38088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform -1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 38088 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform -1 0 1840 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 38088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform -1 0 3220 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform -1 0 1840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 36708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform -1 0 1840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 38088 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 20700 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform -1 0 13248 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 38088 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 38088 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform -1 0 1840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform -1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform -1 0 1840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform -1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform -1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform -1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 36708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform -1 0 17112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 36708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12328 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 38088 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 30452 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform -1 0 2576 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform -1 0 1840 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 38088 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 4324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform -1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform -1 0 15272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform -1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform -1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform -1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform -1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform -1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform -1 0 5612 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 37996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 37996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 18584 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform -1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform -1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform -1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform -1 0 1932 0 -1 36992
box -38 -48 406 592
<< labels >>
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 ccff_head
port 0 nsew signal input
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 2 nsew signal input
flabel metal3 s 39200 11568 39800 11688 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 3 nsew signal input
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 4 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 5 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_left_in[13]
port 6 nsew signal input
flabel metal2 s 15474 200 15530 800 0 FreeSans 224 90 0 0 chanx_left_in[14]
port 7 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 8 nsew signal input
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 9 nsew signal input
flabel metal3 s 39200 31288 39800 31408 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 10 nsew signal input
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_left_in[18]
port 11 nsew signal input
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_left_in[1]
port 12 nsew signal input
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 13 nsew signal input
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chanx_left_in[3]
port 14 nsew signal input
flabel metal3 s 39200 19728 39800 19848 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 15 nsew signal input
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 16 nsew signal input
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 17 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 18 nsew signal input
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 19 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 20 nsew signal input
flabel metal3 s 39200 34688 39800 34808 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 21 nsew signal tristate
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 22 nsew signal tristate
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chanx_left_out[11]
port 23 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 24 nsew signal tristate
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_left_out[13]
port 25 nsew signal tristate
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 26 nsew signal tristate
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 27 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 28 nsew signal tristate
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 29 nsew signal tristate
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 30 nsew signal tristate
flabel metal3 s 39200 36728 39800 36848 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 31 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 32 nsew signal tristate
flabel metal2 s 23846 39200 23902 39800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 33 nsew signal tristate
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 34 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 35 nsew signal tristate
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 36 nsew signal tristate
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 37 nsew signal tristate
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 38 nsew signal tristate
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 39 nsew signal tristate
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal2 s 20626 39200 20682 39800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal3 s 200 2728 800 2848 0 FreeSans 480 0 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal2 s 34794 39200 34850 39800 0 FreeSans 224 90 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal2 s 2594 200 2650 800 0 FreeSans 224 90 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal3 s 200 16328 800 16448 0 FreeSans 480 0 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal3 s 200 8168 800 8288 0 FreeSans 480 0 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal3 s 200 12928 800 13048 0 FreeSans 480 0 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 78 nsew signal input
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 79 nsew signal input
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 80 nsew signal input
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 81 nsew signal input
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 82 nsew signal input
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 83 nsew signal input
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 84 nsew signal input
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 85 nsew signal input
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 86 nsew signal input
flabel metal2 s 7746 200 7802 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 87 nsew signal input
flabel metal2 s 12254 200 12310 800 0 FreeSans 224 90 0 0 pReset
port 88 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 prog_clk
port 89 nsew signal input
flabel metal3 s 39200 23128 39800 23248 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 90 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 91 nsew signal input
flabel metal2 s 31574 39200 31630 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 92 nsew signal input
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 93 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 94 nsew signal input
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 95 nsew signal input
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 96 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 97 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 98 nsew signal input
flabel metal3 s 39200 18368 39800 18488 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 99 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 5803 16490 5803 16490 0 _0000_
rlabel metal1 4738 9078 4738 9078 0 _0001_
rlabel metal1 4745 16150 4745 16150 0 _0002_
rlabel metal1 3411 16490 3411 16490 0 _0003_
rlabel metal2 2622 22950 2622 22950 0 _0004_
rlabel metal2 2990 7106 2990 7106 0 _0005_
rlabel metal1 4094 6970 4094 6970 0 _0006_
rlabel metal1 4462 7514 4462 7514 0 _0007_
rlabel metal1 4692 5882 4692 5882 0 _0008_
rlabel metal1 4830 21046 4830 21046 0 _0009_
rlabel metal1 5198 27302 5198 27302 0 _0010_
rlabel metal1 3365 18326 3365 18326 0 _0011_
rlabel metal1 2109 21590 2109 21590 0 _0012_
rlabel metal1 1833 17578 1833 17578 0 _0013_
rlabel metal1 4133 19414 4133 19414 0 _0014_
rlabel metal2 2714 11135 2714 11135 0 _0015_
rlabel metal1 5145 17578 5145 17578 0 _0016_
rlabel metal2 2714 23800 2714 23800 0 _0017_
rlabel metal1 1833 13974 1833 13974 0 _0018_
rlabel metal1 10679 15062 10679 15062 0 _0019_
rlabel metal2 8786 22117 8786 22117 0 _0020_
rlabel metal2 6026 23545 6026 23545 0 _0021_
rlabel metal2 4784 21148 4784 21148 0 _0022_
rlabel metal1 5336 3638 5336 3638 0 _0023_
rlabel via2 2714 6851 2714 6851 0 _0024_
rlabel metal1 2346 3706 2346 3706 0 _0025_
rlabel metal1 5290 4794 5290 4794 0 _0026_
rlabel metal1 3174 25330 3174 25330 0 _0027_
rlabel metal1 4922 5134 4922 5134 0 _0028_
rlabel metal1 7905 17238 7905 17238 0 _0029_
rlabel metal1 4554 23562 4554 23562 0 _0030_
rlabel metal1 6394 22066 6394 22066 0 _0031_
rlabel via2 1794 9469 1794 9469 0 _0032_
rlabel metal2 3450 4828 3450 4828 0 _0033_
rlabel metal1 7728 9486 7728 9486 0 _0034_
rlabel metal1 1932 15130 1932 15130 0 _0035_
rlabel metal2 7314 10166 7314 10166 0 _0036_
rlabel metal1 6072 9486 6072 9486 0 _0037_
rlabel metal1 4968 21862 4968 21862 0 _0038_
rlabel metal1 2990 3128 2990 3128 0 _0039_
rlabel metal1 6072 4046 6072 4046 0 _0040_
rlabel via3 13133 16660 13133 16660 0 _0041_
rlabel via3 10051 12852 10051 12852 0 _0042_
rlabel metal2 5014 6392 5014 6392 0 _0043_
rlabel metal1 3174 6766 3174 6766 0 _0044_
rlabel metal1 6394 9350 6394 9350 0 _0045_
rlabel metal1 2599 7310 2599 7310 0 _0046_
rlabel metal1 5704 25398 5704 25398 0 _0047_
rlabel metal2 5198 23562 5198 23562 0 _0048_
rlabel via3 7981 15164 7981 15164 0 _0049_
rlabel metal3 6555 13668 6555 13668 0 _0050_
rlabel metal1 7268 29478 7268 29478 0 _0051_
rlabel metal3 7291 29036 7291 29036 0 _0052_
rlabel metal2 9890 21461 9890 21461 0 _0053_
rlabel metal1 7767 21590 7767 21590 0 _0054_
rlabel metal2 12650 16439 12650 16439 0 _0055_
rlabel metal2 6992 21012 6992 21012 0 _0056_
rlabel metal2 3082 7174 3082 7174 0 _0057_
rlabel metal1 3450 6426 3450 6426 0 _0058_
rlabel metal1 1978 18768 1978 18768 0 _0059_
rlabel metal2 4876 13668 4876 13668 0 _0060_
rlabel metal1 8004 8602 8004 8602 0 _0061_
rlabel metal1 5980 11866 5980 11866 0 _0062_
rlabel metal2 8510 9520 8510 9520 0 _0063_
rlabel metal1 6164 8602 6164 8602 0 _0064_
rlabel metal1 1748 4794 1748 4794 0 _0065_
rlabel metal1 4087 12886 4087 12886 0 _0066_
rlabel metal2 5842 6256 5842 6256 0 _0067_
rlabel metal1 1610 4046 1610 4046 0 _0068_
rlabel metal2 2622 22005 2622 22005 0 _0069_
rlabel metal1 5973 14314 5973 14314 0 _0070_
rlabel metal1 4055 23018 4055 23018 0 _0071_
rlabel metal1 3128 26758 3128 26758 0 _0072_
rlabel metal3 5267 20740 5267 20740 0 _0073_
rlabel metal1 3128 7514 3128 7514 0 _0074_
rlabel metal1 3503 15402 3503 15402 0 _0075_
rlabel metal1 9982 20502 9982 20502 0 _0076_
rlabel metal1 18354 24174 18354 24174 0 _0077_
rlabel metal1 13386 26928 13386 26928 0 _0078_
rlabel metal2 6486 25466 6486 25466 0 _0079_
rlabel metal2 23414 14195 23414 14195 0 _0080_
rlabel metal2 23690 20876 23690 20876 0 _0081_
rlabel metal2 20102 26486 20102 26486 0 _0082_
rlabel metal2 17710 27914 17710 27914 0 _0083_
rlabel metal1 17204 16762 17204 16762 0 _0084_
rlabel metal2 11730 24718 11730 24718 0 _0085_
rlabel metal2 8602 6086 8602 6086 0 _0086_
rlabel metal1 9430 12886 9430 12886 0 _0087_
rlabel metal2 8418 14858 8418 14858 0 _0088_
rlabel metal1 13662 12818 13662 12818 0 _0089_
rlabel metal1 10810 24174 10810 24174 0 _0090_
rlabel metal2 20470 11526 20470 11526 0 _0091_
rlabel metal1 23598 11696 23598 11696 0 _0092_
rlabel metal1 5520 25874 5520 25874 0 _0093_
rlabel metal2 14398 11322 14398 11322 0 _0094_
rlabel metal1 4830 20026 4830 20026 0 _0095_
rlabel metal1 5382 19958 5382 19958 0 _0096_
rlabel metal1 24196 16082 24196 16082 0 _0097_
rlabel metal1 25024 14382 25024 14382 0 _0098_
rlabel metal2 9982 26554 9982 26554 0 _0099_
rlabel metal1 6992 27438 6992 27438 0 _0100_
rlabel metal1 5934 24922 5934 24922 0 _0101_
rlabel metal2 14306 12257 14306 12257 0 _0102_
rlabel metal1 3266 25908 3266 25908 0 _0103_
rlabel metal1 4922 26554 4922 26554 0 _0104_
rlabel metal1 23092 12818 23092 12818 0 _0105_
rlabel metal1 23322 11594 23322 11594 0 _0106_
rlabel metal1 12926 10778 12926 10778 0 _0107_
rlabel metal2 18078 10948 18078 10948 0 _0108_
rlabel metal1 16836 17034 16836 17034 0 _0109_
rlabel metal2 13938 23868 13938 23868 0 _0110_
rlabel metal1 13892 18938 13892 18938 0 _0111_
rlabel metal1 21873 19958 21873 19958 0 _0112_
rlabel metal1 22494 14994 22494 14994 0 _0113_
rlabel metal1 21528 14790 21528 14790 0 _0114_
rlabel metal1 17848 21658 17848 21658 0 _0115_
rlabel metal2 20194 21828 20194 21828 0 _0116_
rlabel metal1 19412 20434 19412 20434 0 _0117_
rlabel metal1 21436 18938 21436 18938 0 _0118_
rlabel metal2 18722 11526 18722 11526 0 _0119_
rlabel metal1 22264 12818 22264 12818 0 _0120_
rlabel metal1 14674 20366 14674 20366 0 _0121_
rlabel metal2 12282 26826 12282 26826 0 _0122_
rlabel metal2 15594 26554 15594 26554 0 _0123_
rlabel metal2 20562 23562 20562 23562 0 _0124_
rlabel metal1 6762 15980 6762 15980 0 _0125_
rlabel metal1 18400 13906 18400 13906 0 _0126_
rlabel metal2 14306 19652 14306 19652 0 _0127_
rlabel metal1 13294 23664 13294 23664 0 _0128_
rlabel metal1 20516 23698 20516 23698 0 _0129_
rlabel metal1 14904 9690 14904 9690 0 _0130_
rlabel metal1 14950 19380 14950 19380 0 _0131_
rlabel metal1 14536 21862 14536 21862 0 _0132_
rlabel metal1 17572 9690 17572 9690 0 _0133_
rlabel metal1 19872 10778 19872 10778 0 _0134_
rlabel metal2 18906 10234 18906 10234 0 _0135_
rlabel metal1 13110 12376 13110 12376 0 _0136_
rlabel metal1 15916 16762 15916 16762 0 _0137_
rlabel metal1 6992 17170 6992 17170 0 _0138_
rlabel metal1 25622 18938 25622 18938 0 _0139_
rlabel metal2 25530 19788 25530 19788 0 _0140_
rlabel metal1 24886 17850 24886 17850 0 _0141_
rlabel metal1 26036 17850 26036 17850 0 _0142_
rlabel metal1 26542 16558 26542 16558 0 _0143_
rlabel metal1 25484 16082 25484 16082 0 _0144_
rlabel metal1 20976 18938 20976 18938 0 _0145_
rlabel metal2 15502 15028 15502 15028 0 _0146_
rlabel metal2 22218 18326 22218 18326 0 _0147_
rlabel metal1 20194 17170 20194 17170 0 _0148_
rlabel metal2 2346 17612 2346 17612 0 _0149_
rlabel metal1 21252 20570 21252 20570 0 _0150_
rlabel metal2 9706 25228 9706 25228 0 _0151_
rlabel metal2 12466 26571 12466 26571 0 _0152_
rlabel metal2 15962 27642 15962 27642 0 _0153_
rlabel metal2 10534 10438 10534 10438 0 _0154_
rlabel metal1 10580 7854 10580 7854 0 _0155_
rlabel metal1 9246 8432 9246 8432 0 _0156_
rlabel metal2 13294 10234 13294 10234 0 _0157_
rlabel metal2 15686 9350 15686 9350 0 _0158_
rlabel metal2 15502 8636 15502 8636 0 _0159_
rlabel metal1 2070 19482 2070 19482 0 _0160_
rlabel metal1 11960 9146 11960 9146 0 _0161_
rlabel metal2 16882 9894 16882 9894 0 _0162_
rlabel metal1 8602 23596 8602 23596 0 _0163_
rlabel metal1 7866 12682 7866 12682 0 _0164_
rlabel metal2 8234 11832 8234 11832 0 _0165_
rlabel metal2 17710 26554 17710 26554 0 _0166_
rlabel metal1 14582 25908 14582 25908 0 _0167_
rlabel metal1 20148 25262 20148 25262 0 _0168_
rlabel metal1 13248 9146 13248 9146 0 _0169_
rlabel metal2 12650 8772 12650 8772 0 _0170_
rlabel metal2 16422 10438 16422 10438 0 _0171_
rlabel metal1 18262 14586 18262 14586 0 _0172_
rlabel metal1 8096 20910 8096 20910 0 _0173_
rlabel metal1 8510 4658 8510 4658 0 _0174_
rlabel metal2 2346 25313 2346 25313 0 _0175_
rlabel metal2 2530 27710 2530 27710 0 _0176_
rlabel metal1 2622 6324 2622 6324 0 _0177_
rlabel metal1 2346 25874 2346 25874 0 _0178_
rlabel metal2 2438 24582 2438 24582 0 _0179_
rlabel metal2 1886 19669 1886 19669 0 _0180_
rlabel metal2 2254 3570 2254 3570 0 _0181_
rlabel metal1 14766 12682 14766 12682 0 _0182_
rlabel metal1 12466 21046 12466 21046 0 _0183_
rlabel metal2 14582 15810 14582 15810 0 _0184_
rlabel metal1 17434 15130 17434 15130 0 _0185_
rlabel metal1 17618 17714 17618 17714 0 _0186_
rlabel metal1 10764 23154 10764 23154 0 _0187_
rlabel metal1 16468 10778 16468 10778 0 _0188_
rlabel metal1 12788 9146 12788 9146 0 _0189_
rlabel metal1 13294 13226 13294 13226 0 _0190_
rlabel metal1 14582 9554 14582 9554 0 _0191_
rlabel metal1 11914 11798 11914 11798 0 _0192_
rlabel metal1 14766 14926 14766 14926 0 _0193_
rlabel metal1 14904 23698 14904 23698 0 _0194_
rlabel metal2 20930 24684 20930 24684 0 _0195_
rlabel metal1 17664 24242 17664 24242 0 _0196_
rlabel metal2 15134 24684 15134 24684 0 _0197_
rlabel metal2 20562 25228 20562 25228 0 _0198_
rlabel metal1 17204 24786 17204 24786 0 _0199_
rlabel metal2 11362 12155 11362 12155 0 _0200_
rlabel metal1 3174 14892 3174 14892 0 _0201_
rlabel metal1 10442 22610 10442 22610 0 _0202_
rlabel metal2 2806 14688 2806 14688 0 _0203_
rlabel metal1 9982 10200 9982 10200 0 _0204_
rlabel metal1 9522 23698 9522 23698 0 _0205_
rlabel metal1 12144 10234 12144 10234 0 _0206_
rlabel metal1 16100 13362 16100 13362 0 _0207_
rlabel metal1 13294 17136 13294 17136 0 _0208_
rlabel metal1 12190 15402 12190 15402 0 _0209_
rlabel metal1 16376 9622 16376 9622 0 _0210_
rlabel metal2 11822 15028 11822 15028 0 _0211_
rlabel metal1 15548 9418 15548 9418 0 _0212_
rlabel metal1 15272 8602 15272 8602 0 _0213_
rlabel metal2 13110 12580 13110 12580 0 _0214_
rlabel metal1 14582 9146 14582 9146 0 _0215_
rlabel metal1 14950 8602 14950 8602 0 _0216_
rlabel metal1 11132 13294 11132 13294 0 _0217_
rlabel metal1 10258 8058 10258 8058 0 _0218_
rlabel metal1 9752 8602 9752 8602 0 _0219_
rlabel metal1 10856 10778 10856 10778 0 _0220_
rlabel metal1 11776 13974 11776 13974 0 _0221_
rlabel metal2 9798 10438 9798 10438 0 _0222_
rlabel metal1 10350 12750 10350 12750 0 _0223_
rlabel metal1 14996 24106 14996 24106 0 _0224_
rlabel metal2 15778 26044 15778 26044 0 _0225_
rlabel metal2 11914 23460 11914 23460 0 _0226_
rlabel metal1 10764 23766 10764 23766 0 _0227_
rlabel metal1 16468 25806 16468 25806 0 _0228_
rlabel metal1 11270 24242 11270 24242 0 _0229_
rlabel metal1 4324 19142 4324 19142 0 _0230_
rlabel metal1 21850 20808 21850 20808 0 _0231_
rlabel metal1 19780 17034 19780 17034 0 _0232_
rlabel metal2 8142 19142 8142 19142 0 _0233_
rlabel metal1 21574 21658 21574 21658 0 _0234_
rlabel metal1 6808 22406 6808 22406 0 _0235_
rlabel metal1 13800 16422 13800 16422 0 _0236_
rlabel metal2 21298 18700 21298 18700 0 _0237_
rlabel metal1 20424 18258 20424 18258 0 _0238_
rlabel metal1 16100 14042 16100 14042 0 _0239_
rlabel metal2 21298 17340 21298 17340 0 _0240_
rlabel metal1 21022 18802 21022 18802 0 _0241_
rlabel metal1 25438 16762 25438 16762 0 _0242_
rlabel metal2 25070 16388 25070 16388 0 _0243_
rlabel metal1 25622 18870 25622 18870 0 _0244_
rlabel metal1 25484 18394 25484 18394 0 _0245_
rlabel metal1 24334 17034 24334 17034 0 _0246_
rlabel metal1 24702 18190 24702 18190 0 _0247_
rlabel metal1 23506 18632 23506 18632 0 _0248_
rlabel metal1 23644 17714 23644 17714 0 _0249_
rlabel metal1 23598 19244 23598 19244 0 _0250_
rlabel metal1 24104 19754 24104 19754 0 _0251_
rlabel metal1 22264 18190 22264 18190 0 _0252_
rlabel metal1 23552 16762 23552 16762 0 _0253_
rlabel metal1 16192 16966 16192 16966 0 _0254_
rlabel metal1 7820 16966 7820 16966 0 _0255_
rlabel metal1 13248 18802 13248 18802 0 _0256_
rlabel metal2 9982 19635 9982 19635 0 _0257_
rlabel metal1 15318 12954 15318 12954 0 _0258_
rlabel metal1 8878 13430 8878 13430 0 _0259_
rlabel metal1 19550 11322 19550 11322 0 _0260_
rlabel metal1 18676 10234 18676 10234 0 _0261_
rlabel metal1 17296 10234 17296 10234 0 _0262_
rlabel metal1 18814 12886 18814 12886 0 _0263_
rlabel metal1 17940 13294 17940 13294 0 _0264_
rlabel metal1 17434 10778 17434 10778 0 _0265_
rlabel metal1 15410 19210 15410 19210 0 _0266_
rlabel metal1 15456 21114 15456 21114 0 _0267_
rlabel metal1 13754 14382 13754 14382 0 _0268_
rlabel metal1 15456 11322 15456 11322 0 _0269_
rlabel metal1 14168 20570 14168 20570 0 _0270_
rlabel metal1 13846 10778 13846 10778 0 _0271_
rlabel metal1 15594 22712 15594 22712 0 _0272_
rlabel metal1 17342 23596 17342 23596 0 _0273_
rlabel metal1 14076 19958 14076 19958 0 _0274_
rlabel metal2 13846 22304 13846 22304 0 _0275_
rlabel metal1 16146 23732 16146 23732 0 _0276_
rlabel metal2 12098 19652 12098 19652 0 _0277_
rlabel metal2 13570 16728 13570 16728 0 _0278_
rlabel metal1 18906 14042 18906 14042 0 _0279_
rlabel metal1 18400 23154 18400 23154 0 _0280_
rlabel metal2 12650 18020 12650 18020 0 _0281_
rlabel metal1 18078 17204 18078 17204 0 _0282_
rlabel metal2 19274 22916 19274 22916 0 _0283_
rlabel metal2 13570 25840 13570 25840 0 _0284_
rlabel metal1 16192 25262 16192 25262 0 _0285_
rlabel metal1 17848 20434 17848 20434 0 _0286_
rlabel metal2 13386 25806 13386 25806 0 _0287_
rlabel metal2 15226 26044 15226 26044 0 _0288_
rlabel metal1 18952 25874 18952 25874 0 _0289_
rlabel metal1 18308 14246 18308 14246 0 _0290_
rlabel metal1 21620 12954 21620 12954 0 _0291_
rlabel metal1 20654 22508 20654 22508 0 _0292_
rlabel metal1 18078 15334 18078 15334 0 _0293_
rlabel metal1 19504 13838 19504 13838 0 _0294_
rlabel metal1 20562 14348 20562 14348 0 _0295_
rlabel metal1 20056 21862 20056 21862 0 _0296_
rlabel metal1 19458 20570 19458 20570 0 _0297_
rlabel metal1 17848 21862 17848 21862 0 _0298_
rlabel metal2 18998 21726 18998 21726 0 _0299_
rlabel metal2 18814 17918 18814 17918 0 _0300_
rlabel metal1 14030 21386 14030 21386 0 _0301_
rlabel metal1 21482 15130 21482 15130 0 _0302_
rlabel metal1 22954 16218 22954 16218 0 _0303_
rlabel metal1 21298 19244 21298 19244 0 _0304_
rlabel metal1 21344 14586 21344 14586 0 _0305_
rlabel metal1 18400 16082 18400 16082 0 _0306_
rlabel metal1 20240 19346 20240 19346 0 _0307_
rlabel metal1 16238 22984 16238 22984 0 _0308_
rlabel metal2 15318 20434 15318 20434 0 _0309_
rlabel metal1 17664 17850 17664 17850 0 _0310_
rlabel metal2 17434 22814 17434 22814 0 _0311_
rlabel metal1 12558 19720 12558 19720 0 _0312_
rlabel metal1 11914 18292 11914 18292 0 _0313_
rlabel metal1 18032 15062 18032 15062 0 _0314_
rlabel metal1 14076 16014 14076 16014 0 _0315_
rlabel metal1 16376 15062 16376 15062 0 _0316_
rlabel metal1 13202 15402 13202 15402 0 _0317_
rlabel metal1 23552 13498 23552 13498 0 _0318_
rlabel metal1 22586 12954 22586 12954 0 _0319_
rlabel metal1 23460 12954 23460 12954 0 _0320_
rlabel metal1 21298 12410 21298 12410 0 _0321_
rlabel metal1 4462 24242 4462 24242 0 _0322_
rlabel metal2 3266 25228 3266 25228 0 _0323_
rlabel metal1 4554 24786 4554 24786 0 _0324_
rlabel metal1 8786 23766 8786 23766 0 _0325_
rlabel metal1 16054 16150 16054 16150 0 _0326_
rlabel metal2 6670 24327 6670 24327 0 _0327_
rlabel metal1 7406 14586 7406 14586 0 _0328_
rlabel metal2 7866 24344 7866 24344 0 _0329_
rlabel metal2 6118 26860 6118 26860 0 _0330_
rlabel metal1 8970 25806 8970 25806 0 _0331_
rlabel metal1 7406 26860 7406 26860 0 _0332_
rlabel metal1 8648 26418 8648 26418 0 _0333_
rlabel metal2 24610 14824 24610 14824 0 _0334_
rlabel metal2 23782 16422 23782 16422 0 _0335_
rlabel metal1 24196 14926 24196 14926 0 _0336_
rlabel metal1 23460 15674 23460 15674 0 _0337_
rlabel metal1 7820 21658 7820 21658 0 _0338_
rlabel metal1 5474 20230 5474 20230 0 _0339_
rlabel metal1 9292 22066 9292 22066 0 _0340_
rlabel metal1 11776 20434 11776 20434 0 _0341_
rlabel metal1 15272 15402 15272 15402 0 _0342_
rlabel metal2 5566 24956 5566 24956 0 _0343_
rlabel metal1 5566 14450 5566 14450 0 _0344_
rlabel metal1 8004 24786 8004 24786 0 _0345_
rlabel metal2 23414 12002 23414 12002 0 _0346_
rlabel metal2 20470 12036 20470 12036 0 _0347_
rlabel metal1 21022 11866 21022 11866 0 _0348_
rlabel metal1 20148 13294 20148 13294 0 _0349_
rlabel metal1 14352 21930 14352 21930 0 _0350_
rlabel metal2 14122 15810 14122 15810 0 _0351_
rlabel metal1 10718 21998 10718 21998 0 _0352_
rlabel metal1 11960 24786 11960 24786 0 _0353_
rlabel metal2 14398 19414 14398 19414 0 _0354_
rlabel metal1 9108 6426 9108 6426 0 _0355_
rlabel metal1 14168 14246 14168 14246 0 _0356_
rlabel metal2 6394 5848 6394 5848 0 _0357_
rlabel metal2 13202 23256 13202 23256 0 _0358_
rlabel metal1 17572 17034 17572 17034 0 _0359_
rlabel metal1 14536 21590 14536 21590 0 _0360_
rlabel metal1 16560 16626 16560 16626 0 _0361_
rlabel metal1 17204 27506 17204 27506 0 _0362_
rlabel metal1 18722 25330 18722 25330 0 _0363_
rlabel metal1 17158 26962 17158 26962 0 _0364_
rlabel metal1 20746 26010 20746 26010 0 _0365_
rlabel metal1 23552 20570 23552 20570 0 _0366_
rlabel metal1 19274 14892 19274 14892 0 _0367_
rlabel metal2 21482 17068 21482 17068 0 _0368_
rlabel metal1 19918 14586 19918 14586 0 _0369_
rlabel metal2 6762 23902 6762 23902 0 _0370_
rlabel metal1 14168 24786 14168 24786 0 _0371_
rlabel metal2 7682 24446 7682 24446 0 _0372_
rlabel metal1 9292 25466 9292 25466 0 _0373_
rlabel metal2 18998 23902 18998 23902 0 _0374_
rlabel metal2 10258 20655 10258 20655 0 _0375_
rlabel metal1 17848 24378 17848 24378 0 _0376_
rlabel metal2 5290 22916 5290 22916 0 _0377_
rlabel metal1 7268 37230 7268 37230 0 ccff_head
rlabel metal1 4002 37094 4002 37094 0 ccff_tail
rlabel metal3 1142 27948 1142 27948 0 chanx_left_in[0]
rlabel metal2 38318 11679 38318 11679 0 chanx_left_in[10]
rlabel via2 38318 25245 38318 25245 0 chanx_left_in[11]
rlabel metal1 22724 37230 22724 37230 0 chanx_left_in[12]
rlabel metal2 10350 1588 10350 1588 0 chanx_left_in[13]
rlabel metal2 15502 1588 15502 1588 0 chanx_left_in[14]
rlabel metal2 32246 1588 32246 1588 0 chanx_left_in[15]
rlabel metal3 2338 1428 2338 1428 0 chanx_left_in[16]
rlabel metal2 38318 31569 38318 31569 0 chanx_left_in[17]
rlabel metal2 4554 1588 4554 1588 0 chanx_left_in[18]
rlabel metal2 34178 1588 34178 1588 0 chanx_left_in[1]
rlabel metal3 1142 32708 1142 32708 0 chanx_left_in[2]
rlabel metal1 33672 37230 33672 37230 0 chanx_left_in[3]
rlabel via2 38318 19805 38318 19805 0 chanx_left_in[4]
rlabel metal1 11776 37230 11776 37230 0 chanx_left_in[5]
rlabel metal3 1832 37468 1832 37468 0 chanx_left_in[6]
rlabel metal3 1142 25908 1142 25908 0 chanx_left_in[7]
rlabel metal2 38686 1554 38686 1554 0 chanx_left_in[8]
rlabel metal3 146 17748 146 17748 0 chanx_left_in[9]
rlabel metal2 38226 34833 38226 34833 0 chanx_left_out[0]
rlabel via2 38226 5525 38226 5525 0 chanx_left_out[10]
rlabel metal1 25944 37094 25944 37094 0 chanx_left_out[11]
rlabel metal2 1702 20859 1702 20859 0 chanx_left_out[12]
rlabel metal1 14950 37094 14950 37094 0 chanx_left_out[13]
rlabel metal1 16836 37094 16836 37094 0 chanx_left_out[14]
rlabel metal1 29486 37094 29486 37094 0 chanx_left_out[15]
rlabel metal3 1188 29308 1188 29308 0 chanx_left_out[16]
rlabel metal1 37720 36346 37720 36346 0 chanx_left_out[17]
rlabel via2 38226 33371 38226 33371 0 chanx_left_out[18]
rlabel metal2 38226 36941 38226 36941 0 chanx_left_out[1]
rlabel metal2 38226 8857 38226 8857 0 chanx_left_out[2]
rlabel metal1 24334 37094 24334 37094 0 chanx_left_out[3]
rlabel metal1 18216 37094 18216 37094 0 chanx_left_out[4]
rlabel metal3 1188 4828 1188 4828 0 chanx_left_out[5]
rlabel metal1 1702 37128 1702 37128 0 chanx_left_out[6]
rlabel metal2 9062 1520 9062 1520 0 chanx_left_out[7]
rlabel metal2 38226 28815 38226 28815 0 chanx_left_out[8]
rlabel metal2 37398 1520 37398 1520 0 chanx_left_out[9]
rlabel metal2 38318 15249 38318 15249 0 chany_top_in[0]
rlabel metal1 20838 37230 20838 37230 0 chany_top_in[10]
rlabel metal1 12972 37230 12972 37230 0 chany_top_in[11]
rlabel metal1 37122 3026 37122 3026 0 chany_top_in[12]
rlabel metal2 38318 30107 38318 30107 0 chany_top_in[13]
rlabel metal1 38180 35666 38180 35666 0 chany_top_in[14]
rlabel metal1 2162 3060 2162 3060 0 chany_top_in[15]
rlabel metal2 13570 1588 13570 1588 0 chany_top_in[16]
rlabel metal3 38786 6868 38786 6868 0 chany_top_in[17]
rlabel metal3 1142 22508 1142 22508 0 chany_top_in[18]
rlabel metal2 3542 2907 3542 2907 0 chany_top_in[1]
rlabel metal3 1142 30668 1142 30668 0 chany_top_in[2]
rlabel metal1 10488 37230 10488 37230 0 chany_top_in[3]
rlabel metal2 29026 1588 29026 1588 0 chany_top_in[4]
rlabel metal1 34960 37230 34960 37230 0 chany_top_in[5]
rlabel metal2 24518 1588 24518 1588 0 chany_top_in[6]
rlabel metal2 2622 1588 2622 1588 0 chany_top_in[7]
rlabel metal1 1610 23664 1610 23664 0 chany_top_in[8]
rlabel metal2 35466 1588 35466 1588 0 chany_top_in[9]
rlabel via2 38226 17051 38226 17051 0 chany_top_out[0]
rlabel metal2 38226 10353 38226 10353 0 chany_top_out[10]
rlabel metal2 27738 1520 27738 1520 0 chany_top_out[11]
rlabel metal3 1188 34068 1188 34068 0 chany_top_out[12]
rlabel metal2 38226 2465 38226 2465 0 chany_top_out[13]
rlabel metal1 5290 37094 5290 37094 0 chany_top_out[14]
rlabel via2 38226 13685 38226 13685 0 chany_top_out[15]
rlabel metal1 1656 16218 1656 16218 0 chany_top_out[16]
rlabel metal2 30958 1520 30958 1520 0 chany_top_out[17]
rlabel metal2 38226 26673 38226 26673 0 chany_top_out[18]
rlabel metal2 18722 1520 18722 1520 0 chany_top_out[1]
rlabel metal3 1188 24548 1188 24548 0 chany_top_out[2]
rlabel metal2 20010 1520 20010 1520 0 chany_top_out[3]
rlabel metal2 46 1520 46 1520 0 chany_top_out[4]
rlabel metal2 23230 1520 23230 1520 0 chany_top_out[5]
rlabel metal1 1656 7514 1656 7514 0 chany_top_out[6]
rlabel metal1 19504 37094 19504 37094 0 chany_top_out[7]
rlabel metal2 4094 13073 4094 13073 0 chany_top_out[8]
rlabel metal1 1196 36890 1196 36890 0 chany_top_out[9]
rlabel metal1 5152 20774 5152 20774 0 clknet_0_prog_clk
rlabel metal2 2162 9452 2162 9452 0 clknet_3_0__leaf_prog_clk
rlabel metal1 1702 10710 1702 10710 0 clknet_3_1__leaf_prog_clk
rlabel metal1 7912 9010 7912 9010 0 clknet_3_2__leaf_prog_clk
rlabel metal1 7544 14450 7544 14450 0 clknet_3_3__leaf_prog_clk
rlabel metal1 1702 16694 1702 16694 0 clknet_3_4__leaf_prog_clk
rlabel metal1 2208 21114 2208 21114 0 clknet_3_5__leaf_prog_clk
rlabel metal1 10626 18292 10626 18292 0 clknet_3_6__leaf_prog_clk
rlabel metal2 9154 20400 9154 20400 0 clknet_3_7__leaf_prog_clk
rlabel metal2 5842 1588 5842 1588 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 1334 1860 1334 1860 0 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 36846 37230 36846 37230 0 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 27232 37230 27232 37230 0 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 16790 1588 16790 1588 0 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 36938 36788 36938 36788 0 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
rlabel via2 38318 3485 38318 3485 0 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal1 1610 5712 1610 5712 0 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 38318 21913 38318 21913 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 7774 1588 7774 1588 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 10258 17408 10258 17408 0 mem_left_track_1.DFFR_0_.D
rlabel metal2 22034 18462 22034 18462 0 mem_left_track_1.DFFR_0_.Q
rlabel metal2 21114 19329 21114 19329 0 mem_left_track_1.DFFR_1_.Q
rlabel metal1 3312 21590 3312 21590 0 mem_left_track_11.DFFR_0_.D
rlabel metal1 1886 21454 1886 21454 0 mem_left_track_11.DFFR_0_.Q
rlabel metal1 4002 17578 4002 17578 0 mem_left_track_11.DFFR_1_.Q
rlabel metal2 17342 19975 17342 19975 0 mem_left_track_13.DFFR_0_.Q
rlabel via2 12650 26979 12650 26979 0 mem_left_track_13.DFFR_1_.Q
rlabel metal1 21298 18734 21298 18734 0 mem_left_track_15.DFFR_0_.Q
rlabel metal2 1702 11424 1702 11424 0 mem_left_track_15.DFFR_1_.Q
rlabel metal1 1978 19720 1978 19720 0 mem_left_track_17.DFFR_0_.Q
rlabel metal1 20010 21488 20010 21488 0 mem_left_track_17.DFFR_1_.Q
rlabel metal1 16928 16082 16928 16082 0 mem_left_track_19.DFFR_0_.Q
rlabel metal1 21482 14416 21482 14416 0 mem_left_track_19.DFFR_1_.Q
rlabel metal1 19642 11662 19642 11662 0 mem_left_track_21.DFFR_0_.Q
rlabel metal1 21160 11730 21160 11730 0 mem_left_track_21.DFFR_1_.Q
rlabel metal1 11408 13498 11408 13498 0 mem_left_track_23.DFFR_0_.Q
rlabel metal2 13478 17306 13478 17306 0 mem_left_track_23.DFFR_1_.Q
rlabel metal2 6762 6018 6762 6018 0 mem_left_track_25.DFFR_0_.Q
rlabel metal1 13570 9588 13570 9588 0 mem_left_track_25.DFFR_1_.Q
rlabel metal2 10902 15266 10902 15266 0 mem_left_track_27.DFFR_0_.Q
rlabel metal2 13202 25670 13202 25670 0 mem_left_track_27.DFFR_1_.Q
rlabel metal1 20056 25874 20056 25874 0 mem_left_track_29.DFFR_0_.Q
rlabel metal1 16008 28526 16008 28526 0 mem_left_track_29.DFFR_1_.Q
rlabel metal1 14766 12886 14766 12886 0 mem_left_track_3.DFFR_0_.Q
rlabel metal1 14490 15912 14490 15912 0 mem_left_track_3.DFFR_1_.Q
rlabel metal2 19458 14586 19458 14586 0 mem_left_track_31.DFFR_0_.Q
rlabel metal2 21574 17714 21574 17714 0 mem_left_track_31.DFFR_1_.Q
rlabel metal1 10488 19754 10488 19754 0 mem_left_track_33.DFFR_0_.Q
rlabel metal2 9246 20740 9246 20740 0 mem_left_track_33.DFFR_1_.Q
rlabel metal1 8142 21318 8142 21318 0 mem_left_track_35.DFFR_0_.Q
rlabel metal1 10304 20774 10304 20774 0 mem_left_track_35.DFFR_1_.Q
rlabel metal2 14858 17986 14858 17986 0 mem_left_track_37.DFFR_0_.Q
rlabel metal1 1748 7786 1748 7786 0 mem_left_track_5.DFFR_0_.Q
rlabel via2 19550 10659 19550 10659 0 mem_left_track_5.DFFR_1_.Q
rlabel metal1 15410 21998 15410 21998 0 mem_left_track_7.DFFR_0_.Q
rlabel metal1 13064 20434 13064 20434 0 mem_left_track_7.DFFR_1_.Q
rlabel metal1 6486 18870 6486 18870 0 mem_left_track_9.DFFR_0_.Q
rlabel metal1 7590 19856 7590 19856 0 mem_top_track_0.DFFR_0_.Q
rlabel metal2 13018 14450 13018 14450 0 mem_top_track_0.DFFR_1_.Q
rlabel metal1 5980 12886 5980 12886 0 mem_top_track_10.DFFR_0_.D
rlabel metal1 14674 8500 14674 8500 0 mem_top_track_10.DFFR_0_.Q
rlabel metal2 1702 9248 1702 9248 0 mem_top_track_10.DFFR_1_.Q
rlabel metal1 5290 7922 5290 7922 0 mem_top_track_12.DFFR_0_.Q
rlabel metal1 7130 8058 7130 8058 0 mem_top_track_12.DFFR_1_.Q
rlabel metal1 15502 25942 15502 25942 0 mem_top_track_14.DFFR_0_.Q
rlabel metal1 1564 21862 1564 21862 0 mem_top_track_14.DFFR_1_.Q
rlabel metal1 21436 20434 21436 20434 0 mem_top_track_16.DFFR_0_.Q
rlabel metal1 3266 19346 3266 19346 0 mem_top_track_16.DFFR_1_.Q
rlabel metal2 2162 18445 2162 18445 0 mem_top_track_18.DFFR_0_.Q
rlabel metal2 9338 15113 9338 15113 0 mem_top_track_18.DFFR_1_.Q
rlabel metal1 1794 12070 1794 12070 0 mem_top_track_2.DFFR_0_.Q
rlabel metal1 13754 8976 13754 8976 0 mem_top_track_2.DFFR_1_.Q
rlabel metal1 10580 13770 10580 13770 0 mem_top_track_20.DFFR_0_.Q
rlabel metal1 16790 11152 16790 11152 0 mem_top_track_20.DFFR_1_.Q
rlabel metal1 21666 12172 21666 12172 0 mem_top_track_22.DFFR_0_.Q
rlabel metal2 22770 10846 22770 10846 0 mem_top_track_22.DFFR_1_.Q
rlabel metal2 6348 18700 6348 18700 0 mem_top_track_24.DFFR_0_.Q
rlabel metal1 4600 21930 4600 21930 0 mem_top_track_24.DFFR_1_.Q
rlabel metal1 7038 17034 7038 17034 0 mem_top_track_26.DFFR_0_.Q
rlabel metal1 5060 17170 5060 17170 0 mem_top_track_26.DFFR_1_.Q
rlabel metal2 9292 21556 9292 21556 0 mem_top_track_28.DFFR_0_.Q
rlabel metal1 7544 20774 7544 20774 0 mem_top_track_28.DFFR_1_.Q
rlabel metal1 24610 16116 24610 16116 0 mem_top_track_30.DFFR_0_.Q
rlabel metal2 1978 10829 1978 10829 0 mem_top_track_30.DFFR_1_.Q
rlabel metal1 4232 19822 4232 19822 0 mem_top_track_32.DFFR_0_.Q
rlabel metal1 7038 18734 7038 18734 0 mem_top_track_32.DFFR_1_.Q
rlabel metal1 7636 25262 7636 25262 0 mem_top_track_34.DFFR_0_.Q
rlabel metal1 13662 11764 13662 11764 0 mem_top_track_34.DFFR_1_.Q
rlabel metal1 1886 15368 1886 15368 0 mem_top_track_36.DFFR_0_.Q
rlabel metal1 16054 25874 16054 25874 0 mem_top_track_4.DFFR_0_.Q
rlabel metal1 13570 26316 13570 26316 0 mem_top_track_4.DFFR_1_.Q
rlabel metal2 8464 19788 8464 19788 0 mem_top_track_6.DFFR_0_.Q
rlabel metal1 6716 12818 6716 12818 0 mem_top_track_6.DFFR_1_.Q
rlabel metal1 1702 19380 1702 19380 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 34914 16558 34914 16558 0 mux_left_track_1.INVTX1_0_.out
rlabel metal2 32154 20094 32154 20094 0 mux_left_track_1.INVTX1_1_.out
rlabel metal3 13455 18020 13455 18020 0 mux_left_track_1.INVTX1_2_.out
rlabel metal2 23138 18598 23138 18598 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23046 18394 23046 18394 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 26818 25874 26818 25874 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 31786 26010 31786 26010 0 mux_left_track_1.out
rlabel metal2 33258 24687 33258 24687 0 mux_left_track_11.INVTX1_0_.out
rlabel metal1 21114 31790 21114 31790 0 mux_left_track_11.INVTX1_1_.out
rlabel via1 17894 17187 17894 17187 0 mux_left_track_11.INVTX1_2_.out
rlabel metal2 18906 22576 18906 22576 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18078 17034 18078 17034 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 12926 17578 12926 17578 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 11270 9894 11270 9894 0 mux_left_track_11.out
rlabel metal2 34086 28288 34086 28288 0 mux_left_track_13.INVTX1_0_.out
rlabel metal2 30498 26010 30498 26010 0 mux_left_track_13.INVTX1_2_.out
rlabel metal1 18492 20570 18492 20570 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14536 25398 14536 25398 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 13018 27778 13018 27778 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6716 35054 6716 35054 0 mux_left_track_13.out
rlabel metal1 23506 6766 23506 6766 0 mux_left_track_15.INVTX1_0_.out
rlabel metal1 19320 13906 19320 13906 0 mux_left_track_15.INVTX1_2_.out
rlabel metal1 20424 14586 20424 14586 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 20010 14416 20010 14416 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17480 14314 17480 14314 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 9614 3468 9614 3468 0 mux_left_track_15.out
rlabel metal1 15548 34510 15548 34510 0 mux_left_track_17.INVTX1_0_.out
rlabel metal2 14582 19533 14582 19533 0 mux_left_track_17.INVTX1_2_.out
rlabel metal1 17618 22066 17618 22066 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19550 21012 19550 21012 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 35650 23324 35650 23324 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 36110 25908 36110 25908 0 mux_left_track_17.out
rlabel metal1 20516 34510 20516 34510 0 mux_left_track_19.INVTX1_0_.out
rlabel metal1 21022 19346 21022 19346 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20424 16150 20424 16150 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 21482 15742 21482 15742 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30222 11526 30222 11526 0 mux_left_track_19.out
rlabel metal1 23598 6664 23598 6664 0 mux_left_track_21.INVTX1_0_.out
rlabel metal1 20976 12750 20976 12750 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23322 12342 23322 12342 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 34224 7854 34224 7854 0 mux_left_track_21.out
rlabel metal1 11730 24684 11730 24684 0 mux_left_track_23.INVTX1_0_.out
rlabel via2 14950 17629 14950 17629 0 mux_left_track_23.INVTX1_1_.out
rlabel metal1 11592 22066 11592 22066 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 14674 22015 14674 22015 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 21988 34578 21988 34578 0 mux_left_track_23.out
rlabel metal1 6302 5780 6302 5780 0 mux_left_track_25.INVTX1_0_.out
rlabel metal1 13018 14382 13018 14382 0 mux_left_track_25.INVTX1_1_.out
rlabel metal1 9660 6834 9660 6834 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16422 19703 16422 19703 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 7958 25942 7958 25942 0 mux_left_track_25.out
rlabel metal2 21620 13838 21620 13838 0 mux_left_track_27.INVTX1_0_.out
rlabel metal2 29210 25024 29210 25024 0 mux_left_track_27.INVTX1_1_.out
rlabel metal1 17940 16490 17940 16490 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13892 33490 13892 33490 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14996 33626 14996 33626 0 mux_left_track_27.out
rlabel metal1 24518 33830 24518 33830 0 mux_left_track_29.INVTX1_0_.out
rlabel metal2 18170 26724 18170 26724 0 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16698 29444 16698 29444 0 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17020 31450 17020 31450 0 mux_left_track_29.out
rlabel metal1 11868 19890 11868 19890 0 mux_left_track_3.INVTX1_0_.out
rlabel metal1 14766 19890 14766 19890 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16606 18530 16606 18530 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 17250 19278 17250 19278 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 31556 27098 31556 27098 0 mux_left_track_3.out
rlabel metal1 24518 7514 24518 7514 0 mux_left_track_31.INVTX1_0_.out
rlabel metal1 20332 15674 20332 15674 0 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24012 29614 24012 29614 0 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 24702 32198 24702 32198 0 mux_left_track_31.out
rlabel metal1 10350 33830 10350 33830 0 mux_left_track_33.INVTX1_0_.out
rlabel metal1 13294 24684 13294 24684 0 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 7084 23766 7084 23766 0 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 3818 26486 3818 26486 0 mux_left_track_33.out
rlabel via1 9246 23018 9246 23018 0 mux_left_track_35.INVTX1_0_.out
rlabel via1 18906 22073 18906 22073 0 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 37582 30770 37582 30770 0 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 37398 36346 37398 36346 0 mux_left_track_35.out
rlabel metal1 10166 14926 10166 14926 0 mux_left_track_37.INVTX1_0_.out
rlabel metal2 17342 18836 17342 18836 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16008 20570 16008 20570 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 33350 25466 33350 25466 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 33396 28730 33396 28730 0 mux_left_track_37.out
rlabel metal2 17664 10948 17664 10948 0 mux_left_track_5.INVTX1_0_.out
rlabel metal1 17802 12682 17802 12682 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18906 12750 18906 12750 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 29072 10642 29072 10642 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 32522 10030 32522 10030 0 mux_left_track_5.out
rlabel metal1 14398 13838 14398 13838 0 mux_left_track_7.INVTX1_0_.out
rlabel metal1 14490 14518 14490 14518 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16790 21318 16790 21318 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17526 20808 17526 20808 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 20654 34646 20654 34646 0 mux_left_track_7.out
rlabel metal3 11983 19380 11983 19380 0 mux_left_track_9.INVTX1_0_.out
rlabel metal1 15456 20774 15456 20774 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16422 23494 16422 23494 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16560 22474 16560 22474 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 17342 29818 17342 29818 0 mux_left_track_9.out
rlabel metal1 20056 18734 20056 18734 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 17756 16014 17756 16014 0 mux_top_track_0.INVTX1_1_.out
rlabel metal1 10304 23086 10304 23086 0 mux_top_track_0.INVTX1_2_.out
rlabel metal1 18078 17510 18078 17510 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14996 20774 14996 20774 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 18538 17986 18538 17986 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 33810 17340 33810 17340 0 mux_top_track_0.out
rlabel metal1 13984 17102 13984 17102 0 mux_top_track_10.INVTX1_0_.out
rlabel metal1 21988 16014 21988 16014 0 mux_top_track_10.INVTX1_1_.out
rlabel metal1 15686 5882 15686 5882 0 mux_top_track_10.INVTX1_2_.out
rlabel metal1 13662 14790 13662 14790 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 15594 11866 15594 11866 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17204 12886 17204 12886 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 20194 7004 20194 7004 0 mux_top_track_10.out
rlabel metal1 11546 12274 11546 12274 0 mux_top_track_12.INVTX1_1_.out
rlabel metal2 9982 8772 9982 8772 0 mux_top_track_12.INVTX1_2_.out
rlabel metal1 11684 13838 11684 13838 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 10764 11526 10764 11526 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 12052 13838 12052 13838 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 4462 5236 4462 5236 0 mux_top_track_12.out
rlabel metal1 10764 19346 10764 19346 0 mux_top_track_14.INVTX1_1_.out
rlabel metal1 18768 33286 18768 33286 0 mux_top_track_14.INVTX1_2_.out
rlabel metal2 12006 23834 12006 23834 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16560 24718 16560 24718 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 14674 26962 14674 26962 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 16698 35054 16698 35054 0 mux_top_track_14.out
rlabel metal1 20194 18156 20194 18156 0 mux_top_track_16.INVTX1_1_.out
rlabel metal2 21942 22780 21942 22780 0 mux_top_track_16.INVTX1_2_.out
rlabel metal2 11086 18972 11086 18972 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20010 21930 20010 21930 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 12742 19142 12742 19142 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 14306 11118 14306 11118 0 mux_top_track_16.out
rlabel metal2 21758 15776 21758 15776 0 mux_top_track_18.INVTX1_2_.out
rlabel metal2 19458 19142 19458 19142 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20792 18054 20792 18054 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 15594 19040 15594 19040 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 9522 34578 9522 34578 0 mux_top_track_18.out
rlabel metal2 27278 27098 27278 27098 0 mux_top_track_2.INVTX1_1_.out
rlabel metal1 9614 6222 9614 6222 0 mux_top_track_2.INVTX1_2_.out
rlabel metal2 15134 14688 15134 14688 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 12926 12954 12926 12954 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15778 13974 15778 13974 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 16882 4590 16882 4590 0 mux_top_track_2.out
rlabel metal1 13202 11254 13202 11254 0 mux_top_track_20.INVTX1_1_.out
rlabel metal2 14306 15776 14306 15776 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18630 14858 18630 14858 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 32936 11730 32936 11730 0 mux_top_track_20.out
rlabel metal1 28520 7242 28520 7242 0 mux_top_track_22.INVTX1_1_.out
rlabel metal2 22402 13702 22402 13702 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24104 8942 24104 8942 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25392 8806 25392 8806 0 mux_top_track_22.out
rlabel metal2 25438 26894 25438 26894 0 mux_top_track_24.INVTX1_0_.out
rlabel metal2 3082 24990 3082 24990 0 mux_top_track_24.INVTX1_1_.out
rlabel metal1 4876 24718 4876 24718 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 4922 26656 4922 26656 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 4094 29716 4094 29716 0 mux_top_track_24.out
rlabel metal1 7222 30022 7222 30022 0 mux_top_track_26.INVTX1_0_.out
rlabel metal1 5796 32198 5796 32198 0 mux_top_track_26.INVTX1_1_.out
rlabel metal2 9936 20740 9936 20740 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 36846 8738 36846 8738 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 37490 5372 37490 5372 0 mux_top_track_26.out
rlabel metal1 9108 33830 9108 33830 0 mux_top_track_28.INVTX1_1_.out
rlabel metal1 7636 26214 7636 26214 0 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 6302 28628 6302 28628 0 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 6072 30906 6072 30906 0 mux_top_track_28.out
rlabel metal2 34270 17374 34270 17374 0 mux_top_track_30.INVTX1_1_.out
rlabel metal2 22678 16320 22678 16320 0 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23138 14892 23138 14892 0 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 29302 14348 29302 14348 0 mux_top_track_30.out
rlabel metal1 20746 33354 20746 33354 0 mux_top_track_32.INVTX1_1_.out
rlabel metal2 12374 20672 12374 20672 0 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 12558 24820 12558 24820 0 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 12742 25738 12742 25738 0 mux_top_track_32.out
rlabel metal2 5382 26622 5382 26622 0 mux_top_track_34.INVTX1_1_.out
rlabel metal1 8786 24582 8786 24582 0 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24196 10030 24196 10030 0 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25162 9962 25162 9962 0 mux_top_track_34.out
rlabel metal1 27186 6630 27186 6630 0 mux_top_track_36.INVTX1_2_.out
rlabel metal2 24702 18972 24702 18972 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24380 16762 24380 16762 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 25346 20162 25346 20162 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 33166 22916 33166 22916 0 mux_top_track_36.out
rlabel metal2 20746 26316 20746 26316 0 mux_top_track_4.INVTX1_2_.out
rlabel metal1 17986 24038 17986 24038 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18952 24106 18952 24106 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 14582 24582 14582 24582 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 4738 25296 4738 25296 0 mux_top_track_4.out
rlabel metal1 9706 6630 9706 6630 0 mux_top_track_6.INVTX1_2_.out
rlabel metal1 11132 22678 11132 22678 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 11730 14450 11730 14450 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 14582 14416 14582 14416 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 16882 6766 16882 6766 0 mux_top_track_6.out
rlabel metal2 16698 9146 16698 9146 0 mux_top_track_8.INVTX1_2_.out
rlabel metal1 13386 17000 13386 17000 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16790 14246 16790 14246 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 11040 14858 11040 14858 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 5244 4590 5244 4590 0 mux_top_track_8.out
rlabel via3 7245 36516 7245 36516 0 net1
rlabel metal2 33810 29988 33810 29988 0 net10
rlabel metal1 12604 20502 12604 20502 0 net100
rlabel metal1 12512 9690 12512 9690 0 net101
rlabel metal2 21114 24480 21114 24480 0 net102
rlabel metal1 6118 13362 6118 13362 0 net103
rlabel metal1 15916 10778 15916 10778 0 net104
rlabel metal2 15042 10336 15042 10336 0 net105
rlabel metal2 10350 9962 10350 9962 0 net106
rlabel metal1 15548 24786 15548 24786 0 net107
rlabel metal2 21942 21216 21942 21216 0 net108
rlabel metal2 22678 18428 22678 18428 0 net109
rlabel metal1 6440 6222 6440 6222 0 net11
rlabel metal1 25392 16626 25392 16626 0 net110
rlabel metal2 22678 17476 22678 17476 0 net111
rlabel metal2 16882 16116 16882 16116 0 net112
rlabel metal2 18906 11492 18906 11492 0 net113
rlabel metal2 16882 21590 16882 21590 0 net114
rlabel metal1 17526 23766 17526 23766 0 net115
rlabel metal2 17986 15572 17986 15572 0 net116
rlabel metal1 16192 25330 16192 25330 0 net117
rlabel metal1 21252 13362 21252 13362 0 net118
rlabel metal1 20148 20570 20148 20570 0 net119
rlabel metal1 32752 2550 32752 2550 0 net12
rlabel metal1 18952 15538 18952 15538 0 net120
rlabel metal1 15134 20434 15134 20434 0 net121
rlabel metal1 17940 11866 17940 11866 0 net122
rlabel metal1 23368 13838 23368 13838 0 net123
rlabel metal1 3404 24242 3404 24242 0 net124
rlabel metal1 16284 11866 16284 11866 0 net125
rlabel metal2 5934 26860 5934 26860 0 net126
rlabel metal2 23322 14654 23322 14654 0 net127
rlabel metal1 11546 23154 11546 23154 0 net128
rlabel metal2 15088 15402 15088 15402 0 net129
rlabel metal1 3220 32742 3220 32742 0 net13
rlabel metal1 22678 12138 22678 12138 0 net130
rlabel metal2 14398 23596 14398 23596 0 net131
rlabel metal1 15180 18394 15180 18394 0 net132
rlabel metal2 13110 24140 13110 24140 0 net133
rlabel metal1 17618 27370 17618 27370 0 net134
rlabel metal2 22862 20706 22862 20706 0 net135
rlabel metal1 6440 22678 6440 22678 0 net136
rlabel metal1 19182 23630 19182 23630 0 net137
rlabel metal1 31510 37162 31510 37162 0 net14
rlabel metal2 35558 18972 35558 18972 0 net15
rlabel metal1 11316 37094 11316 37094 0 net16
rlabel metal1 4232 32402 4232 32402 0 net17
rlabel metal2 1886 25466 1886 25466 0 net18
rlabel metal1 35558 2618 35558 2618 0 net19
rlabel metal1 2852 29002 2852 29002 0 net2
rlabel via3 1909 26316 1909 26316 0 net20
rlabel metal2 38134 16150 38134 16150 0 net21
rlabel metal2 20746 35836 20746 35836 0 net22
rlabel metal1 13984 37094 13984 37094 0 net23
rlabel metal2 35650 4964 35650 4964 0 net24
rlabel metal2 35466 29274 35466 29274 0 net25
rlabel metal2 33258 35020 33258 35020 0 net26
rlabel metal2 6670 5100 6670 5100 0 net27
rlabel metal1 14398 2618 14398 2618 0 net28
rlabel metal2 38134 8534 38134 8534 0 net29
rlabel metal1 37536 11866 37536 11866 0 net3
rlabel metal1 1840 22746 1840 22746 0 net30
rlabel metal1 5336 2890 5336 2890 0 net31
rlabel metal2 9154 29138 9154 29138 0 net32
rlabel metal1 10396 37094 10396 37094 0 net33
rlabel metal1 27232 7378 27232 7378 0 net34
rlabel metal1 32614 36890 32614 36890 0 net35
rlabel metal1 24012 2618 24012 2618 0 net36
rlabel metal1 3082 2618 3082 2618 0 net37
rlabel metal1 1840 23834 1840 23834 0 net38
rlabel metal1 34316 2278 34316 2278 0 net39
rlabel metal2 34822 24412 34822 24412 0 net4
rlabel metal1 7038 2618 7038 2618 0 net40
rlabel metal1 4186 3162 4186 3162 0 net41
rlabel metal1 36340 37094 36340 37094 0 net42
rlabel metal1 25254 31790 25254 31790 0 net43
rlabel metal1 17020 2618 17020 2618 0 net44
rlabel metal2 36754 33082 36754 33082 0 net45
rlabel metal1 34454 3706 34454 3706 0 net46
rlabel metal1 2277 5542 2277 5542 0 net47
rlabel metal2 32246 21386 32246 21386 0 net48
rlabel metal1 8970 2618 8970 2618 0 net49
rlabel metal1 21344 37162 21344 37162 0 net5
rlabel metal2 12650 3536 12650 3536 0 net50
rlabel metal2 34546 22508 34546 22508 0 net51
rlabel metal1 21252 2618 21252 2618 0 net52
rlabel metal1 29854 30158 29854 30158 0 net53
rlabel metal1 28014 29614 28014 29614 0 net54
rlabel metal1 4784 37162 4784 37162 0 net55
rlabel metal1 8740 37094 8740 37094 0 net56
rlabel metal2 25438 6324 25438 6324 0 net57
rlabel metal2 11730 7310 11730 7310 0 net58
rlabel metal1 4232 36006 4232 36006 0 net59
rlabel metal1 10258 2618 10258 2618 0 net6
rlabel metal1 37007 18598 37007 18598 0 net60
rlabel metal3 4761 36652 4761 36652 0 net61
rlabel metal1 35236 30906 35236 30906 0 net62
rlabel metal2 38042 6698 38042 6698 0 net63
rlabel metal1 25346 37230 25346 37230 0 net64
rlabel metal1 2392 20434 2392 20434 0 net65
rlabel metal1 15364 34714 15364 34714 0 net66
rlabel metal2 16882 36516 16882 36516 0 net67
rlabel metal1 28612 37230 28612 37230 0 net68
rlabel metal1 2622 29580 2622 29580 0 net69
rlabel metal1 15548 2618 15548 2618 0 net7
rlabel metal1 37812 36142 37812 36142 0 net70
rlabel metal2 33534 31790 33534 31790 0 net71
rlabel metal1 38042 37196 38042 37196 0 net72
rlabel metal2 38042 9418 38042 9418 0 net73
rlabel metal1 23782 37230 23782 37230 0 net74
rlabel metal1 17940 35258 17940 35258 0 net75
rlabel metal1 1886 5100 1886 5100 0 net76
rlabel metal1 2944 36890 2944 36890 0 net77
rlabel metal2 9430 2618 9430 2618 0 net78
rlabel metal1 37168 26554 37168 26554 0 net79
rlabel metal1 31326 2618 31326 2618 0 net8
rlabel metal1 37490 2448 37490 2448 0 net80
rlabel metal1 36961 17170 36961 17170 0 net81
rlabel metal2 35374 11084 35374 11084 0 net82
rlabel metal2 27830 3740 27830 3740 0 net83
rlabel metal1 2944 34578 2944 34578 0 net84
rlabel metal2 38042 4012 38042 4012 0 net85
rlabel metal1 5658 35802 5658 35802 0 net86
rlabel metal1 36961 13906 36961 13906 0 net87
rlabel metal1 1932 16082 1932 16082 0 net88
rlabel metal1 30544 2414 30544 2414 0 net89
rlabel metal1 4462 3706 4462 3706 0 net9
rlabel metal2 35374 25670 35374 25670 0 net90
rlabel metal1 17894 4454 17894 4454 0 net91
rlabel metal1 1886 24752 1886 24752 0 net92
rlabel metal1 18584 4998 18584 4998 0 net93
rlabel metal1 1886 2448 1886 2448 0 net94
rlabel metal2 23322 3706 23322 3706 0 net95
rlabel metal1 1886 7276 1886 7276 0 net96
rlabel metal1 18860 37230 18860 37230 0 net97
rlabel metal1 4876 13294 4876 13294 0 net98
rlabel metal1 2990 36754 2990 36754 0 net99
rlabel metal2 12282 1588 12282 1588 0 pReset
rlabel metal2 3726 14739 3726 14739 0 prog_clk
rlabel metal2 38318 23443 38318 23443 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 21298 1588 21298 1588 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal1 32154 37230 32154 37230 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 30544 37230 30544 37230 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 2162 37230 2162 37230 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 8878 37230 8878 37230 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 26450 1588 26450 1588 0 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 2116 6426 2116 6426 0 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal3 1142 36108 1142 36108 0 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 38318 18581 38318 18581 0 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
