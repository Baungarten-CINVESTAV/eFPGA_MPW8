VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2808.930 BY 2948.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.940 0.000 1243.220 3.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.980 2945.000 1024.260 2948.000 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.140 0.000 2241.420 3.000 ;
    END
  END clk
  PIN gfpga_pad_GPIO_PAD_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.080 0.000 2489.360 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[0]
  PIN gfpga_pad_GPIO_PAD_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.760 0.000 1826.040 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[10]
  PIN gfpga_pad_GPIO_PAD_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.920 2945.000 1272.200 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[11]
  PIN gfpga_pad_GPIO_PAD_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 97.640 2808.930 98.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[12]
  PIN gfpga_pad_GPIO_PAD_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2552.440 2808.930 2553.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[13]
  PIN gfpga_pad_GPIO_PAD_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2769.220 2945.000 2769.500 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[14]
  PIN gfpga_pad_GPIO_PAD_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.300 2945.000 1687.580 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[15]
  PIN gfpga_pad_GPIO_PAD_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.060 0.000 747.340 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[16]
  PIN gfpga_pad_GPIO_PAD_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 611.040 3.930 611.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[17]
  PIN gfpga_pad_GPIO_PAD_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 699.440 3.930 700.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[18]
  PIN gfpga_pad_GPIO_PAD_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 522.640 3.930 523.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[19]
  PIN gfpga_pad_GPIO_PAD_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.360 2945.000 1439.640 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[1]
  PIN gfpga_pad_GPIO_PAD_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.940 2945.000 277.220 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[20]
  PIN gfpga_pad_GPIO_PAD_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2290.640 2808.930 2291.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[21]
  PIN gfpga_pad_GPIO_PAD_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2103.640 3.930 2104.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[22]
  PIN gfpga_pad_GPIO_PAD_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2379.040 2808.930 2379.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[23]
  PIN gfpga_pad_GPIO_PAD_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.560 0.000 827.840 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[24]
  PIN gfpga_pad_GPIO_PAD_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.780 2945.000 2602.060 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[25]
  PIN gfpga_pad_GPIO_PAD_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.740 2945.000 1855.020 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[26]
  PIN gfpga_pad_GPIO_PAD_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.660 2945.000 360.940 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[27]
  PIN gfpga_pad_GPIO_PAD_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.640 2945.000 1355.920 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[28]
  PIN gfpga_pad_GPIO_PAD_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2365.440 3.930 2366.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[29]
  PIN gfpga_pad_GPIO_PAD_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1151.640 2808.930 1152.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[2]
  PIN gfpga_pad_GPIO_PAD_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1665.040 3.930 1665.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[30]
  PIN gfpga_pad_GPIO_PAD_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 9.240 2808.930 9.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[31]
  PIN gfpga_pad_GPIO_PAD_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.500 2945.000 109.780 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[32]
  PIN gfpga_pad_GPIO_PAD_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.280 0.000 911.560 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[33]
  PIN gfpga_pad_GPIO_PAD_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1240.040 2808.930 1240.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[34]
  PIN gfpga_pad_GPIO_PAD_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.440 0.000 1162.720 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[35]
  PIN gfpga_pad_GPIO_PAD_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1226.440 3.930 1227.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[36]
  PIN gfpga_pad_GPIO_PAD_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.160 2945.000 441.440 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[37]
  PIN gfpga_pad_GPIO_PAD_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.080 2945.000 1523.360 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[38]
  PIN gfpga_pad_GPIO_PAD_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.840 2945.000 2354.120 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[39]
  PIN gfpga_pad_GPIO_PAD_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1763.640 2808.930 1764.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[3]
  PIN gfpga_pad_GPIO_PAD_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1852.040 2808.930 1852.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[40]
  PIN gfpga_pad_GPIO_PAD_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.600 2945.000 608.880 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[41]
  PIN gfpga_pad_GPIO_PAD_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.120 2945.000 2270.400 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[42]
  PIN gfpga_pad_GPIO_PAD_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.040 0.000 1742.320 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[43]
  PIN gfpga_pad_GPIO_PAD_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.380 0.000 1410.660 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[44]
  PIN gfpga_pad_GPIO_PAD_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2028.840 2808.930 2029.440 ;
    END
  END gfpga_pad_GPIO_PAD_in[45]
  PIN gfpga_pad_GPIO_PAD_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2740.240 0.000 2740.520 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[46]
  PIN gfpga_pad_GPIO_PAD_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.360 0.000 2405.640 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[47]
  PIN gfpga_pad_GPIO_PAD_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1325.040 2808.930 1325.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[48]
  PIN gfpga_pad_GPIO_PAD_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.340 2945.000 2434.620 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[49]
  PIN gfpga_pad_GPIO_PAD_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.100 0.000 1494.380 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[4]
  PIN gfpga_pad_GPIO_PAD_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 886.440 2808.930 887.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[50]
  PIN gfpga_pad_GPIO_PAD_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.340 0.000 663.620 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[51]
  PIN gfpga_pad_GPIO_PAD_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.520 0.000 80.800 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[52]
  PIN gfpga_pad_GPIO_PAD_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 801.440 2808.930 802.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[53]
  PIN gfpga_pad_GPIO_PAD_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.260 2945.000 940.540 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[54]
  PIN gfpga_pad_GPIO_PAD_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1488.240 3.930 1488.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[55]
  PIN gfpga_pad_GPIO_PAD_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1926.840 3.930 1927.440 ;
    END
  END gfpga_pad_GPIO_PAD_in[56]
  PIN gfpga_pad_GPIO_PAD_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 362.840 2808.930 363.440 ;
    END
  END gfpga_pad_GPIO_PAD_in[57]
  PIN gfpga_pad_GPIO_PAD_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.700 0.000 2073.980 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[58]
  PIN gfpga_pad_GPIO_PAD_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2202.240 2808.930 2202.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[59]
  PIN gfpga_pad_GPIO_PAD_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1399.840 3.930 1400.440 ;
    END
  END gfpga_pad_GPIO_PAD_in[5]
  PIN gfpga_pad_GPIO_PAD_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.720 0.000 1079.000 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[60]
  PIN gfpga_pad_GPIO_PAD_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.180 0.000 412.460 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[61]
  PIN gfpga_pad_GPIO_PAD_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.500 2945.000 2685.780 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[62]
  PIN gfpga_pad_GPIO_PAD_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1311.440 3.930 1312.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[63]
  PIN gfpga_pad_GPIO_PAD_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 349.240 3.930 349.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[6]
  PIN gfpga_pad_GPIO_PAD_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1590.240 2808.930 1590.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[7]
  PIN gfpga_pad_GPIO_PAD_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.320 2945.000 692.600 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[8]
  PIN gfpga_pad_GPIO_PAD_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2906.040 2808.930 2906.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[9]
  PIN gfpga_pad_GPIO_PAD_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2015.240 3.930 2015.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[0]
  PIN gfpga_pad_GPIO_PAD_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1750.040 3.930 1750.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[10]
  PIN gfpga_pad_GPIO_PAD_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.220 2945.000 193.500 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[11]
  PIN gfpga_pad_GPIO_PAD_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.540 2945.000 856.820 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[12]
  PIN gfpga_pad_GPIO_PAD_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.700 2945.000 1107.980 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[13]
  PIN gfpga_pad_GPIO_PAD_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2188.640 3.930 2189.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[14]
  PIN gfpga_pad_GPIO_PAD_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 434.240 3.930 434.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[15]
  PIN gfpga_pad_GPIO_PAD_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 974.840 2808.930 975.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[16]
  PIN gfpga_pad_GPIO_PAD_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2729.240 2808.930 2729.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[17]
  PIN gfpga_pad_GPIO_PAD_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.960 0.000 248.240 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[18]
  PIN gfpga_pad_GPIO_PAD_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 186.040 2808.930 186.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[19]
  PIN gfpga_pad_GPIO_PAD_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1063.240 2808.930 1063.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[1]
  PIN gfpga_pad_GPIO_PAD_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.460 2945.000 1938.740 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[20]
  PIN gfpga_pad_GPIO_PAD_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 624.640 2808.930 625.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[21]
  PIN gfpga_pad_GPIO_PAD_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2892.440 3.930 2893.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[22]
  PIN gfpga_pad_GPIO_PAD_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1576.640 3.930 1577.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[23]
  PIN gfpga_pad_GPIO_PAD_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1501.840 2808.930 1502.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[24]
  PIN gfpga_pad_GPIO_PAD_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2817.640 2808.930 2818.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[25]
  PIN gfpga_pad_GPIO_PAD_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1138.040 3.930 1138.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[26]
  PIN gfpga_pad_GPIO_PAD_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 447.840 2808.930 448.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[27]
  PIN gfpga_pad_GPIO_PAD_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.320 0.000 1658.600 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[28]
  PIN gfpga_pad_GPIO_PAD_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.520 0.000 2656.800 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[29]
  PIN gfpga_pad_GPIO_PAD_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.420 2945.000 1191.700 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[2]
  PIN gfpga_pad_GPIO_PAD_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.420 0.000 2157.700 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[30]
  PIN gfpga_pad_GPIO_PAD_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.680 0.000 331.960 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[31]
  PIN gfpga_pad_GPIO_PAD_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1049.640 3.930 1050.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[32]
  PIN gfpga_pad_GPIO_PAD_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 274.440 2808.930 275.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[33]
  PIN gfpga_pad_GPIO_PAD_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2113.840 2808.930 2114.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[34]
  PIN gfpga_pad_GPIO_PAD_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 84.040 3.930 84.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[35]
  PIN gfpga_pad_GPIO_PAD_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.860 0.000 2325.140 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[36]
  PIN gfpga_pad_GPIO_PAD_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 1838.440 3.930 1839.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[37]
  PIN gfpga_pad_GPIO_PAD_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 713.040 2808.930 713.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[38]
  PIN gfpga_pad_GPIO_PAD_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2453.840 3.930 2454.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[39]
  PIN gfpga_pad_GPIO_PAD_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1678.640 2808.930 1679.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[3]
  PIN gfpga_pad_GPIO_PAD_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2467.440 2808.930 2468.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[40]
  PIN gfpga_pad_GPIO_PAD_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2572.800 0.000 2573.080 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[41]
  PIN gfpga_pad_GPIO_PAD_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 2640.840 2808.930 2641.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[42]
  PIN gfpga_pad_GPIO_PAD_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 172.440 3.930 173.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[43]
  PIN gfpga_pad_GPIO_PAD_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2627.240 3.930 2627.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[44]
  PIN gfpga_pad_GPIO_PAD_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 961.240 3.930 961.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[45]
  PIN gfpga_pad_GPIO_PAD_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[46]
  PIN gfpga_pad_GPIO_PAD_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.480 0.000 1909.760 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[47]
  PIN gfpga_pad_GPIO_PAD_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2804.040 3.930 2804.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[48]
  PIN gfpga_pad_GPIO_PAD_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.040 2945.000 776.320 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[49]
  PIN gfpga_pad_GPIO_PAD_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.020 2945.000 1771.300 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[4]
  PIN gfpga_pad_GPIO_PAD_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2277.040 3.930 2277.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[50]
  PIN gfpga_pad_GPIO_PAD_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.900 0.000 496.180 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[51]
  PIN gfpga_pad_GPIO_PAD_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.240 0.000 164.520 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[52]
  PIN gfpga_pad_GPIO_PAD_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.400 2945.000 2186.680 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[53]
  PIN gfpga_pad_GPIO_PAD_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.800 2945.000 1607.080 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[54]
  PIN gfpga_pad_GPIO_PAD_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.660 0.000 1326.940 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[55]
  PIN gfpga_pad_GPIO_PAD_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.060 2945.000 2518.340 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[56]
  PIN gfpga_pad_GPIO_PAD_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 536.240 2808.930 536.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[57]
  PIN gfpga_pad_GPIO_PAD_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2715.640 3.930 2716.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[58]
  PIN gfpga_pad_GPIO_PAD_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 872.840 3.930 873.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[59]
  PIN gfpga_pad_GPIO_PAD_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.620 0.000 579.900 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[5]
  PIN gfpga_pad_GPIO_PAD_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.000 0.000 995.280 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[60]
  PIN gfpga_pad_GPIO_PAD_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 260.840 3.930 261.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[61]
  PIN gfpga_pad_GPIO_PAD_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1940.440 2808.930 1941.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[62]
  PIN gfpga_pad_GPIO_PAD_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.820 0.000 1578.100 3.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[63]
  PIN gfpga_pad_GPIO_PAD_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.680 2945.000 2102.960 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[6]
  PIN gfpga_pad_GPIO_PAD_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.960 2945.000 2019.240 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[7]
  PIN gfpga_pad_GPIO_PAD_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.780 2945.000 26.060 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[8]
  PIN gfpga_pad_GPIO_PAD_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.880 2945.000 525.160 2948.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[9]
  PIN pReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.200 0.000 1993.480 3.000 ;
    END
  END pReset
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 787.840 3.930 788.440 ;
    END
  END prog_clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.930 2538.840 3.930 2539.440 ;
    END
  END reset
  PIN set
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2805.930 1413.440 2808.930 1414.040 ;
    END
  END set
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 41.650 9.640 43.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.650 9.640 113.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.650 9.640 183.250 302.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.650 492.045 183.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.650 9.640 253.250 302.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.650 492.045 253.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.650 9.640 323.250 554.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.650 746.125 323.250 1064.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.650 1256.125 323.250 1574.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.650 1766.125 323.250 2151.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.650 2248.245 323.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.650 9.640 393.250 554.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.650 746.125 393.250 1064.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.650 1256.125 393.250 1574.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.650 1766.125 393.250 2151.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.650 2248.245 393.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.650 9.640 463.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.650 9.640 533.250 799.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.650 1016.260 533.250 1309.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.650 1526.260 533.250 1819.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.650 2036.260 533.250 2329.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.650 2546.260 533.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.650 9.640 603.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.650 989.325 603.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.650 1499.325 603.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.650 2009.325 603.250 2080.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.650 2274.765 603.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.650 2519.325 603.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.650 9.640 673.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.650 989.325 673.250 1064.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.650 1124.885 673.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.650 1499.325 673.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.650 2009.325 673.250 2080.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.650 2274.765 673.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.650 2519.325 673.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.650 9.640 743.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.650 9.640 813.250 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.650 482.525 813.250 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.650 732.325 813.250 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.650 1242.325 813.250 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.650 1752.325 813.250 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.650 2244.645 813.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.650 9.640 883.250 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.650 482.525 883.250 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.650 732.325 883.250 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.650 1242.325 883.250 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.650 1752.325 883.250 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.650 2244.645 883.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.650 9.640 953.250 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.650 732.325 953.250 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.650 1242.325 953.250 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.650 1752.325 953.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.650 9.640 1023.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.650 989.325 1023.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.650 1499.325 1023.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.650 2009.325 1023.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.650 2519.325 1023.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.650 9.640 1093.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.650 989.325 1093.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.650 1499.325 1093.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.650 2009.325 1093.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.650 2519.325 1093.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 9.640 1163.250 281.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 377.525 1163.250 554.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 614.885 1163.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 989.325 1163.250 1064.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 1124.885 1163.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 1499.325 1163.250 1574.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 1634.885 1163.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 2009.325 1163.250 2080.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 2274.765 1163.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.650 2519.325 1163.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.650 9.640 1233.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.650 9.640 1303.250 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.650 482.525 1303.250 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.650 732.325 1303.250 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.650 1242.325 1303.250 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.650 1752.325 1303.250 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.650 2244.645 1303.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.650 9.640 1373.250 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.650 482.525 1373.250 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.650 732.325 1373.250 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.650 1242.325 1373.250 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.650 1752.325 1373.250 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.650 2244.645 1373.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.650 9.640 1443.250 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.650 732.325 1443.250 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.650 1242.325 1443.250 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.650 1752.325 1443.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1511.650 9.640 1513.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.650 9.640 1583.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.650 989.325 1583.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.650 1499.325 1583.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.650 2009.325 1583.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.650 2519.325 1583.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.650 9.640 1653.250 281.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.650 377.525 1653.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.650 989.325 1653.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.650 1499.325 1653.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.650 2009.325 1653.250 2080.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.650 2274.765 1653.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.650 2519.325 1653.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.650 9.640 1723.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.650 989.325 1723.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.650 1499.325 1723.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.650 2009.325 1723.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.650 2519.325 1723.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1791.650 9.640 1793.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.650 9.640 1863.250 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.650 482.525 1863.250 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.650 732.325 1863.250 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.650 1242.325 1863.250 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.650 1752.325 1863.250 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.650 2244.645 1863.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.650 9.640 1933.250 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.650 482.525 1933.250 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.650 732.325 1933.250 826.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.650 927.445 1933.250 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.650 1242.325 1933.250 1336.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.650 1437.445 1933.250 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.650 1752.325 1933.250 1846.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.650 1947.445 1933.250 2356.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.650 2457.445 1933.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2001.650 9.640 2003.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.650 9.640 2073.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.650 989.325 2073.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.650 1499.325 2073.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.650 2009.325 2073.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.650 2519.325 2073.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.650 9.640 2143.250 281.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.650 377.525 2143.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.650 989.325 2143.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.650 1499.325 2143.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.650 2009.325 2143.250 2080.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.650 2274.765 2143.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.650 2519.325 2143.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.650 9.640 2213.250 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.650 989.325 2213.250 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.650 1499.325 2213.250 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.650 2009.325 2213.250 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.650 2519.325 2213.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.650 9.640 2283.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.650 9.640 2353.250 308.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.650 492.725 2353.250 541.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.650 729.325 2353.250 774.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.650 868.645 2353.250 1021.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.650 1209.325 2353.250 1284.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.650 1378.645 2353.250 1531.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.650 1719.325 2353.250 1794.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.650 1888.645 2353.250 2304.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.650 2398.645 2353.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.650 9.640 2423.250 308.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.650 492.725 2423.250 541.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.650 729.325 2423.250 1021.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.650 1209.325 2423.250 1531.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.650 1719.325 2423.250 2043.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.650 2176.285 2423.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2491.650 9.640 2493.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2561.650 9.640 2563.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2631.650 9.640 2633.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2701.650 9.640 2703.250 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2771.650 9.640 2773.250 2936.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 46.080 2804.330 47.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 121.080 2804.330 122.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 196.080 2804.330 197.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 271.080 2804.330 272.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 346.080 2804.330 347.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 421.080 2804.330 422.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 496.080 2804.330 497.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 571.080 2804.330 572.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 646.080 2804.330 647.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 721.080 2804.330 722.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 796.080 2804.330 797.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 871.080 2804.330 872.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 946.080 2804.330 947.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1021.080 2804.330 1022.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1096.080 2804.330 1097.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1171.080 2804.330 1172.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1246.080 2804.330 1247.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1321.080 2804.330 1322.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1396.080 2804.330 1397.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1471.080 2804.330 1472.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1546.080 2804.330 1547.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1621.080 2804.330 1622.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1696.080 2804.330 1697.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1771.080 2804.330 1772.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1846.080 2804.330 1847.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1921.080 2804.330 1922.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1996.080 2804.330 1997.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2071.080 2804.330 2072.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2146.080 2804.330 2147.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2221.080 2804.330 2222.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2296.080 2804.330 2297.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2371.080 2804.330 2372.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2446.080 2804.330 2447.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2521.080 2804.330 2522.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2596.080 2804.330 2597.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2671.080 2804.330 2672.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2746.080 2804.330 2747.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2821.080 2804.330 2822.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2896.080 2804.330 2897.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.470 523.720 14.070 752.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 512.030 1045.960 513.630 1272.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1256.310 1568.200 1257.910 1780.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.070 2074.120 1766.670 2292.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.150 784.840 2018.750 804.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.350 1274.440 2533.950 1487.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2789.950 1785.800 2791.550 2012.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.470 1035.080 14.070 1264.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.670 534.600 506.270 763.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 997.790 784.840 999.390 1013.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1256.310 2074.120 1257.910 2292.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.070 1565.480 1766.670 1783.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.510 284.360 2026.110 494.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.350 1785.800 2533.950 1998.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2789.950 1274.440 2791.550 1503.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.470 1543.720 14.070 1772.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.670 2065.960 506.270 2292.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1256.310 1056.840 1257.910 1269.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1769.670 284.360 1771.270 494.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.150 804.660 2018.750 1013.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.350 2294.440 2533.950 2507.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.470 2055.080 14.070 2284.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.670 1554.600 506.270 1783.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1256.310 545.480 1257.910 763.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.430 784.840 1774.030 1013.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.150 1293.480 2018.750 1313.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2789.950 2294.440 2791.550 2523.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 997.790 1293.480 999.390 1522.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.990 284.360 1261.590 494.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.070 545.480 1766.670 774.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.510 1054.120 2026.110 1277.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.750 784.840 1264.350 1013.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.070 1054.120 1766.670 1272.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.510 545.480 2026.110 763.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 997.790 1804.840 999.390 2033.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.750 1293.480 1264.350 1522.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.430 2313.480 1774.030 2542.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.510 1565.480 2026.110 1783.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.350 765.800 2533.950 978.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.750 1804.840 1264.350 2033.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.430 1293.480 1774.030 1522.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.150 2313.480 2018.750 2333.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2789.950 765.800 2791.550 992.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 997.790 2313.480 999.390 2542.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.430 1804.840 1774.030 2033.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.150 1313.300 2018.750 1522.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 2281.650 747.900 2426.550 749.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.750 2313.480 1264.350 2542.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.150 1804.840 2018.750 1824.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.150 1824.660 2018.750 2033.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.510 2074.120 2026.110 2292.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.150 2333.300 2018.750 2542.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 44.950 9.640 46.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.950 9.640 116.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.950 9.640 186.550 302.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.950 492.045 186.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.950 9.640 256.550 302.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.950 492.045 256.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.950 9.640 326.550 554.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.950 746.125 326.550 1064.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.950 1256.125 326.550 1574.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.950 1766.125 326.550 2151.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.950 2248.245 326.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.950 9.640 396.550 554.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.950 746.125 396.550 1064.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.950 1256.125 396.550 1574.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.950 1766.125 396.550 2151.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.950 2248.245 396.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.950 9.640 466.550 549.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.950 747.220 466.550 1059.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.950 1257.220 466.550 1569.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.950 1767.220 466.550 2079.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.950 2277.220 466.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.950 9.640 536.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.950 989.325 536.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.950 1499.325 536.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.950 2009.325 536.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.950 2519.325 536.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.950 9.640 606.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.950 989.325 606.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.950 1499.325 606.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.950 2009.325 606.550 2080.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.950 2274.765 606.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.950 2519.325 606.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.950 9.640 676.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.950 989.325 676.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.950 1499.325 676.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.950 2009.325 676.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.950 2519.325 676.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.950 9.640 746.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.950 9.640 816.550 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.950 482.525 816.550 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.950 732.325 816.550 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.950 1242.325 816.550 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.950 1752.325 816.550 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.950 2244.645 816.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 884.950 9.640 886.550 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 884.950 482.525 886.550 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 884.950 732.325 886.550 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 884.950 1242.325 886.550 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 884.950 1752.325 886.550 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 884.950 2244.645 886.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 9.640 956.550 299.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 497.220 956.550 559.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 757.220 956.550 799.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 997.220 956.550 1069.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 1267.220 956.550 1309.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 1507.220 956.550 1579.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 1777.220 956.550 1819.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 2017.220 956.550 2089.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 2287.220 956.550 2329.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.950 2527.220 956.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1024.950 9.640 1026.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1024.950 989.325 1026.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1024.950 1499.325 1026.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1024.950 2009.325 1026.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1024.950 2519.325 1026.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1094.950 9.640 1096.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1094.950 989.325 1096.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1094.950 1499.325 1096.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1094.950 2009.325 1096.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1094.950 2519.325 1096.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.950 9.640 1166.550 554.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.950 614.885 1166.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.950 989.325 1166.550 1064.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.950 1124.885 1166.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.950 1499.325 1166.550 1574.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.950 1634.885 1166.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.950 2009.325 1166.550 2080.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.950 2274.765 1166.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.950 2519.325 1166.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.950 9.640 1236.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.950 9.640 1306.550 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.950 482.525 1306.550 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.950 732.325 1306.550 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.950 1242.325 1306.550 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.950 1752.325 1306.550 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.950 2244.645 1306.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.950 9.640 1376.550 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.950 482.525 1376.550 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.950 732.325 1376.550 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.950 1242.325 1376.550 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.950 1752.325 1376.550 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.950 2244.645 1376.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.950 9.640 1446.550 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.950 732.325 1446.550 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.950 1242.325 1446.550 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1444.950 1752.325 1446.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1514.950 9.640 1516.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.950 9.640 1586.550 29.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.950 227.220 1586.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.950 989.325 1586.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.950 1499.325 1586.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.950 2009.325 1586.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.950 2519.325 1586.550 2609.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1584.950 2807.220 1586.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.950 9.640 1656.550 281.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.950 377.525 1656.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.950 989.325 1656.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.950 1499.325 1656.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.950 2009.325 1656.550 2080.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.950 2274.765 1656.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.950 2519.325 1656.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1724.950 9.640 1726.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1724.950 989.325 1726.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1724.950 1499.325 1726.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1724.950 2009.325 1726.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 1724.950 2519.325 1726.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1794.950 9.640 1796.550 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1794.950 2244.645 1796.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.950 9.640 1866.550 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.950 482.525 1866.550 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.950 732.325 1866.550 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.950 1242.325 1866.550 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.950 1752.325 1866.550 2091.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.950 2244.645 1866.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.950 9.640 1936.550 335.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.950 482.525 1936.550 560.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.950 732.325 1936.550 826.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.950 927.445 1936.550 1070.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.950 1242.325 1936.550 1336.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.950 1437.445 1936.550 1580.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.950 1752.325 1936.550 1846.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.950 1947.445 1936.550 2356.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.950 2457.445 1936.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.950 9.640 2006.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 9.640 2076.550 279.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 477.220 2076.550 549.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 747.220 2076.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 989.325 2076.550 1062.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 1260.220 2076.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 1499.325 2076.550 1569.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 1767.220 2076.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 2009.325 2076.550 2079.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 2277.220 2076.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2074.950 2519.325 2076.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.950 9.640 2146.550 281.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.950 377.525 2146.550 803.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.950 989.325 2146.550 1313.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.950 1499.325 2146.550 1823.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.950 2009.325 2146.550 2080.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.950 2274.765 2146.550 2333.835 ;
    END
    PORT
      LAYER met4 ;
        RECT 2144.950 2519.325 2146.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.950 9.640 2216.550 799.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.950 1016.260 2216.550 1309.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.950 1526.260 2216.550 1819.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.950 2036.260 2216.550 2329.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.950 2546.260 2216.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2284.950 9.640 2286.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.950 9.640 2356.550 308.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.950 492.725 2356.550 541.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.950 729.325 2356.550 774.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.950 868.645 2356.550 1021.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.950 1209.325 2356.550 1284.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.950 1378.645 2356.550 1531.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.950 1719.325 2356.550 1794.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.950 1888.645 2356.550 2304.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.950 2398.645 2356.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2424.950 9.640 2426.550 308.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2424.950 492.725 2426.550 541.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2424.950 729.325 2426.550 1021.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2424.950 1209.325 2426.550 1531.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2424.950 1719.325 2426.550 2039.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2424.950 2188.260 2426.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.950 9.640 2496.550 2039.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.950 2188.260 2496.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2564.950 9.640 2566.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2634.950 9.640 2636.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.950 9.640 2706.550 2936.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2774.950 9.640 2776.550 2936.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 49.380 2804.330 50.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 124.380 2804.330 125.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 199.380 2804.330 200.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 274.380 2804.330 275.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 349.380 2804.330 350.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 424.380 2804.330 425.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 499.380 2804.330 500.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 574.380 2804.330 575.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 649.380 2804.330 650.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 724.380 2804.330 725.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 799.380 2804.330 800.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 874.380 2804.330 875.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 949.380 2804.330 950.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1024.380 2804.330 1025.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1099.380 2804.330 1100.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1174.380 2804.330 1175.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1249.380 2804.330 1250.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1324.380 2804.330 1325.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1399.380 2804.330 1400.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1474.380 2804.330 1475.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1549.380 2804.330 1550.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1624.380 2804.330 1625.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1699.380 2804.330 1700.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1774.380 2804.330 1775.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1849.380 2804.330 1850.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1924.380 2804.330 1925.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 1999.380 2804.330 2000.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2074.380 2804.330 2075.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2149.380 2804.330 2150.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2224.380 2804.330 2225.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2299.380 2804.330 2300.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2374.380 2804.330 2375.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2449.380 2804.330 2450.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2524.380 2804.330 2525.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2599.380 2804.330 2600.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2674.380 2804.330 2675.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2749.380 2804.330 2750.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2824.380 2804.330 2825.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.210 2899.380 2804.330 2900.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.150 523.720 17.750 752.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 515.710 1045.960 517.310 1272.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1006.990 287.080 1008.590 494.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.750 2074.120 1770.350 2292.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.830 784.840 2022.430 804.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.030 1274.440 2537.630 1487.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2793.630 1785.800 2795.230 2012.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.150 1035.080 17.750 1264.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.350 534.600 509.950 763.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.470 784.840 1003.070 1013.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.750 1565.480 1770.350 1783.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.190 284.360 2029.790 494.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.030 1785.800 2537.630 1998.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2793.630 1274.440 2795.230 1503.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.150 1543.720 17.750 1772.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.350 2065.960 509.950 2292.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1006.990 548.200 1008.590 760.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1773.350 284.360 1774.950 494.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.830 804.660 2022.430 1013.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.030 2294.440 2537.630 2507.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.150 2055.080 17.750 2284.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.350 1554.600 509.950 1783.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1006.990 1054.120 1008.590 1272.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.110 784.840 1777.710 1013.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.830 1293.480 2022.430 1313.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2793.630 2294.440 2795.230 2523.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.470 1293.480 1003.070 1522.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.670 284.360 1265.270 494.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.750 545.480 1770.350 774.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.190 1054.120 2029.790 1277.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1006.990 1565.480 1008.590 1783.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1266.430 784.840 1268.030 1013.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.750 1054.120 1770.350 1272.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.190 545.480 2029.790 763.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.470 1804.840 1003.070 2033.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1266.430 1293.480 1268.030 1522.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.110 2313.480 1777.710 2542.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.190 1565.480 2029.790 1783.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.030 765.800 2537.630 978.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1006.990 2076.840 1008.590 2289.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1266.430 1804.840 1268.030 2033.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.110 1293.480 1777.710 1522.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.830 2313.480 2022.430 2333.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2793.630 765.800 2795.230 992.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.470 2313.480 1003.070 2542.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.110 1804.840 1777.710 2033.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.830 1313.300 2022.430 1522.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 2281.650 751.300 2426.550 752.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1266.430 2313.480 1268.030 2542.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.830 1804.840 2022.430 1824.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.830 1824.660 2022.430 2033.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.190 2074.120 2029.790 2292.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.830 2333.300 2022.430 2542.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.450 9.795 2804.090 2936.685 ;
      LAYER met1 ;
        RECT 0.000 7.880 2804.390 2936.840 ;
      LAYER met2 ;
        RECT 0.030 2944.720 25.500 2945.170 ;
        RECT 26.340 2944.720 109.220 2945.170 ;
        RECT 110.060 2944.720 192.940 2945.170 ;
        RECT 193.780 2944.720 276.660 2945.170 ;
        RECT 277.500 2944.720 360.380 2945.170 ;
        RECT 361.220 2944.720 440.880 2945.170 ;
        RECT 441.720 2944.720 524.600 2945.170 ;
        RECT 525.440 2944.720 608.320 2945.170 ;
        RECT 609.160 2944.720 692.040 2945.170 ;
        RECT 692.880 2944.720 775.760 2945.170 ;
        RECT 776.600 2944.720 856.260 2945.170 ;
        RECT 857.100 2944.720 939.980 2945.170 ;
        RECT 940.820 2944.720 1023.700 2945.170 ;
        RECT 1024.540 2944.720 1107.420 2945.170 ;
        RECT 1108.260 2944.720 1191.140 2945.170 ;
        RECT 1191.980 2944.720 1271.640 2945.170 ;
        RECT 1272.480 2944.720 1355.360 2945.170 ;
        RECT 1356.200 2944.720 1439.080 2945.170 ;
        RECT 1439.920 2944.720 1522.800 2945.170 ;
        RECT 1523.640 2944.720 1606.520 2945.170 ;
        RECT 1607.360 2944.720 1687.020 2945.170 ;
        RECT 1687.860 2944.720 1770.740 2945.170 ;
        RECT 1771.580 2944.720 1854.460 2945.170 ;
        RECT 1855.300 2944.720 1938.180 2945.170 ;
        RECT 1939.020 2944.720 2018.680 2945.170 ;
        RECT 2019.520 2944.720 2102.400 2945.170 ;
        RECT 2103.240 2944.720 2186.120 2945.170 ;
        RECT 2186.960 2944.720 2269.840 2945.170 ;
        RECT 2270.680 2944.720 2353.560 2945.170 ;
        RECT 2354.400 2944.720 2434.060 2945.170 ;
        RECT 2434.900 2944.720 2517.780 2945.170 ;
        RECT 2518.620 2944.720 2601.500 2945.170 ;
        RECT 2602.340 2944.720 2685.220 2945.170 ;
        RECT 2686.060 2944.720 2768.940 2945.170 ;
        RECT 2769.780 2944.720 2801.690 2945.170 ;
        RECT 0.030 3.280 2801.690 2944.720 ;
        RECT 0.580 2.670 80.240 3.280 ;
        RECT 81.080 2.670 163.960 3.280 ;
        RECT 164.800 2.670 247.680 3.280 ;
        RECT 248.520 2.670 331.400 3.280 ;
        RECT 332.240 2.670 411.900 3.280 ;
        RECT 412.740 2.670 495.620 3.280 ;
        RECT 496.460 2.670 579.340 3.280 ;
        RECT 580.180 2.670 663.060 3.280 ;
        RECT 663.900 2.670 746.780 3.280 ;
        RECT 747.620 2.670 827.280 3.280 ;
        RECT 828.120 2.670 911.000 3.280 ;
        RECT 911.840 2.670 994.720 3.280 ;
        RECT 995.560 2.670 1078.440 3.280 ;
        RECT 1079.280 2.670 1162.160 3.280 ;
        RECT 1163.000 2.670 1242.660 3.280 ;
        RECT 1243.500 2.670 1326.380 3.280 ;
        RECT 1327.220 2.670 1410.100 3.280 ;
        RECT 1410.940 2.670 1493.820 3.280 ;
        RECT 1494.660 2.670 1577.540 3.280 ;
        RECT 1578.380 2.670 1658.040 3.280 ;
        RECT 1658.880 2.670 1741.760 3.280 ;
        RECT 1742.600 2.670 1825.480 3.280 ;
        RECT 1826.320 2.670 1909.200 3.280 ;
        RECT 1910.040 2.670 1992.920 3.280 ;
        RECT 1993.760 2.670 2073.420 3.280 ;
        RECT 2074.260 2.670 2157.140 3.280 ;
        RECT 2157.980 2.670 2240.860 3.280 ;
        RECT 2241.700 2.670 2324.580 3.280 ;
        RECT 2325.420 2.670 2405.080 3.280 ;
        RECT 2405.920 2.670 2488.800 3.280 ;
        RECT 2489.640 2.670 2572.520 3.280 ;
        RECT 2573.360 2.670 2656.240 3.280 ;
        RECT 2657.080 2.670 2739.960 3.280 ;
        RECT 2740.800 2.670 2801.690 3.280 ;
      LAYER met3 ;
        RECT 3.930 2907.040 2805.930 2936.765 ;
        RECT 3.930 2905.640 2805.530 2907.040 ;
        RECT 3.930 2893.440 2805.930 2905.640 ;
        RECT 4.330 2892.040 2805.930 2893.440 ;
        RECT 3.930 2818.640 2805.930 2892.040 ;
        RECT 3.930 2817.240 2805.530 2818.640 ;
        RECT 3.930 2805.040 2805.930 2817.240 ;
        RECT 4.330 2803.640 2805.930 2805.040 ;
        RECT 3.930 2730.240 2805.930 2803.640 ;
        RECT 3.930 2728.840 2805.530 2730.240 ;
        RECT 3.930 2716.640 2805.930 2728.840 ;
        RECT 4.330 2715.240 2805.930 2716.640 ;
        RECT 3.930 2641.840 2805.930 2715.240 ;
        RECT 3.930 2640.440 2805.530 2641.840 ;
        RECT 3.930 2628.240 2805.930 2640.440 ;
        RECT 4.330 2626.840 2805.930 2628.240 ;
        RECT 3.930 2553.440 2805.930 2626.840 ;
        RECT 3.930 2552.040 2805.530 2553.440 ;
        RECT 3.930 2539.840 2805.930 2552.040 ;
        RECT 4.330 2538.440 2805.930 2539.840 ;
        RECT 3.930 2468.440 2805.930 2538.440 ;
        RECT 3.930 2467.040 2805.530 2468.440 ;
        RECT 3.930 2454.840 2805.930 2467.040 ;
        RECT 4.330 2453.440 2805.930 2454.840 ;
        RECT 3.930 2380.040 2805.930 2453.440 ;
        RECT 3.930 2378.640 2805.530 2380.040 ;
        RECT 3.930 2366.440 2805.930 2378.640 ;
        RECT 4.330 2365.040 2805.930 2366.440 ;
        RECT 3.930 2291.640 2805.930 2365.040 ;
        RECT 3.930 2290.240 2805.530 2291.640 ;
        RECT 3.930 2278.040 2805.930 2290.240 ;
        RECT 4.330 2276.640 2805.930 2278.040 ;
        RECT 3.930 2203.240 2805.930 2276.640 ;
        RECT 3.930 2201.840 2805.530 2203.240 ;
        RECT 3.930 2189.640 2805.930 2201.840 ;
        RECT 4.330 2188.240 2805.930 2189.640 ;
        RECT 3.930 2114.840 2805.930 2188.240 ;
        RECT 3.930 2113.440 2805.530 2114.840 ;
        RECT 3.930 2104.640 2805.930 2113.440 ;
        RECT 4.330 2103.240 2805.930 2104.640 ;
        RECT 3.930 2029.840 2805.930 2103.240 ;
        RECT 3.930 2028.440 2805.530 2029.840 ;
        RECT 3.930 2016.240 2805.930 2028.440 ;
        RECT 4.330 2014.840 2805.930 2016.240 ;
        RECT 3.930 1941.440 2805.930 2014.840 ;
        RECT 3.930 1940.040 2805.530 1941.440 ;
        RECT 3.930 1927.840 2805.930 1940.040 ;
        RECT 4.330 1926.440 2805.930 1927.840 ;
        RECT 3.930 1853.040 2805.930 1926.440 ;
        RECT 3.930 1851.640 2805.530 1853.040 ;
        RECT 3.930 1839.440 2805.930 1851.640 ;
        RECT 4.330 1838.040 2805.930 1839.440 ;
        RECT 3.930 1764.640 2805.930 1838.040 ;
        RECT 3.930 1763.240 2805.530 1764.640 ;
        RECT 3.930 1751.040 2805.930 1763.240 ;
        RECT 4.330 1749.640 2805.930 1751.040 ;
        RECT 3.930 1679.640 2805.930 1749.640 ;
        RECT 3.930 1678.240 2805.530 1679.640 ;
        RECT 3.930 1666.040 2805.930 1678.240 ;
        RECT 4.330 1664.640 2805.930 1666.040 ;
        RECT 3.930 1591.240 2805.930 1664.640 ;
        RECT 3.930 1589.840 2805.530 1591.240 ;
        RECT 3.930 1577.640 2805.930 1589.840 ;
        RECT 4.330 1576.240 2805.930 1577.640 ;
        RECT 3.930 1502.840 2805.930 1576.240 ;
        RECT 3.930 1501.440 2805.530 1502.840 ;
        RECT 3.930 1489.240 2805.930 1501.440 ;
        RECT 4.330 1487.840 2805.930 1489.240 ;
        RECT 3.930 1414.440 2805.930 1487.840 ;
        RECT 3.930 1413.040 2805.530 1414.440 ;
        RECT 3.930 1400.840 2805.930 1413.040 ;
        RECT 4.330 1399.440 2805.930 1400.840 ;
        RECT 3.930 1326.040 2805.930 1399.440 ;
        RECT 3.930 1324.640 2805.530 1326.040 ;
        RECT 3.930 1312.440 2805.930 1324.640 ;
        RECT 4.330 1311.040 2805.930 1312.440 ;
        RECT 3.930 1241.040 2805.930 1311.040 ;
        RECT 3.930 1239.640 2805.530 1241.040 ;
        RECT 3.930 1227.440 2805.930 1239.640 ;
        RECT 4.330 1226.040 2805.930 1227.440 ;
        RECT 3.930 1152.640 2805.930 1226.040 ;
        RECT 3.930 1151.240 2805.530 1152.640 ;
        RECT 3.930 1139.040 2805.930 1151.240 ;
        RECT 4.330 1137.640 2805.930 1139.040 ;
        RECT 3.930 1064.240 2805.930 1137.640 ;
        RECT 3.930 1062.840 2805.530 1064.240 ;
        RECT 3.930 1050.640 2805.930 1062.840 ;
        RECT 4.330 1049.240 2805.930 1050.640 ;
        RECT 3.930 975.840 2805.930 1049.240 ;
        RECT 3.930 974.440 2805.530 975.840 ;
        RECT 3.930 962.240 2805.930 974.440 ;
        RECT 4.330 960.840 2805.930 962.240 ;
        RECT 3.930 887.440 2805.930 960.840 ;
        RECT 3.930 886.040 2805.530 887.440 ;
        RECT 3.930 873.840 2805.930 886.040 ;
        RECT 4.330 872.440 2805.930 873.840 ;
        RECT 3.930 802.440 2805.930 872.440 ;
        RECT 3.930 801.040 2805.530 802.440 ;
        RECT 3.930 788.840 2805.930 801.040 ;
        RECT 4.330 787.440 2805.930 788.840 ;
        RECT 3.930 714.040 2805.930 787.440 ;
        RECT 3.930 712.640 2805.530 714.040 ;
        RECT 3.930 700.440 2805.930 712.640 ;
        RECT 4.330 699.040 2805.930 700.440 ;
        RECT 3.930 625.640 2805.930 699.040 ;
        RECT 3.930 624.240 2805.530 625.640 ;
        RECT 3.930 612.040 2805.930 624.240 ;
        RECT 4.330 610.640 2805.930 612.040 ;
        RECT 3.930 537.240 2805.930 610.640 ;
        RECT 3.930 535.840 2805.530 537.240 ;
        RECT 3.930 523.640 2805.930 535.840 ;
        RECT 4.330 522.240 2805.930 523.640 ;
        RECT 3.930 448.840 2805.930 522.240 ;
        RECT 3.930 447.440 2805.530 448.840 ;
        RECT 3.930 435.240 2805.930 447.440 ;
        RECT 4.330 433.840 2805.930 435.240 ;
        RECT 3.930 363.840 2805.930 433.840 ;
        RECT 3.930 362.440 2805.530 363.840 ;
        RECT 3.930 350.240 2805.930 362.440 ;
        RECT 4.330 348.840 2805.930 350.240 ;
        RECT 3.930 275.440 2805.930 348.840 ;
        RECT 3.930 274.040 2805.530 275.440 ;
        RECT 3.930 261.840 2805.930 274.040 ;
        RECT 4.330 260.440 2805.930 261.840 ;
        RECT 3.930 187.040 2805.930 260.440 ;
        RECT 3.930 185.640 2805.530 187.040 ;
        RECT 3.930 173.440 2805.930 185.640 ;
        RECT 4.330 172.040 2805.930 173.440 ;
        RECT 3.930 98.640 2805.930 172.040 ;
        RECT 3.930 97.240 2805.530 98.640 ;
        RECT 3.930 85.040 2805.930 97.240 ;
        RECT 4.330 83.640 2805.930 85.040 ;
        RECT 3.930 10.240 2805.930 83.640 ;
        RECT 3.930 8.840 2805.530 10.240 ;
        RECT 3.930 8.695 2805.930 8.840 ;
      LAYER met4 ;
        RECT 26.905 9.240 41.250 2935.745 ;
        RECT 43.650 9.240 44.550 2935.745 ;
        RECT 46.950 9.240 111.250 2935.745 ;
        RECT 113.650 9.240 114.550 2935.745 ;
        RECT 116.950 491.645 181.250 2935.745 ;
        RECT 183.650 491.645 184.550 2935.745 ;
        RECT 186.950 491.645 251.250 2935.745 ;
        RECT 253.650 491.645 254.550 2935.745 ;
        RECT 256.950 2247.845 321.250 2935.745 ;
        RECT 323.650 2247.845 324.550 2935.745 ;
        RECT 326.950 2247.845 391.250 2935.745 ;
        RECT 393.650 2247.845 394.550 2935.745 ;
        RECT 396.950 2247.845 461.250 2935.745 ;
        RECT 256.950 2151.555 461.250 2247.845 ;
        RECT 256.950 1765.725 321.250 2151.555 ;
        RECT 323.650 1765.725 324.550 2151.555 ;
        RECT 326.950 1765.725 391.250 2151.555 ;
        RECT 393.650 1765.725 394.550 2151.555 ;
        RECT 396.950 1765.725 461.250 2151.555 ;
        RECT 256.950 1574.915 461.250 1765.725 ;
        RECT 256.950 1255.725 321.250 1574.915 ;
        RECT 323.650 1255.725 324.550 1574.915 ;
        RECT 326.950 1255.725 391.250 1574.915 ;
        RECT 393.650 1255.725 394.550 1574.915 ;
        RECT 396.950 1255.725 461.250 1574.915 ;
        RECT 256.950 1064.915 461.250 1255.725 ;
        RECT 256.950 745.725 321.250 1064.915 ;
        RECT 323.650 745.725 324.550 1064.915 ;
        RECT 326.950 745.725 391.250 1064.915 ;
        RECT 393.650 745.725 394.550 1064.915 ;
        RECT 396.950 745.725 461.250 1064.915 ;
        RECT 256.950 554.915 461.250 745.725 ;
        RECT 256.950 491.645 321.250 554.915 ;
        RECT 116.950 302.875 321.250 491.645 ;
        RECT 116.950 9.240 181.250 302.875 ;
        RECT 183.650 9.240 184.550 302.875 ;
        RECT 186.950 9.240 251.250 302.875 ;
        RECT 253.650 9.240 254.550 302.875 ;
        RECT 256.950 9.240 321.250 302.875 ;
        RECT 323.650 9.240 324.550 554.915 ;
        RECT 326.950 9.240 391.250 554.915 ;
        RECT 393.650 9.240 394.550 554.915 ;
        RECT 396.950 9.240 461.250 554.915 ;
        RECT 463.650 2276.820 464.550 2935.745 ;
        RECT 466.950 2545.860 531.250 2935.745 ;
        RECT 533.650 2545.860 534.550 2935.745 ;
        RECT 466.950 2518.925 534.550 2545.860 ;
        RECT 536.950 2518.925 601.250 2935.745 ;
        RECT 603.650 2518.925 604.550 2935.745 ;
        RECT 606.950 2518.925 671.250 2935.745 ;
        RECT 673.650 2518.925 674.550 2935.745 ;
        RECT 676.950 2518.925 741.250 2935.745 ;
        RECT 466.950 2334.235 741.250 2518.925 ;
        RECT 466.950 2329.740 534.550 2334.235 ;
        RECT 466.950 2292.600 531.250 2329.740 ;
        RECT 466.950 2276.820 504.270 2292.600 ;
        RECT 463.650 2079.740 504.270 2276.820 ;
        RECT 463.650 1766.820 464.550 2079.740 ;
        RECT 466.950 2065.560 504.270 2079.740 ;
        RECT 506.670 2065.560 507.950 2292.600 ;
        RECT 510.350 2065.560 531.250 2292.600 ;
        RECT 466.950 2035.860 531.250 2065.560 ;
        RECT 533.650 2035.860 534.550 2329.740 ;
        RECT 466.950 2008.925 534.550 2035.860 ;
        RECT 536.950 2274.365 601.250 2334.235 ;
        RECT 603.650 2274.365 604.550 2334.235 ;
        RECT 606.950 2274.365 671.250 2334.235 ;
        RECT 673.650 2274.365 674.550 2334.235 ;
        RECT 536.950 2080.835 674.550 2274.365 ;
        RECT 536.950 2008.925 601.250 2080.835 ;
        RECT 603.650 2008.925 604.550 2080.835 ;
        RECT 606.950 2008.925 671.250 2080.835 ;
        RECT 673.650 2008.925 674.550 2080.835 ;
        RECT 676.950 2008.925 741.250 2334.235 ;
        RECT 466.950 1824.235 741.250 2008.925 ;
        RECT 466.950 1819.740 534.550 1824.235 ;
        RECT 466.950 1783.960 531.250 1819.740 ;
        RECT 466.950 1766.820 504.270 1783.960 ;
        RECT 463.650 1569.740 504.270 1766.820 ;
        RECT 463.650 1256.820 464.550 1569.740 ;
        RECT 466.950 1554.200 504.270 1569.740 ;
        RECT 506.670 1554.200 507.950 1783.960 ;
        RECT 510.350 1554.200 531.250 1783.960 ;
        RECT 466.950 1525.860 531.250 1554.200 ;
        RECT 533.650 1525.860 534.550 1819.740 ;
        RECT 466.950 1498.925 534.550 1525.860 ;
        RECT 536.950 1498.925 601.250 1824.235 ;
        RECT 603.650 1498.925 604.550 1824.235 ;
        RECT 606.950 1498.925 671.250 1824.235 ;
        RECT 673.650 1498.925 674.550 1824.235 ;
        RECT 676.950 1498.925 741.250 1824.235 ;
        RECT 466.950 1314.235 741.250 1498.925 ;
        RECT 466.950 1309.740 534.550 1314.235 ;
        RECT 466.950 1272.600 531.250 1309.740 ;
        RECT 466.950 1256.820 511.630 1272.600 ;
        RECT 463.650 1059.740 511.630 1256.820 ;
        RECT 463.650 746.820 464.550 1059.740 ;
        RECT 466.950 1045.560 511.630 1059.740 ;
        RECT 514.030 1045.560 515.310 1272.600 ;
        RECT 517.710 1045.560 531.250 1272.600 ;
        RECT 466.950 1015.860 531.250 1045.560 ;
        RECT 533.650 1015.860 534.550 1309.740 ;
        RECT 466.950 988.925 534.550 1015.860 ;
        RECT 536.950 988.925 601.250 1314.235 ;
        RECT 603.650 988.925 604.550 1314.235 ;
        RECT 606.950 1124.485 671.250 1314.235 ;
        RECT 673.650 1124.485 674.550 1314.235 ;
        RECT 606.950 1064.915 674.550 1124.485 ;
        RECT 606.950 988.925 671.250 1064.915 ;
        RECT 673.650 988.925 674.550 1064.915 ;
        RECT 676.950 988.925 741.250 1314.235 ;
        RECT 466.950 804.235 741.250 988.925 ;
        RECT 466.950 799.740 534.550 804.235 ;
        RECT 466.950 763.960 531.250 799.740 ;
        RECT 466.950 746.820 504.270 763.960 ;
        RECT 463.650 549.740 504.270 746.820 ;
        RECT 463.650 9.240 464.550 549.740 ;
        RECT 466.950 534.200 504.270 549.740 ;
        RECT 506.670 534.200 507.950 763.960 ;
        RECT 510.350 534.200 531.250 763.960 ;
        RECT 466.950 9.240 531.250 534.200 ;
        RECT 533.650 9.240 534.550 799.740 ;
        RECT 536.950 9.240 601.250 804.235 ;
        RECT 603.650 9.240 604.550 804.235 ;
        RECT 606.950 9.240 671.250 804.235 ;
        RECT 673.650 9.240 674.550 804.235 ;
        RECT 676.950 9.240 741.250 804.235 ;
        RECT 743.650 9.240 744.550 2935.745 ;
        RECT 746.950 2244.245 811.250 2935.745 ;
        RECT 813.650 2244.245 814.550 2935.745 ;
        RECT 816.950 2244.245 881.250 2935.745 ;
        RECT 883.650 2244.245 884.550 2935.745 ;
        RECT 886.950 2244.245 951.250 2935.745 ;
        RECT 746.950 2092.195 951.250 2244.245 ;
        RECT 746.950 1751.925 811.250 2092.195 ;
        RECT 813.650 1751.925 814.550 2092.195 ;
        RECT 816.950 1751.925 881.250 2092.195 ;
        RECT 883.650 1751.925 884.550 2092.195 ;
        RECT 886.950 1751.925 951.250 2092.195 ;
        RECT 953.650 2526.820 954.550 2935.745 ;
        RECT 956.950 2542.840 1021.250 2935.745 ;
        RECT 956.950 2526.820 997.390 2542.840 ;
        RECT 953.650 2329.740 997.390 2526.820 ;
        RECT 953.650 2286.820 954.550 2329.740 ;
        RECT 956.950 2313.080 997.390 2329.740 ;
        RECT 999.790 2313.080 1001.070 2542.840 ;
        RECT 1003.470 2518.925 1021.250 2542.840 ;
        RECT 1023.650 2518.925 1024.550 2935.745 ;
        RECT 1026.950 2518.925 1091.250 2935.745 ;
        RECT 1093.650 2518.925 1094.550 2935.745 ;
        RECT 1096.950 2518.925 1161.250 2935.745 ;
        RECT 1163.650 2518.925 1164.550 2935.745 ;
        RECT 1166.950 2518.925 1231.250 2935.745 ;
        RECT 1003.470 2334.235 1231.250 2518.925 ;
        RECT 1003.470 2313.080 1021.250 2334.235 ;
        RECT 956.950 2289.880 1021.250 2313.080 ;
        RECT 956.950 2286.820 1006.590 2289.880 ;
        RECT 953.650 2089.740 1006.590 2286.820 ;
        RECT 953.650 2016.820 954.550 2089.740 ;
        RECT 956.950 2076.440 1006.590 2089.740 ;
        RECT 1008.990 2076.440 1021.250 2289.880 ;
        RECT 956.950 2034.200 1021.250 2076.440 ;
        RECT 956.950 2016.820 997.390 2034.200 ;
        RECT 953.650 1819.740 997.390 2016.820 ;
        RECT 953.650 1776.820 954.550 1819.740 ;
        RECT 956.950 1804.440 997.390 1819.740 ;
        RECT 999.790 1804.440 1001.070 2034.200 ;
        RECT 1003.470 2008.925 1021.250 2034.200 ;
        RECT 1023.650 2008.925 1024.550 2334.235 ;
        RECT 1026.950 2008.925 1091.250 2334.235 ;
        RECT 1093.650 2008.925 1094.550 2334.235 ;
        RECT 1096.950 2274.365 1161.250 2334.235 ;
        RECT 1163.650 2274.365 1164.550 2334.235 ;
        RECT 1166.950 2274.365 1231.250 2334.235 ;
        RECT 1096.950 2080.835 1231.250 2274.365 ;
        RECT 1096.950 2008.925 1161.250 2080.835 ;
        RECT 1163.650 2008.925 1164.550 2080.835 ;
        RECT 1166.950 2008.925 1231.250 2080.835 ;
        RECT 1003.470 1824.235 1231.250 2008.925 ;
        RECT 1003.470 1804.440 1021.250 1824.235 ;
        RECT 956.950 1783.960 1021.250 1804.440 ;
        RECT 956.950 1776.820 1006.590 1783.960 ;
        RECT 953.650 1751.925 1006.590 1776.820 ;
        RECT 746.950 1580.835 1006.590 1751.925 ;
        RECT 746.950 1241.925 811.250 1580.835 ;
        RECT 813.650 1241.925 814.550 1580.835 ;
        RECT 816.950 1241.925 881.250 1580.835 ;
        RECT 883.650 1241.925 884.550 1580.835 ;
        RECT 886.950 1241.925 951.250 1580.835 ;
        RECT 953.650 1579.740 1006.590 1580.835 ;
        RECT 953.650 1506.820 954.550 1579.740 ;
        RECT 956.950 1565.080 1006.590 1579.740 ;
        RECT 1008.990 1565.080 1021.250 1783.960 ;
        RECT 956.950 1522.840 1021.250 1565.080 ;
        RECT 956.950 1506.820 997.390 1522.840 ;
        RECT 953.650 1309.740 997.390 1506.820 ;
        RECT 953.650 1266.820 954.550 1309.740 ;
        RECT 956.950 1293.080 997.390 1309.740 ;
        RECT 999.790 1293.080 1001.070 1522.840 ;
        RECT 1003.470 1498.925 1021.250 1522.840 ;
        RECT 1023.650 1498.925 1024.550 1824.235 ;
        RECT 1026.950 1498.925 1091.250 1824.235 ;
        RECT 1093.650 1498.925 1094.550 1824.235 ;
        RECT 1096.950 1634.485 1161.250 1824.235 ;
        RECT 1163.650 1634.485 1164.550 1824.235 ;
        RECT 1166.950 1634.485 1231.250 1824.235 ;
        RECT 1096.950 1574.915 1231.250 1634.485 ;
        RECT 1096.950 1498.925 1161.250 1574.915 ;
        RECT 1163.650 1498.925 1164.550 1574.915 ;
        RECT 1166.950 1498.925 1231.250 1574.915 ;
        RECT 1003.470 1314.235 1231.250 1498.925 ;
        RECT 1003.470 1293.080 1021.250 1314.235 ;
        RECT 956.950 1272.600 1021.250 1293.080 ;
        RECT 956.950 1266.820 1006.590 1272.600 ;
        RECT 953.650 1241.925 1006.590 1266.820 ;
        RECT 746.950 1070.835 1006.590 1241.925 ;
        RECT 746.950 731.925 811.250 1070.835 ;
        RECT 813.650 731.925 814.550 1070.835 ;
        RECT 816.950 731.925 881.250 1070.835 ;
        RECT 883.650 731.925 884.550 1070.835 ;
        RECT 886.950 731.925 951.250 1070.835 ;
        RECT 953.650 1069.740 1006.590 1070.835 ;
        RECT 953.650 996.820 954.550 1069.740 ;
        RECT 956.950 1053.720 1006.590 1069.740 ;
        RECT 1008.990 1053.720 1021.250 1272.600 ;
        RECT 956.950 1014.200 1021.250 1053.720 ;
        RECT 956.950 996.820 997.390 1014.200 ;
        RECT 953.650 799.740 997.390 996.820 ;
        RECT 953.650 756.820 954.550 799.740 ;
        RECT 956.950 784.440 997.390 799.740 ;
        RECT 999.790 784.440 1001.070 1014.200 ;
        RECT 1003.470 988.925 1021.250 1014.200 ;
        RECT 1023.650 988.925 1024.550 1314.235 ;
        RECT 1026.950 988.925 1091.250 1314.235 ;
        RECT 1093.650 988.925 1094.550 1314.235 ;
        RECT 1096.950 1124.485 1161.250 1314.235 ;
        RECT 1163.650 1124.485 1164.550 1314.235 ;
        RECT 1166.950 1124.485 1231.250 1314.235 ;
        RECT 1096.950 1064.915 1231.250 1124.485 ;
        RECT 1096.950 988.925 1161.250 1064.915 ;
        RECT 1163.650 988.925 1164.550 1064.915 ;
        RECT 1166.950 988.925 1231.250 1064.915 ;
        RECT 1003.470 804.235 1231.250 988.925 ;
        RECT 1003.470 784.440 1021.250 804.235 ;
        RECT 956.950 761.240 1021.250 784.440 ;
        RECT 956.950 756.820 1006.590 761.240 ;
        RECT 953.650 731.925 1006.590 756.820 ;
        RECT 746.950 560.835 1006.590 731.925 ;
        RECT 746.950 482.125 811.250 560.835 ;
        RECT 813.650 482.125 814.550 560.835 ;
        RECT 816.950 482.125 881.250 560.835 ;
        RECT 883.650 482.125 884.550 560.835 ;
        RECT 886.950 482.125 951.250 560.835 ;
        RECT 746.950 336.195 951.250 482.125 ;
        RECT 746.950 9.240 811.250 336.195 ;
        RECT 813.650 9.240 814.550 336.195 ;
        RECT 816.950 9.240 881.250 336.195 ;
        RECT 883.650 9.240 884.550 336.195 ;
        RECT 886.950 9.240 951.250 336.195 ;
        RECT 953.650 559.740 1006.590 560.835 ;
        RECT 953.650 496.820 954.550 559.740 ;
        RECT 956.950 547.800 1006.590 559.740 ;
        RECT 1008.990 547.800 1021.250 761.240 ;
        RECT 956.950 496.820 1021.250 547.800 ;
        RECT 953.650 494.680 1021.250 496.820 ;
        RECT 953.650 299.740 1006.590 494.680 ;
        RECT 953.650 9.240 954.550 299.740 ;
        RECT 956.950 286.680 1006.590 299.740 ;
        RECT 1008.990 286.680 1021.250 494.680 ;
        RECT 956.950 9.240 1021.250 286.680 ;
        RECT 1023.650 9.240 1024.550 804.235 ;
        RECT 1026.950 9.240 1091.250 804.235 ;
        RECT 1093.650 9.240 1094.550 804.235 ;
        RECT 1096.950 614.485 1161.250 804.235 ;
        RECT 1163.650 614.485 1164.550 804.235 ;
        RECT 1166.950 614.485 1231.250 804.235 ;
        RECT 1096.950 554.915 1231.250 614.485 ;
        RECT 1096.950 377.125 1161.250 554.915 ;
        RECT 1163.650 377.125 1164.550 554.915 ;
        RECT 1096.950 281.515 1164.550 377.125 ;
        RECT 1096.950 9.240 1161.250 281.515 ;
        RECT 1163.650 9.240 1164.550 281.515 ;
        RECT 1166.950 9.240 1231.250 554.915 ;
        RECT 1233.650 9.240 1234.550 2935.745 ;
        RECT 1236.950 2542.840 1301.250 2935.745 ;
        RECT 1236.950 2313.080 1262.350 2542.840 ;
        RECT 1264.750 2313.080 1266.030 2542.840 ;
        RECT 1268.430 2313.080 1301.250 2542.840 ;
        RECT 1236.950 2292.600 1301.250 2313.080 ;
        RECT 1236.950 2073.720 1255.910 2292.600 ;
        RECT 1258.310 2244.245 1301.250 2292.600 ;
        RECT 1303.650 2244.245 1304.550 2935.745 ;
        RECT 1306.950 2244.245 1371.250 2935.745 ;
        RECT 1373.650 2244.245 1374.550 2935.745 ;
        RECT 1376.950 2244.245 1441.250 2935.745 ;
        RECT 1258.310 2092.195 1441.250 2244.245 ;
        RECT 1258.310 2073.720 1301.250 2092.195 ;
        RECT 1236.950 2034.200 1301.250 2073.720 ;
        RECT 1236.950 1804.440 1262.350 2034.200 ;
        RECT 1264.750 1804.440 1266.030 2034.200 ;
        RECT 1268.430 1804.440 1301.250 2034.200 ;
        RECT 1236.950 1781.240 1301.250 1804.440 ;
        RECT 1236.950 1567.800 1255.910 1781.240 ;
        RECT 1258.310 1751.925 1301.250 1781.240 ;
        RECT 1303.650 1751.925 1304.550 2092.195 ;
        RECT 1306.950 1751.925 1371.250 2092.195 ;
        RECT 1373.650 1751.925 1374.550 2092.195 ;
        RECT 1376.950 1751.925 1441.250 2092.195 ;
        RECT 1443.650 1751.925 1444.550 2935.745 ;
        RECT 1446.950 1751.925 1511.250 2935.745 ;
        RECT 1258.310 1580.835 1511.250 1751.925 ;
        RECT 1258.310 1567.800 1301.250 1580.835 ;
        RECT 1236.950 1522.840 1301.250 1567.800 ;
        RECT 1236.950 1293.080 1262.350 1522.840 ;
        RECT 1264.750 1293.080 1266.030 1522.840 ;
        RECT 1268.430 1293.080 1301.250 1522.840 ;
        RECT 1236.950 1269.880 1301.250 1293.080 ;
        RECT 1236.950 1056.440 1255.910 1269.880 ;
        RECT 1258.310 1241.925 1301.250 1269.880 ;
        RECT 1303.650 1241.925 1304.550 1580.835 ;
        RECT 1306.950 1241.925 1371.250 1580.835 ;
        RECT 1373.650 1241.925 1374.550 1580.835 ;
        RECT 1376.950 1241.925 1441.250 1580.835 ;
        RECT 1443.650 1241.925 1444.550 1580.835 ;
        RECT 1446.950 1241.925 1511.250 1580.835 ;
        RECT 1258.310 1070.835 1511.250 1241.925 ;
        RECT 1258.310 1056.440 1301.250 1070.835 ;
        RECT 1236.950 1014.200 1301.250 1056.440 ;
        RECT 1236.950 784.440 1262.350 1014.200 ;
        RECT 1264.750 784.440 1266.030 1014.200 ;
        RECT 1268.430 784.440 1301.250 1014.200 ;
        RECT 1236.950 763.960 1301.250 784.440 ;
        RECT 1236.950 545.080 1255.910 763.960 ;
        RECT 1258.310 731.925 1301.250 763.960 ;
        RECT 1303.650 731.925 1304.550 1070.835 ;
        RECT 1306.950 731.925 1371.250 1070.835 ;
        RECT 1373.650 731.925 1374.550 1070.835 ;
        RECT 1376.950 731.925 1441.250 1070.835 ;
        RECT 1443.650 731.925 1444.550 1070.835 ;
        RECT 1446.950 731.925 1511.250 1070.835 ;
        RECT 1258.310 560.835 1511.250 731.925 ;
        RECT 1258.310 545.080 1301.250 560.835 ;
        RECT 1236.950 494.680 1301.250 545.080 ;
        RECT 1236.950 283.960 1259.590 494.680 ;
        RECT 1261.990 283.960 1263.270 494.680 ;
        RECT 1265.670 482.125 1301.250 494.680 ;
        RECT 1303.650 482.125 1304.550 560.835 ;
        RECT 1306.950 482.125 1371.250 560.835 ;
        RECT 1373.650 482.125 1374.550 560.835 ;
        RECT 1376.950 482.125 1441.250 560.835 ;
        RECT 1265.670 336.195 1441.250 482.125 ;
        RECT 1265.670 283.960 1301.250 336.195 ;
        RECT 1236.950 9.240 1301.250 283.960 ;
        RECT 1303.650 9.240 1304.550 336.195 ;
        RECT 1306.950 9.240 1371.250 336.195 ;
        RECT 1373.650 9.240 1374.550 336.195 ;
        RECT 1376.950 9.240 1441.250 336.195 ;
        RECT 1443.650 9.240 1444.550 560.835 ;
        RECT 1446.950 9.240 1511.250 560.835 ;
        RECT 1513.650 9.240 1514.550 2935.745 ;
        RECT 1516.950 2518.925 1581.250 2935.745 ;
        RECT 1583.650 2806.820 1584.550 2935.745 ;
        RECT 1586.950 2806.820 1651.250 2935.745 ;
        RECT 1583.650 2609.740 1651.250 2806.820 ;
        RECT 1583.650 2518.925 1584.550 2609.740 ;
        RECT 1586.950 2518.925 1651.250 2609.740 ;
        RECT 1653.650 2518.925 1654.550 2935.745 ;
        RECT 1656.950 2518.925 1721.250 2935.745 ;
        RECT 1723.650 2518.925 1724.550 2935.745 ;
        RECT 1726.950 2542.840 1791.250 2935.745 ;
        RECT 1726.950 2518.925 1772.030 2542.840 ;
        RECT 1516.950 2334.235 1772.030 2518.925 ;
        RECT 1516.950 2008.925 1581.250 2334.235 ;
        RECT 1583.650 2008.925 1584.550 2334.235 ;
        RECT 1586.950 2274.365 1651.250 2334.235 ;
        RECT 1653.650 2274.365 1654.550 2334.235 ;
        RECT 1656.950 2274.365 1721.250 2334.235 ;
        RECT 1586.950 2080.835 1721.250 2274.365 ;
        RECT 1586.950 2008.925 1651.250 2080.835 ;
        RECT 1653.650 2008.925 1654.550 2080.835 ;
        RECT 1656.950 2008.925 1721.250 2080.835 ;
        RECT 1723.650 2008.925 1724.550 2334.235 ;
        RECT 1726.950 2313.080 1772.030 2334.235 ;
        RECT 1774.430 2313.080 1775.710 2542.840 ;
        RECT 1778.110 2313.080 1791.250 2542.840 ;
        RECT 1726.950 2292.600 1791.250 2313.080 ;
        RECT 1726.950 2073.720 1764.670 2292.600 ;
        RECT 1767.070 2073.720 1768.350 2292.600 ;
        RECT 1770.750 2073.720 1791.250 2292.600 ;
        RECT 1726.950 2034.200 1791.250 2073.720 ;
        RECT 1726.950 2008.925 1772.030 2034.200 ;
        RECT 1516.950 1824.235 1772.030 2008.925 ;
        RECT 1516.950 1498.925 1581.250 1824.235 ;
        RECT 1583.650 1498.925 1584.550 1824.235 ;
        RECT 1586.950 1498.925 1651.250 1824.235 ;
        RECT 1653.650 1498.925 1654.550 1824.235 ;
        RECT 1656.950 1498.925 1721.250 1824.235 ;
        RECT 1723.650 1498.925 1724.550 1824.235 ;
        RECT 1726.950 1804.440 1772.030 1824.235 ;
        RECT 1774.430 1804.440 1775.710 2034.200 ;
        RECT 1778.110 1804.440 1791.250 2034.200 ;
        RECT 1726.950 1783.960 1791.250 1804.440 ;
        RECT 1726.950 1565.080 1764.670 1783.960 ;
        RECT 1767.070 1565.080 1768.350 1783.960 ;
        RECT 1770.750 1565.080 1791.250 1783.960 ;
        RECT 1726.950 1522.840 1791.250 1565.080 ;
        RECT 1726.950 1498.925 1772.030 1522.840 ;
        RECT 1516.950 1314.235 1772.030 1498.925 ;
        RECT 1516.950 988.925 1581.250 1314.235 ;
        RECT 1583.650 988.925 1584.550 1314.235 ;
        RECT 1586.950 988.925 1651.250 1314.235 ;
        RECT 1653.650 988.925 1654.550 1314.235 ;
        RECT 1656.950 988.925 1721.250 1314.235 ;
        RECT 1723.650 988.925 1724.550 1314.235 ;
        RECT 1726.950 1293.080 1772.030 1314.235 ;
        RECT 1774.430 1293.080 1775.710 1522.840 ;
        RECT 1778.110 1293.080 1791.250 1522.840 ;
        RECT 1726.950 1272.600 1791.250 1293.080 ;
        RECT 1726.950 1053.720 1764.670 1272.600 ;
        RECT 1767.070 1053.720 1768.350 1272.600 ;
        RECT 1770.750 1053.720 1791.250 1272.600 ;
        RECT 1726.950 1014.200 1791.250 1053.720 ;
        RECT 1726.950 988.925 1772.030 1014.200 ;
        RECT 1516.950 804.235 1772.030 988.925 ;
        RECT 1516.950 9.240 1581.250 804.235 ;
        RECT 1583.650 226.820 1584.550 804.235 ;
        RECT 1586.950 377.125 1651.250 804.235 ;
        RECT 1653.650 377.125 1654.550 804.235 ;
        RECT 1656.950 377.125 1721.250 804.235 ;
        RECT 1586.950 281.515 1721.250 377.125 ;
        RECT 1586.950 226.820 1651.250 281.515 ;
        RECT 1583.650 29.740 1651.250 226.820 ;
        RECT 1583.650 9.240 1584.550 29.740 ;
        RECT 1586.950 9.240 1651.250 29.740 ;
        RECT 1653.650 9.240 1654.550 281.515 ;
        RECT 1656.950 9.240 1721.250 281.515 ;
        RECT 1723.650 9.240 1724.550 804.235 ;
        RECT 1726.950 784.440 1772.030 804.235 ;
        RECT 1774.430 784.440 1775.710 1014.200 ;
        RECT 1778.110 784.440 1791.250 1014.200 ;
        RECT 1726.950 774.840 1791.250 784.440 ;
        RECT 1726.950 545.080 1764.670 774.840 ;
        RECT 1767.070 545.080 1768.350 774.840 ;
        RECT 1770.750 545.080 1791.250 774.840 ;
        RECT 1726.950 494.680 1791.250 545.080 ;
        RECT 1726.950 283.960 1769.270 494.680 ;
        RECT 1771.670 283.960 1772.950 494.680 ;
        RECT 1775.350 283.960 1791.250 494.680 ;
        RECT 1726.950 9.240 1791.250 283.960 ;
        RECT 1793.650 2244.245 1794.550 2935.745 ;
        RECT 1796.950 2244.245 1861.250 2935.745 ;
        RECT 1863.650 2244.245 1864.550 2935.745 ;
        RECT 1866.950 2457.045 1931.250 2935.745 ;
        RECT 1933.650 2457.045 1934.550 2935.745 ;
        RECT 1936.950 2457.045 2001.250 2935.745 ;
        RECT 1866.950 2356.675 2001.250 2457.045 ;
        RECT 1866.950 2244.245 1931.250 2356.675 ;
        RECT 1793.650 2092.195 1931.250 2244.245 ;
        RECT 1793.650 9.240 1794.550 2092.195 ;
        RECT 1796.950 1751.925 1861.250 2092.195 ;
        RECT 1863.650 1751.925 1864.550 2092.195 ;
        RECT 1866.950 1947.045 1931.250 2092.195 ;
        RECT 1933.650 1947.045 1934.550 2356.675 ;
        RECT 1936.950 1947.045 2001.250 2356.675 ;
        RECT 1866.950 1846.675 2001.250 1947.045 ;
        RECT 1866.950 1751.925 1931.250 1846.675 ;
        RECT 1933.650 1751.925 1934.550 1846.675 ;
        RECT 1936.950 1751.925 2001.250 1846.675 ;
        RECT 1796.950 1580.835 2001.250 1751.925 ;
        RECT 1796.950 1241.925 1861.250 1580.835 ;
        RECT 1863.650 1241.925 1864.550 1580.835 ;
        RECT 1866.950 1437.045 1931.250 1580.835 ;
        RECT 1933.650 1437.045 1934.550 1580.835 ;
        RECT 1936.950 1437.045 2001.250 1580.835 ;
        RECT 1866.950 1336.675 2001.250 1437.045 ;
        RECT 1866.950 1241.925 1931.250 1336.675 ;
        RECT 1933.650 1241.925 1934.550 1336.675 ;
        RECT 1936.950 1241.925 2001.250 1336.675 ;
        RECT 1796.950 1070.835 2001.250 1241.925 ;
        RECT 1796.950 731.925 1861.250 1070.835 ;
        RECT 1863.650 731.925 1864.550 1070.835 ;
        RECT 1866.950 927.045 1931.250 1070.835 ;
        RECT 1933.650 927.045 1934.550 1070.835 ;
        RECT 1936.950 927.045 2001.250 1070.835 ;
        RECT 1866.950 826.675 2001.250 927.045 ;
        RECT 1866.950 731.925 1931.250 826.675 ;
        RECT 1933.650 731.925 1934.550 826.675 ;
        RECT 1936.950 731.925 2001.250 826.675 ;
        RECT 1796.950 560.835 2001.250 731.925 ;
        RECT 1796.950 482.125 1861.250 560.835 ;
        RECT 1863.650 482.125 1864.550 560.835 ;
        RECT 1866.950 482.125 1931.250 560.835 ;
        RECT 1933.650 482.125 1934.550 560.835 ;
        RECT 1936.950 482.125 2001.250 560.835 ;
        RECT 1796.950 336.195 2001.250 482.125 ;
        RECT 1796.950 9.240 1861.250 336.195 ;
        RECT 1863.650 9.240 1864.550 336.195 ;
        RECT 1866.950 9.240 1931.250 336.195 ;
        RECT 1933.650 9.240 1934.550 336.195 ;
        RECT 1936.950 9.240 2001.250 336.195 ;
        RECT 2003.650 9.240 2004.550 2935.745 ;
        RECT 2006.950 2542.840 2071.250 2935.745 ;
        RECT 2006.950 2313.080 2016.750 2542.840 ;
        RECT 2019.150 2313.080 2020.430 2542.840 ;
        RECT 2022.830 2518.925 2071.250 2542.840 ;
        RECT 2073.650 2518.925 2074.550 2935.745 ;
        RECT 2076.950 2518.925 2141.250 2935.745 ;
        RECT 2143.650 2518.925 2144.550 2935.745 ;
        RECT 2146.950 2518.925 2211.250 2935.745 ;
        RECT 2213.650 2545.860 2214.550 2935.745 ;
        RECT 2216.950 2545.860 2281.250 2935.745 ;
        RECT 2213.650 2518.925 2281.250 2545.860 ;
        RECT 2022.830 2334.235 2281.250 2518.925 ;
        RECT 2022.830 2313.080 2071.250 2334.235 ;
        RECT 2006.950 2292.600 2071.250 2313.080 ;
        RECT 2006.950 2073.720 2024.110 2292.600 ;
        RECT 2026.510 2073.720 2027.790 2292.600 ;
        RECT 2030.190 2073.720 2071.250 2292.600 ;
        RECT 2006.950 2034.200 2071.250 2073.720 ;
        RECT 2006.950 1804.440 2016.750 2034.200 ;
        RECT 2019.150 1804.440 2020.430 2034.200 ;
        RECT 2022.830 2008.925 2071.250 2034.200 ;
        RECT 2073.650 2276.820 2074.550 2334.235 ;
        RECT 2076.950 2276.820 2141.250 2334.235 ;
        RECT 2073.650 2274.365 2141.250 2276.820 ;
        RECT 2143.650 2274.365 2144.550 2334.235 ;
        RECT 2146.950 2274.365 2211.250 2334.235 ;
        RECT 2073.650 2080.835 2211.250 2274.365 ;
        RECT 2073.650 2079.740 2141.250 2080.835 ;
        RECT 2073.650 2008.925 2074.550 2079.740 ;
        RECT 2076.950 2008.925 2141.250 2079.740 ;
        RECT 2143.650 2008.925 2144.550 2080.835 ;
        RECT 2146.950 2008.925 2211.250 2080.835 ;
        RECT 2213.650 2329.740 2281.250 2334.235 ;
        RECT 2213.650 2035.860 2214.550 2329.740 ;
        RECT 2216.950 2035.860 2281.250 2329.740 ;
        RECT 2213.650 2008.925 2281.250 2035.860 ;
        RECT 2022.830 1824.235 2281.250 2008.925 ;
        RECT 2022.830 1804.440 2071.250 1824.235 ;
        RECT 2006.950 1783.960 2071.250 1804.440 ;
        RECT 2006.950 1565.080 2024.110 1783.960 ;
        RECT 2026.510 1565.080 2027.790 1783.960 ;
        RECT 2030.190 1565.080 2071.250 1783.960 ;
        RECT 2006.950 1522.840 2071.250 1565.080 ;
        RECT 2006.950 1293.080 2016.750 1522.840 ;
        RECT 2019.150 1293.080 2020.430 1522.840 ;
        RECT 2022.830 1498.925 2071.250 1522.840 ;
        RECT 2073.650 1766.820 2074.550 1824.235 ;
        RECT 2076.950 1766.820 2141.250 1824.235 ;
        RECT 2073.650 1569.740 2141.250 1766.820 ;
        RECT 2073.650 1498.925 2074.550 1569.740 ;
        RECT 2076.950 1498.925 2141.250 1569.740 ;
        RECT 2143.650 1498.925 2144.550 1824.235 ;
        RECT 2146.950 1498.925 2211.250 1824.235 ;
        RECT 2213.650 1819.740 2281.250 1824.235 ;
        RECT 2213.650 1525.860 2214.550 1819.740 ;
        RECT 2216.950 1525.860 2281.250 1819.740 ;
        RECT 2213.650 1498.925 2281.250 1525.860 ;
        RECT 2022.830 1314.235 2281.250 1498.925 ;
        RECT 2022.830 1293.080 2071.250 1314.235 ;
        RECT 2006.950 1278.040 2071.250 1293.080 ;
        RECT 2006.950 1053.720 2024.110 1278.040 ;
        RECT 2026.510 1053.720 2027.790 1278.040 ;
        RECT 2030.190 1053.720 2071.250 1278.040 ;
        RECT 2006.950 1014.200 2071.250 1053.720 ;
        RECT 2006.950 784.440 2016.750 1014.200 ;
        RECT 2019.150 784.440 2020.430 1014.200 ;
        RECT 2022.830 988.925 2071.250 1014.200 ;
        RECT 2073.650 1259.820 2074.550 1314.235 ;
        RECT 2076.950 1259.820 2141.250 1314.235 ;
        RECT 2073.650 1062.740 2141.250 1259.820 ;
        RECT 2073.650 988.925 2074.550 1062.740 ;
        RECT 2076.950 988.925 2141.250 1062.740 ;
        RECT 2143.650 988.925 2144.550 1314.235 ;
        RECT 2146.950 988.925 2211.250 1314.235 ;
        RECT 2213.650 1309.740 2281.250 1314.235 ;
        RECT 2213.650 1015.860 2214.550 1309.740 ;
        RECT 2216.950 1015.860 2281.250 1309.740 ;
        RECT 2213.650 988.925 2281.250 1015.860 ;
        RECT 2022.830 804.235 2281.250 988.925 ;
        RECT 2022.830 784.440 2071.250 804.235 ;
        RECT 2006.950 763.960 2071.250 784.440 ;
        RECT 2006.950 545.080 2024.110 763.960 ;
        RECT 2026.510 545.080 2027.790 763.960 ;
        RECT 2030.190 545.080 2071.250 763.960 ;
        RECT 2006.950 494.680 2071.250 545.080 ;
        RECT 2006.950 283.960 2024.110 494.680 ;
        RECT 2026.510 283.960 2027.790 494.680 ;
        RECT 2030.190 283.960 2071.250 494.680 ;
        RECT 2006.950 9.240 2071.250 283.960 ;
        RECT 2073.650 746.820 2074.550 804.235 ;
        RECT 2076.950 746.820 2141.250 804.235 ;
        RECT 2073.650 549.740 2141.250 746.820 ;
        RECT 2073.650 476.820 2074.550 549.740 ;
        RECT 2076.950 476.820 2141.250 549.740 ;
        RECT 2073.650 377.125 2141.250 476.820 ;
        RECT 2143.650 377.125 2144.550 804.235 ;
        RECT 2146.950 377.125 2211.250 804.235 ;
        RECT 2073.650 281.515 2211.250 377.125 ;
        RECT 2073.650 279.740 2141.250 281.515 ;
        RECT 2073.650 9.240 2074.550 279.740 ;
        RECT 2076.950 9.240 2141.250 279.740 ;
        RECT 2143.650 9.240 2144.550 281.515 ;
        RECT 2146.950 9.240 2211.250 281.515 ;
        RECT 2213.650 799.740 2281.250 804.235 ;
        RECT 2213.650 9.240 2214.550 799.740 ;
        RECT 2216.950 9.240 2281.250 799.740 ;
        RECT 2283.650 9.240 2284.550 2935.745 ;
        RECT 2286.950 2398.245 2351.250 2935.745 ;
        RECT 2353.650 2398.245 2354.550 2935.745 ;
        RECT 2356.950 2398.245 2421.250 2935.745 ;
        RECT 2286.950 2304.675 2421.250 2398.245 ;
        RECT 2286.950 1888.245 2351.250 2304.675 ;
        RECT 2353.650 1888.245 2354.550 2304.675 ;
        RECT 2356.950 2175.885 2421.250 2304.675 ;
        RECT 2423.650 2187.860 2424.550 2935.745 ;
        RECT 2426.950 2187.860 2491.250 2935.745 ;
        RECT 2423.650 2175.885 2491.250 2187.860 ;
        RECT 2356.950 2044.235 2491.250 2175.885 ;
        RECT 2356.950 1888.245 2421.250 2044.235 ;
        RECT 2286.950 1794.675 2421.250 1888.245 ;
        RECT 2286.950 1718.925 2351.250 1794.675 ;
        RECT 2353.650 1718.925 2354.550 1794.675 ;
        RECT 2356.950 1718.925 2421.250 1794.675 ;
        RECT 2423.650 2039.740 2491.250 2044.235 ;
        RECT 2423.650 1718.925 2424.550 2039.740 ;
        RECT 2426.950 1718.925 2491.250 2039.740 ;
        RECT 2286.950 1532.195 2491.250 1718.925 ;
        RECT 2286.950 1378.245 2351.250 1532.195 ;
        RECT 2353.650 1378.245 2354.550 1532.195 ;
        RECT 2356.950 1378.245 2421.250 1532.195 ;
        RECT 2286.950 1284.675 2421.250 1378.245 ;
        RECT 2286.950 1208.925 2351.250 1284.675 ;
        RECT 2353.650 1208.925 2354.550 1284.675 ;
        RECT 2356.950 1208.925 2421.250 1284.675 ;
        RECT 2423.650 1208.925 2424.550 1532.195 ;
        RECT 2426.950 1208.925 2491.250 1532.195 ;
        RECT 2286.950 1022.195 2491.250 1208.925 ;
        RECT 2286.950 868.245 2351.250 1022.195 ;
        RECT 2353.650 868.245 2354.550 1022.195 ;
        RECT 2356.950 868.245 2421.250 1022.195 ;
        RECT 2286.950 774.675 2421.250 868.245 ;
        RECT 2286.950 728.925 2351.250 774.675 ;
        RECT 2353.650 728.925 2354.550 774.675 ;
        RECT 2356.950 728.925 2421.250 774.675 ;
        RECT 2423.650 728.925 2424.550 1022.195 ;
        RECT 2426.950 728.925 2491.250 1022.195 ;
        RECT 2286.950 542.195 2491.250 728.925 ;
        RECT 2286.950 492.325 2351.250 542.195 ;
        RECT 2353.650 492.325 2354.550 542.195 ;
        RECT 2356.950 492.325 2421.250 542.195 ;
        RECT 2423.650 492.325 2424.550 542.195 ;
        RECT 2426.950 492.325 2491.250 542.195 ;
        RECT 2286.950 308.995 2491.250 492.325 ;
        RECT 2286.950 9.240 2351.250 308.995 ;
        RECT 2353.650 9.240 2354.550 308.995 ;
        RECT 2356.950 9.240 2421.250 308.995 ;
        RECT 2423.650 9.240 2424.550 308.995 ;
        RECT 2426.950 9.240 2491.250 308.995 ;
        RECT 2493.650 2187.860 2494.550 2935.745 ;
        RECT 2496.950 2507.480 2561.250 2935.745 ;
        RECT 2496.950 2294.040 2531.950 2507.480 ;
        RECT 2534.350 2294.040 2535.630 2507.480 ;
        RECT 2538.030 2294.040 2561.250 2507.480 ;
        RECT 2496.950 2187.860 2561.250 2294.040 ;
        RECT 2493.650 2039.740 2561.250 2187.860 ;
        RECT 2493.650 9.240 2494.550 2039.740 ;
        RECT 2496.950 1998.840 2561.250 2039.740 ;
        RECT 2496.950 1785.400 2531.950 1998.840 ;
        RECT 2534.350 1785.400 2535.630 1998.840 ;
        RECT 2538.030 1785.400 2561.250 1998.840 ;
        RECT 2496.950 1487.480 2561.250 1785.400 ;
        RECT 2496.950 1274.040 2531.950 1487.480 ;
        RECT 2534.350 1274.040 2535.630 1487.480 ;
        RECT 2538.030 1274.040 2561.250 1487.480 ;
        RECT 2496.950 978.840 2561.250 1274.040 ;
        RECT 2496.950 765.400 2531.950 978.840 ;
        RECT 2534.350 765.400 2535.630 978.840 ;
        RECT 2538.030 765.400 2561.250 978.840 ;
        RECT 2496.950 9.240 2561.250 765.400 ;
        RECT 2563.650 9.240 2564.550 2935.745 ;
        RECT 2566.950 9.240 2631.250 2935.745 ;
        RECT 2633.650 9.240 2634.550 2935.745 ;
        RECT 2636.950 9.240 2701.250 2935.745 ;
        RECT 2703.650 9.240 2704.550 2935.745 ;
        RECT 2706.950 9.240 2766.995 2935.745 ;
        RECT 26.905 8.695 2766.995 9.240 ;
  END
END fpga_top
END LIBRARY

