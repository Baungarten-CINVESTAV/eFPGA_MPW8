VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_4__4_
  CLASS BLOCK ;
  FOREIGN sb_4__4_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 146.000 26.130 149.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 146.000 16.470 149.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
  PIN bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 102.040 4.000 102.640 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 44.240 149.000 44.840 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 91.840 149.000 92.440 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 146.000 84.090 149.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1.000 39.010 4.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1.000 58.330 4.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1.000 122.730 4.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 3.440 4.000 4.040 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 115.640 149.000 116.240 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 1.000 16.470 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1.000 129.170 4.000 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 122.440 4.000 123.040 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 146.000 125.950 149.000 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.840 149.000 75.440 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 146.000 45.450 149.000 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 139.440 4.000 140.040 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 98.640 4.000 99.240 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1.000 145.270 4.000 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 68.040 4.000 68.640 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 129.240 149.000 129.840 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 17.040 149.000 17.640 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 146.000 96.970 149.000 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 78.240 4.000 78.840 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 146.000 55.110 149.000 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 146.000 61.550 149.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 146.000 109.850 149.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 108.840 4.000 109.440 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 142.840 149.000 143.440 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 122.440 149.000 123.040 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 136.040 149.000 136.640 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 30.640 149.000 31.240 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 146.000 90.530 149.000 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 146.000 67.990 149.000 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 17.040 4.000 17.640 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 146.240 4.000 146.840 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1.000 32.570 4.000 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 105.440 149.000 106.040 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 1.000 138.830 4.000 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 54.440 149.000 55.040 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 146.000 80.870 149.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 146.000 51.890 149.000 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 0.040 149.000 0.640 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 112.240 149.000 112.840 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 146.000 145.270 149.000 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 23.840 4.000 24.440 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 1.000 51.890 4.000 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 23.840 149.000 24.440 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 85.040 4.000 85.640 ;
    END
  END chanx_left_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 10.240 4.000 10.840 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 115.640 4.000 116.240 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 146.000 39.010 149.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1.000 109.850 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 146.000 132.390 149.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 1.000 93.750 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 1.000 10.030 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 71.440 4.000 72.040 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 1.000 132.390 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 61.240 149.000 61.840 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 37.440 149.000 38.040 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1.000 103.410 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 129.240 4.000 129.840 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 6.840 149.000 7.440 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 146.000 19.690 149.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 47.640 149.000 48.240 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 61.240 4.000 61.840 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 1.000 116.290 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 98.640 149.000 99.240 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1.000 67.990 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 91.840 4.000 92.440 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 1.000 74.430 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1.000 87.310 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 30.640 4.000 31.240 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 146.000 74.430 149.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 47.640 4.000 48.240 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 146.000 3.590 149.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1.000 22.910 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 1.000 3.590 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 146.000 138.830 149.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 146.000 103.410 149.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1.000 64.770 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 146.000 148.490 149.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 10.240 149.000 10.840 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 34.040 4.000 34.640 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 78.240 149.000 78.840 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 1.000 29.350 4.000 ;
    END
  END chany_bottom_out[9]
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 1.000 45.450 4.000 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 54.440 4.000 55.040 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 85.040 149.000 85.640 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1.000 80.870 4.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 146.000 119.510 149.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 146.000 116.290 149.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 146.000 10.030 149.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 146.000 32.570 149.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 1.000 96.970 4.000 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
  PIN left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 40.840 4.000 41.440 ;
    END
  END left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
  PIN pReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 136.040 4.000 136.640 ;
    END
  END pReset
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 68.040 149.000 68.640 ;
    END
  END prog_clk
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 10.640 23.685 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 10.640 58.415 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 10.640 93.145 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 10.640 127.875 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.450 10.640 41.050 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.180 10.640 75.780 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.910 10.640 110.510 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.640 10.640 145.240 138.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 0.070 6.840 149.890 138.960 ;
      LAYER met2 ;
        RECT 0.100 145.720 3.030 146.725 ;
        RECT 3.870 145.720 9.470 146.725 ;
        RECT 10.310 145.720 15.910 146.725 ;
        RECT 16.750 145.720 19.130 146.725 ;
        RECT 19.970 145.720 25.570 146.725 ;
        RECT 26.410 145.720 32.010 146.725 ;
        RECT 32.850 145.720 38.450 146.725 ;
        RECT 39.290 145.720 44.890 146.725 ;
        RECT 45.730 145.720 51.330 146.725 ;
        RECT 52.170 145.720 54.550 146.725 ;
        RECT 55.390 145.720 60.990 146.725 ;
        RECT 61.830 145.720 67.430 146.725 ;
        RECT 68.270 145.720 73.870 146.725 ;
        RECT 74.710 145.720 80.310 146.725 ;
        RECT 81.150 145.720 83.530 146.725 ;
        RECT 84.370 145.720 89.970 146.725 ;
        RECT 90.810 145.720 96.410 146.725 ;
        RECT 97.250 145.720 102.850 146.725 ;
        RECT 103.690 145.720 109.290 146.725 ;
        RECT 110.130 145.720 115.730 146.725 ;
        RECT 116.570 145.720 118.950 146.725 ;
        RECT 119.790 145.720 125.390 146.725 ;
        RECT 126.230 145.720 131.830 146.725 ;
        RECT 132.670 145.720 138.270 146.725 ;
        RECT 139.110 145.720 144.710 146.725 ;
        RECT 145.550 145.720 147.930 146.725 ;
        RECT 148.770 145.720 149.870 146.725 ;
        RECT 0.100 4.280 149.870 145.720 ;
        RECT 0.650 0.720 3.030 4.280 ;
        RECT 3.870 0.720 9.470 4.280 ;
        RECT 10.310 0.720 15.910 4.280 ;
        RECT 16.750 0.720 22.350 4.280 ;
        RECT 23.190 0.720 28.790 4.280 ;
        RECT 29.630 0.720 32.010 4.280 ;
        RECT 32.850 0.720 38.450 4.280 ;
        RECT 39.290 0.720 44.890 4.280 ;
        RECT 45.730 0.720 51.330 4.280 ;
        RECT 52.170 0.720 57.770 4.280 ;
        RECT 58.610 0.720 64.210 4.280 ;
        RECT 65.050 0.720 67.430 4.280 ;
        RECT 68.270 0.720 73.870 4.280 ;
        RECT 74.710 0.720 80.310 4.280 ;
        RECT 81.150 0.720 86.750 4.280 ;
        RECT 87.590 0.720 93.190 4.280 ;
        RECT 94.030 0.720 96.410 4.280 ;
        RECT 97.250 0.720 102.850 4.280 ;
        RECT 103.690 0.720 109.290 4.280 ;
        RECT 110.130 0.720 115.730 4.280 ;
        RECT 116.570 0.720 122.170 4.280 ;
        RECT 123.010 0.720 128.610 4.280 ;
        RECT 129.450 0.720 131.830 4.280 ;
        RECT 132.670 0.720 138.270 4.280 ;
        RECT 139.110 0.720 144.710 4.280 ;
        RECT 145.550 0.720 149.870 4.280 ;
        RECT 0.100 0.155 149.870 0.720 ;
      LAYER met3 ;
        RECT 4.400 145.840 149.895 146.705 ;
        RECT 4.000 143.840 149.895 145.840 ;
        RECT 4.000 142.440 145.600 143.840 ;
        RECT 149.400 142.440 149.895 143.840 ;
        RECT 4.000 140.440 149.895 142.440 ;
        RECT 4.400 139.040 149.895 140.440 ;
        RECT 4.000 137.040 149.895 139.040 ;
        RECT 4.400 135.640 145.600 137.040 ;
        RECT 149.400 135.640 149.895 137.040 ;
        RECT 4.000 130.240 149.895 135.640 ;
        RECT 4.400 128.840 145.600 130.240 ;
        RECT 149.400 128.840 149.895 130.240 ;
        RECT 4.000 123.440 149.895 128.840 ;
        RECT 4.400 122.040 145.600 123.440 ;
        RECT 149.400 122.040 149.895 123.440 ;
        RECT 4.000 116.640 149.895 122.040 ;
        RECT 4.400 115.240 145.600 116.640 ;
        RECT 149.400 115.240 149.895 116.640 ;
        RECT 4.000 113.240 149.895 115.240 ;
        RECT 4.000 111.840 145.600 113.240 ;
        RECT 149.400 111.840 149.895 113.240 ;
        RECT 4.000 109.840 149.895 111.840 ;
        RECT 4.400 108.440 149.895 109.840 ;
        RECT 4.000 106.440 149.895 108.440 ;
        RECT 4.000 105.040 145.600 106.440 ;
        RECT 149.400 105.040 149.895 106.440 ;
        RECT 4.000 103.040 149.895 105.040 ;
        RECT 4.400 101.640 149.895 103.040 ;
        RECT 4.000 99.640 149.895 101.640 ;
        RECT 4.400 98.240 145.600 99.640 ;
        RECT 149.400 98.240 149.895 99.640 ;
        RECT 4.000 92.840 149.895 98.240 ;
        RECT 4.400 91.440 145.600 92.840 ;
        RECT 149.400 91.440 149.895 92.840 ;
        RECT 4.000 86.040 149.895 91.440 ;
        RECT 4.400 84.640 145.600 86.040 ;
        RECT 149.400 84.640 149.895 86.040 ;
        RECT 4.000 79.240 149.895 84.640 ;
        RECT 4.400 77.840 145.600 79.240 ;
        RECT 149.400 77.840 149.895 79.240 ;
        RECT 4.000 75.840 149.895 77.840 ;
        RECT 4.000 74.440 145.600 75.840 ;
        RECT 149.400 74.440 149.895 75.840 ;
        RECT 4.000 72.440 149.895 74.440 ;
        RECT 4.400 71.040 149.895 72.440 ;
        RECT 4.000 69.040 149.895 71.040 ;
        RECT 4.400 67.640 145.600 69.040 ;
        RECT 149.400 67.640 149.895 69.040 ;
        RECT 4.000 62.240 149.895 67.640 ;
        RECT 4.400 60.840 145.600 62.240 ;
        RECT 149.400 60.840 149.895 62.240 ;
        RECT 4.000 55.440 149.895 60.840 ;
        RECT 4.400 54.040 145.600 55.440 ;
        RECT 149.400 54.040 149.895 55.440 ;
        RECT 4.000 48.640 149.895 54.040 ;
        RECT 4.400 47.240 145.600 48.640 ;
        RECT 149.400 47.240 149.895 48.640 ;
        RECT 4.000 45.240 149.895 47.240 ;
        RECT 4.000 43.840 145.600 45.240 ;
        RECT 149.400 43.840 149.895 45.240 ;
        RECT 4.000 41.840 149.895 43.840 ;
        RECT 4.400 40.440 149.895 41.840 ;
        RECT 4.000 38.440 149.895 40.440 ;
        RECT 4.000 37.040 145.600 38.440 ;
        RECT 149.400 37.040 149.895 38.440 ;
        RECT 4.000 35.040 149.895 37.040 ;
        RECT 4.400 33.640 149.895 35.040 ;
        RECT 4.000 31.640 149.895 33.640 ;
        RECT 4.400 30.240 145.600 31.640 ;
        RECT 149.400 30.240 149.895 31.640 ;
        RECT 4.000 24.840 149.895 30.240 ;
        RECT 4.400 23.440 145.600 24.840 ;
        RECT 149.400 23.440 149.895 24.840 ;
        RECT 4.000 18.040 149.895 23.440 ;
        RECT 4.400 16.640 145.600 18.040 ;
        RECT 149.400 16.640 149.895 18.040 ;
        RECT 4.000 11.240 149.895 16.640 ;
        RECT 4.400 9.840 145.600 11.240 ;
        RECT 149.400 9.840 149.895 11.240 ;
        RECT 4.000 7.840 149.895 9.840 ;
        RECT 4.000 6.440 145.600 7.840 ;
        RECT 149.400 6.440 149.895 7.840 ;
        RECT 4.000 4.440 149.895 6.440 ;
        RECT 4.400 3.040 149.895 4.440 ;
        RECT 4.000 1.040 149.895 3.040 ;
        RECT 4.000 0.175 145.600 1.040 ;
        RECT 149.400 0.175 149.895 1.040 ;
      LAYER met4 ;
        RECT 64.695 15.135 73.780 126.985 ;
        RECT 76.180 15.135 91.145 126.985 ;
        RECT 93.545 15.135 108.510 126.985 ;
        RECT 110.910 15.135 119.305 126.985 ;
  END
END sb_4__4_
END LIBRARY

