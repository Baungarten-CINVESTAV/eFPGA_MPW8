magic
tech sky130A
magscale 1 2
timestamp 1672416658
<< viali >>
rect 16221 37417 16255 37451
rect 26617 37417 26651 37451
rect 34253 37417 34287 37451
rect 9781 37281 9815 37315
rect 11161 37281 11195 37315
rect 11897 37281 11931 37315
rect 12357 37281 12391 37315
rect 16865 37281 16899 37315
rect 19625 37281 19659 37315
rect 20085 37281 20119 37315
rect 24041 37281 24075 37315
rect 24593 37281 24627 37315
rect 27169 37281 27203 37315
rect 34897 37281 34931 37315
rect 1869 37213 1903 37247
rect 2329 37213 2363 37247
rect 3985 37213 4019 37247
rect 5549 37213 5583 37247
rect 7481 37213 7515 37247
rect 9137 37213 9171 37247
rect 10885 37213 10919 37247
rect 12633 37213 12667 37247
rect 14289 37213 14323 37247
rect 17141 37213 17175 37247
rect 18153 37213 18187 37247
rect 20361 37213 20395 37247
rect 22017 37213 22051 37247
rect 23765 37213 23799 37247
rect 25237 37213 25271 37247
rect 27353 37213 27387 37247
rect 29745 37213 29779 37247
rect 30481 37213 30515 37247
rect 32321 37213 32355 37247
rect 35081 37213 35115 37247
rect 36461 37213 36495 37247
rect 38025 37213 38059 37247
rect 3065 37145 3099 37179
rect 1685 37077 1719 37111
rect 2513 37077 2547 37111
rect 4169 37077 4203 37111
rect 5365 37077 5399 37111
rect 7297 37077 7331 37111
rect 8033 37077 8067 37111
rect 9321 37077 9355 37111
rect 14473 37077 14507 37111
rect 18337 37077 18371 37111
rect 22201 37077 22235 37111
rect 25421 37077 25455 37111
rect 29929 37077 29963 37111
rect 30665 37077 30699 37111
rect 32505 37077 32539 37111
rect 36277 37077 36311 37111
rect 38209 37077 38243 37111
rect 3433 36873 3467 36907
rect 11713 36873 11747 36907
rect 17877 36873 17911 36907
rect 20729 36873 20763 36907
rect 21373 36873 21407 36907
rect 30113 36873 30147 36907
rect 38209 36873 38243 36907
rect 1685 36805 1719 36839
rect 3617 36737 3651 36771
rect 17693 36737 17727 36771
rect 21189 36737 21223 36771
rect 24041 36737 24075 36771
rect 24685 36737 24719 36771
rect 25973 36737 26007 36771
rect 27169 36737 27203 36771
rect 30021 36737 30055 36771
rect 30665 36737 30699 36771
rect 38025 36737 38059 36771
rect 25421 36669 25455 36703
rect 1869 36601 1903 36635
rect 26157 36601 26191 36635
rect 27353 36601 27387 36635
rect 2329 36533 2363 36567
rect 4169 36533 4203 36567
rect 24225 36533 24259 36567
rect 36553 36533 36587 36567
rect 2329 36329 2363 36363
rect 1869 36125 1903 36159
rect 38025 36125 38059 36159
rect 1685 35989 1719 36023
rect 38209 35989 38243 36023
rect 1961 35785 1995 35819
rect 38209 35785 38243 35819
rect 2053 35649 2087 35683
rect 38025 35649 38059 35683
rect 2513 35445 2547 35479
rect 1869 34561 1903 34595
rect 38025 34561 38059 34595
rect 2329 34493 2363 34527
rect 37473 34493 37507 34527
rect 1685 34357 1719 34391
rect 38209 34357 38243 34391
rect 1685 32385 1719 32419
rect 25513 32385 25547 32419
rect 38025 32385 38059 32419
rect 38301 32317 38335 32351
rect 1869 32249 1903 32283
rect 25421 32181 25455 32215
rect 1593 31977 1627 32011
rect 38301 31977 38335 32011
rect 23857 31433 23891 31467
rect 23673 31297 23707 31331
rect 25513 31297 25547 31331
rect 24317 31093 24351 31127
rect 25421 31093 25455 31127
rect 1869 30685 1903 30719
rect 10977 30685 11011 30719
rect 22937 30685 22971 30719
rect 11253 30617 11287 30651
rect 1685 30549 1719 30583
rect 2329 30549 2363 30583
rect 23029 30549 23063 30583
rect 18797 30209 18831 30243
rect 38025 30141 38059 30175
rect 38301 30141 38335 30175
rect 18889 30005 18923 30039
rect 38301 29801 38335 29835
rect 14197 29257 14231 29291
rect 1869 29121 1903 29155
rect 14013 29121 14047 29155
rect 22753 29121 22787 29155
rect 23397 29121 23431 29155
rect 38025 29121 38059 29155
rect 1685 28985 1719 29019
rect 14749 28985 14783 29019
rect 22845 28985 22879 29019
rect 38209 28985 38243 29019
rect 23029 28509 23063 28543
rect 23673 28509 23707 28543
rect 23213 28373 23247 28407
rect 23121 28169 23155 28203
rect 26157 28169 26191 28203
rect 22569 28033 22603 28067
rect 25513 28033 25547 28067
rect 22477 27829 22511 27863
rect 25605 27829 25639 27863
rect 1593 26877 1627 26911
rect 1869 26877 1903 26911
rect 38025 26877 38059 26911
rect 38301 26877 38335 26911
rect 1593 26537 1627 26571
rect 23121 26537 23155 26571
rect 38301 26537 38335 26571
rect 16037 26469 16071 26503
rect 16773 26401 16807 26435
rect 16221 26333 16255 26367
rect 22477 26333 22511 26367
rect 22569 26265 22603 26299
rect 1869 24769 1903 24803
rect 37565 24769 37599 24803
rect 38209 24769 38243 24803
rect 38025 24633 38059 24667
rect 1685 24565 1719 24599
rect 25789 24361 25823 24395
rect 28733 23817 28767 23851
rect 23857 23749 23891 23783
rect 24777 23749 24811 23783
rect 26249 23749 26283 23783
rect 22385 23681 22419 23715
rect 23029 23681 23063 23715
rect 25605 23681 25639 23715
rect 26341 23681 26375 23715
rect 27169 23681 27203 23715
rect 28549 23681 28583 23715
rect 29193 23681 29227 23715
rect 22569 23613 22603 23647
rect 24869 23613 24903 23647
rect 25421 23545 25455 23579
rect 7297 23273 7331 23307
rect 23305 23273 23339 23307
rect 25973 23273 26007 23307
rect 22661 23137 22695 23171
rect 7481 23069 7515 23103
rect 22845 23069 22879 23103
rect 25513 23069 25547 23103
rect 1685 22933 1719 22967
rect 8033 22933 8067 22967
rect 25421 22933 25455 22967
rect 25421 22661 25455 22695
rect 25513 22661 25547 22695
rect 1685 22593 1719 22627
rect 38025 22593 38059 22627
rect 23029 22525 23063 22559
rect 1869 22457 1903 22491
rect 24961 22457 24995 22491
rect 38209 22457 38243 22491
rect 22385 22185 22419 22219
rect 23305 22185 23339 22219
rect 25053 22185 25087 22219
rect 22937 22049 22971 22083
rect 2237 21981 2271 22015
rect 21833 21981 21867 22015
rect 22293 21981 22327 22015
rect 23121 21981 23155 22015
rect 24961 21981 24995 22015
rect 25605 21981 25639 22015
rect 2053 21845 2087 21879
rect 2789 21845 2823 21879
rect 22477 21641 22511 21675
rect 23121 21641 23155 21675
rect 24777 21641 24811 21675
rect 22385 21505 22419 21539
rect 23213 21505 23247 21539
rect 24133 21505 24167 21539
rect 24225 21301 24259 21335
rect 30297 21029 30331 21063
rect 23489 20893 23523 20927
rect 24685 20893 24719 20927
rect 30113 20893 30147 20927
rect 30757 20893 30791 20927
rect 38025 20893 38059 20927
rect 1685 20825 1719 20859
rect 1869 20825 1903 20859
rect 19809 20825 19843 20859
rect 20361 20825 20395 20859
rect 19717 20757 19751 20791
rect 22753 20757 22787 20791
rect 23397 20757 23431 20791
rect 24041 20757 24075 20791
rect 38209 20757 38243 20791
rect 22201 20553 22235 20587
rect 38025 20553 38059 20587
rect 1593 20485 1627 20519
rect 23489 20485 23523 20519
rect 25329 20485 25363 20519
rect 22661 20417 22695 20451
rect 27353 20417 27387 20451
rect 37841 20417 37875 20451
rect 23397 20349 23431 20383
rect 24041 20349 24075 20383
rect 24961 20349 24995 20383
rect 25421 20349 25455 20383
rect 22753 20213 22787 20247
rect 27261 20213 27295 20247
rect 27905 20213 27939 20247
rect 23673 20009 23707 20043
rect 24869 20009 24903 20043
rect 9137 19941 9171 19975
rect 16589 19805 16623 19839
rect 17233 19805 17267 19839
rect 22477 19805 22511 19839
rect 22661 19805 22695 19839
rect 23765 19805 23799 19839
rect 24777 19805 24811 19839
rect 9321 19737 9355 19771
rect 16681 19737 16715 19771
rect 22017 19737 22051 19771
rect 25421 19737 25455 19771
rect 9873 19669 9907 19703
rect 23121 19669 23155 19703
rect 25973 19669 26007 19703
rect 37657 19669 37691 19703
rect 23305 19465 23339 19499
rect 22201 19397 22235 19431
rect 24225 19397 24259 19431
rect 25145 19397 25179 19431
rect 25237 19397 25271 19431
rect 26341 19397 26375 19431
rect 26433 19397 26467 19431
rect 1869 19329 1903 19363
rect 23397 19329 23431 19363
rect 38025 19329 38059 19363
rect 1593 19261 1627 19295
rect 22109 19261 22143 19295
rect 22661 19193 22695 19227
rect 25881 19193 25915 19227
rect 38209 19125 38243 19159
rect 1593 18921 1627 18955
rect 25973 18921 26007 18955
rect 38025 18921 38059 18955
rect 10333 18853 10367 18887
rect 21649 18785 21683 18819
rect 22293 18785 22327 18819
rect 23121 18785 23155 18819
rect 23397 18785 23431 18819
rect 10241 18717 10275 18751
rect 10885 18717 10919 18751
rect 24777 18717 24811 18751
rect 25421 18717 25455 18751
rect 25881 18717 25915 18751
rect 26525 18717 26559 18751
rect 27629 18717 27663 18751
rect 37841 18717 37875 18751
rect 21741 18649 21775 18683
rect 23213 18649 23247 18683
rect 27077 18649 27111 18683
rect 21097 18581 21131 18615
rect 24685 18581 24719 18615
rect 25329 18581 25363 18615
rect 21373 18377 21407 18411
rect 22753 18309 22787 18343
rect 25421 18309 25455 18343
rect 25513 18309 25547 18343
rect 26433 18309 26467 18343
rect 21281 18241 21315 18275
rect 23765 18241 23799 18275
rect 23949 18241 23983 18275
rect 22661 18173 22695 18207
rect 23121 18173 23155 18207
rect 24133 18105 24167 18139
rect 22109 18037 22143 18071
rect 27169 18037 27203 18071
rect 38117 18037 38151 18071
rect 21741 17833 21775 17867
rect 22385 17833 22419 17867
rect 27537 17833 27571 17867
rect 29837 17833 29871 17867
rect 24961 17765 24995 17799
rect 26893 17765 26927 17799
rect 20637 17697 20671 17731
rect 23029 17697 23063 17731
rect 24041 17697 24075 17731
rect 25697 17697 25731 17731
rect 21833 17629 21867 17663
rect 22477 17629 22511 17663
rect 24593 17629 24627 17663
rect 24777 17629 24811 17663
rect 25881 17629 25915 17663
rect 26985 17629 27019 17663
rect 27629 17629 27663 17663
rect 29745 17629 29779 17663
rect 23121 17561 23155 17595
rect 21189 17493 21223 17527
rect 26341 17493 26375 17527
rect 28181 17493 28215 17527
rect 24317 17289 24351 17323
rect 27905 17289 27939 17323
rect 22477 17221 22511 17255
rect 23213 17221 23247 17255
rect 25237 17221 25271 17255
rect 25329 17221 25363 17255
rect 26249 17221 26283 17255
rect 1869 17153 1903 17187
rect 20913 17153 20947 17187
rect 22385 17153 22419 17187
rect 24225 17153 24259 17187
rect 27813 17153 27847 17187
rect 37657 17153 37691 17187
rect 38301 17153 38335 17187
rect 23121 17085 23155 17119
rect 27169 17085 27203 17119
rect 1685 17017 1719 17051
rect 23673 17017 23707 17051
rect 28457 17017 28491 17051
rect 21373 16949 21407 16983
rect 38117 16949 38151 16983
rect 2421 16745 2455 16779
rect 28181 16745 28215 16779
rect 23121 16677 23155 16711
rect 10793 16609 10827 16643
rect 20085 16609 20119 16643
rect 25329 16609 25363 16643
rect 26157 16609 26191 16643
rect 1961 16541 1995 16575
rect 10149 16541 10183 16575
rect 21189 16541 21223 16575
rect 22017 16541 22051 16575
rect 23949 16541 23983 16575
rect 24593 16541 24627 16575
rect 26985 16541 27019 16575
rect 27629 16541 27663 16575
rect 10241 16473 10275 16507
rect 20269 16473 20303 16507
rect 21281 16473 21315 16507
rect 22569 16473 22603 16507
rect 22661 16473 22695 16507
rect 23673 16473 23707 16507
rect 25421 16473 25455 16507
rect 1777 16405 1811 16439
rect 21833 16405 21867 16439
rect 24685 16405 24719 16439
rect 26893 16405 26927 16439
rect 27537 16405 27571 16439
rect 21373 16201 21407 16235
rect 20545 16133 20579 16167
rect 23581 16133 23615 16167
rect 26065 16133 26099 16167
rect 21465 16065 21499 16099
rect 22937 16065 22971 16099
rect 24593 16065 24627 16099
rect 24777 16065 24811 16099
rect 26617 16065 26651 16099
rect 27169 16065 27203 16099
rect 22753 15997 22787 16031
rect 23489 15997 23523 16031
rect 25973 15997 26007 16031
rect 24041 15929 24075 15963
rect 22569 15861 22603 15895
rect 25237 15861 25271 15895
rect 27261 15861 27295 15895
rect 27905 15861 27939 15895
rect 6929 15657 6963 15691
rect 22201 15657 22235 15691
rect 27537 15657 27571 15691
rect 21557 15589 21591 15623
rect 25237 15589 25271 15623
rect 23121 15521 23155 15555
rect 24593 15521 24627 15555
rect 24777 15521 24811 15555
rect 25697 15521 25731 15555
rect 26157 15521 26191 15555
rect 1869 15453 1903 15487
rect 7113 15453 7147 15487
rect 22201 15453 22235 15487
rect 26341 15453 26375 15487
rect 26801 15453 26835 15487
rect 27629 15453 27663 15487
rect 28273 15453 28307 15487
rect 38025 15453 38059 15487
rect 7665 15385 7699 15419
rect 22845 15385 22879 15419
rect 22937 15385 22971 15419
rect 28825 15385 28859 15419
rect 1685 15317 1719 15351
rect 23949 15317 23983 15351
rect 26893 15317 26927 15351
rect 28181 15317 28215 15351
rect 38209 15317 38243 15351
rect 12173 15113 12207 15147
rect 22753 15113 22787 15147
rect 25789 15113 25823 15147
rect 28365 15113 28399 15147
rect 22201 15045 22235 15079
rect 23489 15045 23523 15079
rect 24041 15045 24075 15079
rect 24593 15045 24627 15079
rect 24685 15045 24719 15079
rect 26433 15045 26467 15079
rect 12357 14977 12391 15011
rect 21465 14977 21499 15011
rect 22661 14977 22695 15011
rect 25881 14977 25915 15011
rect 26525 14977 26559 15011
rect 27353 14977 27387 15011
rect 28457 14977 28491 15011
rect 23397 14909 23431 14943
rect 25237 14909 25271 14943
rect 27169 14909 27203 14943
rect 12909 14841 12943 14875
rect 27721 14773 27755 14807
rect 1961 14569 1995 14603
rect 35725 14569 35759 14603
rect 22109 14433 22143 14467
rect 22753 14433 22787 14467
rect 25237 14433 25271 14467
rect 26433 14433 26467 14467
rect 26801 14433 26835 14467
rect 27997 14433 28031 14467
rect 12081 14365 12115 14399
rect 12725 14365 12759 14399
rect 23397 14365 23431 14399
rect 23581 14365 23615 14399
rect 24041 14365 24075 14399
rect 24777 14365 24811 14399
rect 25421 14365 25455 14399
rect 35541 14365 35575 14399
rect 1869 14297 1903 14331
rect 2513 14297 2547 14331
rect 12173 14297 12207 14331
rect 22201 14297 22235 14331
rect 26709 14297 26743 14331
rect 27353 14297 27387 14331
rect 27905 14297 27939 14331
rect 38117 14229 38151 14263
rect 22201 14025 22235 14059
rect 23305 14025 23339 14059
rect 23949 14025 23983 14059
rect 27261 14025 27295 14059
rect 38025 14025 38059 14059
rect 25053 13957 25087 13991
rect 25145 13957 25179 13991
rect 25881 13957 25915 13991
rect 25973 13957 26007 13991
rect 19165 13889 19199 13923
rect 19809 13889 19843 13923
rect 21465 13889 21499 13923
rect 22293 13889 22327 13923
rect 23397 13889 23431 13923
rect 24041 13889 24075 13923
rect 26525 13889 26559 13923
rect 27353 13889 27387 13923
rect 37841 13889 37875 13923
rect 19257 13821 19291 13855
rect 24501 13821 24535 13855
rect 23949 13481 23983 13515
rect 26249 13481 26283 13515
rect 26985 13481 27019 13515
rect 22937 13413 22971 13447
rect 22385 13345 22419 13379
rect 1869 13277 1903 13311
rect 10517 13277 10551 13311
rect 11161 13277 11195 13311
rect 21649 13277 21683 13311
rect 24041 13277 24075 13311
rect 25789 13277 25823 13311
rect 25973 13277 26007 13311
rect 27077 13277 27111 13311
rect 38025 13277 38059 13311
rect 22477 13209 22511 13243
rect 24593 13209 24627 13243
rect 25145 13209 25179 13243
rect 25237 13209 25271 13243
rect 1685 13141 1719 13175
rect 10609 13141 10643 13175
rect 21097 13141 21131 13175
rect 21741 13141 21775 13175
rect 38209 13141 38243 13175
rect 25697 12937 25731 12971
rect 26341 12937 26375 12971
rect 27261 12937 27295 12971
rect 27905 12937 27939 12971
rect 20821 12869 20855 12903
rect 23765 12869 23799 12903
rect 24409 12869 24443 12903
rect 24961 12869 24995 12903
rect 22661 12801 22695 12835
rect 25605 12801 25639 12835
rect 26433 12801 26467 12835
rect 27353 12801 27387 12835
rect 27997 12801 28031 12835
rect 28641 12801 28675 12835
rect 20729 12733 20763 12767
rect 21373 12733 21407 12767
rect 23213 12733 23247 12767
rect 23857 12733 23891 12767
rect 25053 12733 25087 12767
rect 22661 12665 22695 12699
rect 20177 12597 20211 12631
rect 28549 12597 28583 12631
rect 29193 12597 29227 12631
rect 4353 12393 4387 12427
rect 20729 12393 20763 12427
rect 28457 12393 28491 12427
rect 17233 12257 17267 12291
rect 22293 12257 22327 12291
rect 24961 12257 24995 12291
rect 25973 12257 26007 12291
rect 26525 12257 26559 12291
rect 27169 12257 27203 12291
rect 4445 12189 4479 12223
rect 17141 12189 17175 12223
rect 17785 12189 17819 12223
rect 20177 12189 20211 12223
rect 20637 12189 20671 12223
rect 27905 12189 27939 12223
rect 28549 12189 28583 12223
rect 21465 12121 21499 12155
rect 22017 12121 22051 12155
rect 22109 12121 22143 12155
rect 23213 12121 23247 12155
rect 23305 12121 23339 12155
rect 23857 12121 23891 12155
rect 25881 12121 25915 12155
rect 27077 12121 27111 12155
rect 4997 12053 5031 12087
rect 27813 12053 27847 12087
rect 26065 11849 26099 11883
rect 27261 11849 27295 11883
rect 22201 11781 22235 11815
rect 22293 11781 22327 11815
rect 24501 11781 24535 11815
rect 24593 11781 24627 11815
rect 20821 11713 20855 11747
rect 21465 11713 21499 11747
rect 23305 11713 23339 11747
rect 26157 11713 26191 11747
rect 27353 11713 27387 11747
rect 27813 11713 27847 11747
rect 24869 11645 24903 11679
rect 22753 11577 22787 11611
rect 23489 11577 23523 11611
rect 27905 11577 27939 11611
rect 21281 11509 21315 11543
rect 16405 11305 16439 11339
rect 22385 11305 22419 11339
rect 23029 11305 23063 11339
rect 23673 11305 23707 11339
rect 24961 11169 24995 11203
rect 26433 11169 26467 11203
rect 38025 11169 38059 11203
rect 1869 11101 1903 11135
rect 15761 11101 15795 11135
rect 21097 11101 21131 11135
rect 21557 11101 21591 11135
rect 22477 11101 22511 11135
rect 23121 11101 23155 11135
rect 23765 11101 23799 11135
rect 27353 11101 27387 11135
rect 38301 11101 38335 11135
rect 21833 11033 21867 11067
rect 24685 11033 24719 11067
rect 24777 11033 24811 11067
rect 26709 11033 26743 11067
rect 26801 11033 26835 11067
rect 27997 11033 28031 11067
rect 1685 10965 1719 10999
rect 15945 10965 15979 10999
rect 23305 10761 23339 10795
rect 24225 10761 24259 10795
rect 36277 10761 36311 10795
rect 38301 10761 38335 10795
rect 2053 10693 2087 10727
rect 15761 10693 15795 10727
rect 22098 10693 22132 10727
rect 22201 10693 22235 10727
rect 25421 10693 25455 10727
rect 26341 10693 26375 10727
rect 29193 10693 29227 10727
rect 31217 10693 31251 10727
rect 1869 10625 1903 10659
rect 21373 10625 21407 10659
rect 21465 10625 21499 10659
rect 23397 10625 23431 10659
rect 24133 10625 24167 10659
rect 29101 10625 29135 10659
rect 36185 10625 36219 10659
rect 15669 10557 15703 10591
rect 25329 10557 25363 10591
rect 31309 10557 31343 10591
rect 16221 10489 16255 10523
rect 22661 10489 22695 10523
rect 30757 10489 30791 10523
rect 14381 10217 14415 10251
rect 17233 10217 17267 10251
rect 17877 10217 17911 10251
rect 33609 10217 33643 10251
rect 23397 10149 23431 10183
rect 1869 10081 1903 10115
rect 22937 10081 22971 10115
rect 25605 10081 25639 10115
rect 26617 10081 26651 10115
rect 1593 10013 1627 10047
rect 14289 10013 14323 10047
rect 17325 10013 17359 10047
rect 24593 10013 24627 10047
rect 27353 10013 27387 10047
rect 33701 10013 33735 10047
rect 22293 9945 22327 9979
rect 22385 9945 22419 9979
rect 26525 9945 26559 9979
rect 24685 9877 24719 9911
rect 27261 9877 27295 9911
rect 22293 9673 22327 9707
rect 1593 9605 1627 9639
rect 24685 9605 24719 9639
rect 25329 9605 25363 9639
rect 26249 9605 26283 9639
rect 22201 9537 22235 9571
rect 24133 9469 24167 9503
rect 24777 9469 24811 9503
rect 26341 9469 26375 9503
rect 20913 9129 20947 9163
rect 23489 9129 23523 9163
rect 25053 9129 25087 9163
rect 38117 9129 38151 9163
rect 25697 9061 25731 9095
rect 22109 8993 22143 9027
rect 26433 8993 26467 9027
rect 20821 8925 20855 8959
rect 23581 8925 23615 8959
rect 25145 8925 25179 8959
rect 25789 8925 25823 8959
rect 30757 8925 30791 8959
rect 21465 8857 21499 8891
rect 22017 8857 22051 8891
rect 37565 8857 37599 8891
rect 38209 8857 38243 8891
rect 27261 8789 27295 8823
rect 29837 8789 29871 8823
rect 25421 8585 25455 8619
rect 26065 8585 26099 8619
rect 27537 8585 27571 8619
rect 22293 8517 22327 8551
rect 23397 8517 23431 8551
rect 29009 8517 29043 8551
rect 22385 8449 22419 8483
rect 25513 8449 25547 8483
rect 26157 8449 26191 8483
rect 29285 8449 29319 8483
rect 31493 8449 31527 8483
rect 23121 8381 23155 8415
rect 24869 8381 24903 8415
rect 31217 8381 31251 8415
rect 21097 8313 21131 8347
rect 29745 8313 29779 8347
rect 24685 8041 24719 8075
rect 31493 8041 31527 8075
rect 25513 7973 25547 8007
rect 32045 7973 32079 8007
rect 21465 7905 21499 7939
rect 21741 7905 21775 7939
rect 32689 7905 32723 7939
rect 38025 7905 38059 7939
rect 1869 7837 1903 7871
rect 22293 7837 22327 7871
rect 24777 7837 24811 7871
rect 27261 7837 27295 7871
rect 29745 7837 29779 7871
rect 32137 7837 32171 7871
rect 32781 7837 32815 7871
rect 38301 7837 38335 7871
rect 21649 7769 21683 7803
rect 22569 7769 22603 7803
rect 26985 7769 27019 7803
rect 30021 7769 30055 7803
rect 1685 7701 1719 7735
rect 24041 7701 24075 7735
rect 27721 7701 27755 7735
rect 28549 7701 28583 7735
rect 29101 7701 29135 7735
rect 14105 7497 14139 7531
rect 21373 7497 21407 7531
rect 22477 7497 22511 7531
rect 23489 7497 23523 7531
rect 33057 7497 33091 7531
rect 33701 7497 33735 7531
rect 38301 7497 38335 7531
rect 30665 7429 30699 7463
rect 14289 7361 14323 7395
rect 21465 7361 21499 7395
rect 22569 7361 22603 7395
rect 31769 7361 31803 7395
rect 32505 7361 32539 7395
rect 33149 7361 33183 7395
rect 24961 7293 24995 7327
rect 25237 7293 25271 7327
rect 28630 7293 28664 7327
rect 28089 7225 28123 7259
rect 32413 7225 32447 7259
rect 14841 7157 14875 7191
rect 25789 7157 25823 7191
rect 26249 7157 26283 7191
rect 27629 7157 27663 7191
rect 28904 7157 28938 7191
rect 31677 7157 31711 7191
rect 22556 6953 22590 6987
rect 24856 6953 24890 6987
rect 28475 6953 28509 6987
rect 20637 6817 20671 6851
rect 22293 6817 22327 6851
rect 26341 6817 26375 6851
rect 28733 6817 28767 6851
rect 32781 6817 32815 6851
rect 34069 6817 34103 6851
rect 24593 6749 24627 6783
rect 29745 6749 29779 6783
rect 32137 6749 32171 6783
rect 32229 6749 32263 6783
rect 32873 6749 32907 6783
rect 33517 6749 33551 6783
rect 20821 6681 20855 6715
rect 20913 6681 20947 6715
rect 30021 6681 30055 6715
rect 33425 6681 33459 6715
rect 24041 6613 24075 6647
rect 26985 6613 27019 6647
rect 31493 6613 31527 6647
rect 34897 6613 34931 6647
rect 21373 6409 21407 6443
rect 31677 6409 31711 6443
rect 32413 6409 32447 6443
rect 22201 6341 22235 6375
rect 25053 6341 25087 6375
rect 27905 6341 27939 6375
rect 30389 6341 30423 6375
rect 33057 6341 33091 6375
rect 21465 6273 21499 6307
rect 29929 6273 29963 6307
rect 31125 6273 31159 6307
rect 31769 6273 31803 6307
rect 32505 6273 32539 6307
rect 33149 6273 33183 6307
rect 33609 6273 33643 6307
rect 34437 6273 34471 6307
rect 22109 6205 22143 6239
rect 25329 6205 25363 6239
rect 29653 6205 29687 6239
rect 22661 6137 22695 6171
rect 34345 6137 34379 6171
rect 23581 6069 23615 6103
rect 25789 6069 25823 6103
rect 26341 6069 26375 6103
rect 27169 6069 27203 6103
rect 31033 6069 31067 6103
rect 33701 6069 33735 6103
rect 34897 6069 34931 6103
rect 35541 6069 35575 6103
rect 36093 6069 36127 6103
rect 37657 6069 37691 6103
rect 38209 6069 38243 6103
rect 33885 5865 33919 5899
rect 38117 5865 38151 5899
rect 26985 5797 27019 5831
rect 29193 5797 29227 5831
rect 25513 5729 25547 5763
rect 27721 5729 27755 5763
rect 34989 5729 35023 5763
rect 1869 5661 1903 5695
rect 4997 5661 5031 5695
rect 5089 5661 5123 5695
rect 25237 5661 25271 5695
rect 27445 5661 27479 5695
rect 31493 5661 31527 5695
rect 32137 5661 32171 5695
rect 32873 5661 32907 5695
rect 33977 5661 34011 5695
rect 34897 5661 34931 5695
rect 37657 5661 37691 5695
rect 38301 5661 38335 5695
rect 31217 5593 31251 5627
rect 33149 5593 33183 5627
rect 36645 5593 36679 5627
rect 1685 5525 1719 5559
rect 5641 5525 5675 5559
rect 21833 5525 21867 5559
rect 22293 5525 22327 5559
rect 24593 5525 24627 5559
rect 29745 5525 29779 5559
rect 32045 5525 32079 5559
rect 35541 5525 35575 5559
rect 36093 5525 36127 5559
rect 22109 5321 22143 5355
rect 25697 5321 25731 5355
rect 26525 5321 26559 5355
rect 27169 5321 27203 5355
rect 27721 5321 27755 5355
rect 30113 5321 30147 5355
rect 28641 5253 28675 5287
rect 33149 5253 33183 5287
rect 35357 5253 35391 5287
rect 35909 5253 35943 5287
rect 36461 5253 36495 5287
rect 20361 5185 20395 5219
rect 21097 5185 21131 5219
rect 21189 5185 21223 5219
rect 22201 5185 22235 5219
rect 22845 5185 22879 5219
rect 28365 5185 28399 5219
rect 31125 5185 31159 5219
rect 31769 5185 31803 5219
rect 32873 5185 32907 5219
rect 34253 5185 34287 5219
rect 34897 5185 34931 5219
rect 20545 5117 20579 5151
rect 23397 5117 23431 5151
rect 23673 5117 23707 5151
rect 25145 5117 25179 5151
rect 31033 5117 31067 5151
rect 33977 5117 34011 5151
rect 20177 5049 20211 5083
rect 22753 4981 22787 5015
rect 31677 4981 31711 5015
rect 32321 4981 32355 5015
rect 34805 4981 34839 5015
rect 37473 4981 37507 5015
rect 38301 4981 38335 5015
rect 21649 4777 21683 4811
rect 24041 4777 24075 4811
rect 26341 4777 26375 4811
rect 29009 4777 29043 4811
rect 31493 4777 31527 4811
rect 32137 4777 32171 4811
rect 34069 4777 34103 4811
rect 36553 4777 36587 4811
rect 28549 4709 28583 4743
rect 32781 4709 32815 4743
rect 22109 4641 22143 4675
rect 24869 4641 24903 4675
rect 27077 4641 27111 4675
rect 29745 4641 29779 4675
rect 37105 4641 37139 4675
rect 22293 4573 22327 4607
rect 24593 4573 24627 4607
rect 26801 4573 26835 4607
rect 32229 4573 32263 4607
rect 32873 4573 32907 4607
rect 33517 4573 33551 4607
rect 34161 4573 34195 4607
rect 37841 4573 37875 4607
rect 30021 4505 30055 4539
rect 20637 4437 20671 4471
rect 22937 4437 22971 4471
rect 23397 4437 23431 4471
rect 33425 4437 33459 4471
rect 34897 4437 34931 4471
rect 35449 4437 35483 4471
rect 36001 4437 36035 4471
rect 38025 4437 38059 4471
rect 20361 4233 20395 4267
rect 25881 4233 25915 4267
rect 36001 4233 36035 4267
rect 31677 4165 31711 4199
rect 20269 4097 20303 4131
rect 21097 4097 21131 4131
rect 22385 4097 22419 4131
rect 22937 4097 22971 4131
rect 25421 4097 25455 4131
rect 26433 4097 26467 4131
rect 30205 4097 30239 4131
rect 31125 4097 31159 4131
rect 31769 4097 31803 4131
rect 32321 4097 32355 4131
rect 33149 4097 33183 4131
rect 33793 4097 33827 4131
rect 34437 4097 34471 4131
rect 38025 4097 38059 4131
rect 23397 4029 23431 4063
rect 23673 4029 23707 4063
rect 28457 4029 28491 4063
rect 29929 4029 29963 4063
rect 34345 4029 34379 4063
rect 36553 4029 36587 4063
rect 33057 3961 33091 3995
rect 37473 3961 37507 3995
rect 1593 3893 1627 3927
rect 21005 3893 21039 3927
rect 27261 3893 27295 3927
rect 27721 3893 27755 3927
rect 31033 3893 31067 3927
rect 32413 3893 32447 3927
rect 33701 3893 33735 3927
rect 34897 3893 34931 3927
rect 35449 3893 35483 3927
rect 38209 3893 38243 3927
rect 20453 3689 20487 3723
rect 21373 3689 21407 3723
rect 28641 3689 28675 3723
rect 34253 3689 34287 3723
rect 34989 3689 35023 3723
rect 35541 3689 35575 3723
rect 36093 3689 36127 3723
rect 31493 3621 31527 3655
rect 33701 3621 33735 3655
rect 20637 3553 20671 3587
rect 24869 3553 24903 3587
rect 26893 3553 26927 3587
rect 30021 3553 30055 3587
rect 32229 3553 32263 3587
rect 1869 3485 1903 3519
rect 19717 3485 19751 3519
rect 20821 3485 20855 3519
rect 22293 3485 22327 3519
rect 24593 3485 24627 3519
rect 29745 3485 29779 3519
rect 31953 3485 31987 3519
rect 34345 3485 34379 3519
rect 34897 3485 34931 3519
rect 38025 3485 38059 3519
rect 38301 3485 38335 3519
rect 2329 3417 2363 3451
rect 22569 3417 22603 3451
rect 27169 3417 27203 3451
rect 1685 3349 1719 3383
rect 19533 3349 19567 3383
rect 24041 3349 24075 3383
rect 26341 3349 26375 3383
rect 29101 3349 29135 3383
rect 36645 3349 36679 3383
rect 20637 3145 20671 3179
rect 21373 3145 21407 3179
rect 26525 3145 26559 3179
rect 27261 3145 27295 3179
rect 28089 3145 28123 3179
rect 35357 3145 35391 3179
rect 36369 3145 36403 3179
rect 3341 3077 3375 3111
rect 19533 3077 19567 3111
rect 22569 3077 22603 3111
rect 23581 3077 23615 3111
rect 25329 3077 25363 3111
rect 28181 3077 28215 3111
rect 34621 3077 34655 3111
rect 17509 3009 17543 3043
rect 19993 3009 20027 3043
rect 20821 3009 20855 3043
rect 21465 3009 21499 3043
rect 22109 3009 22143 3043
rect 22753 3009 22787 3043
rect 23305 3009 23339 3043
rect 25789 3009 25823 3043
rect 30757 3009 30791 3043
rect 31401 3009 31435 3043
rect 34713 3009 34747 3043
rect 35173 3009 35207 3043
rect 38025 3009 38059 3043
rect 38301 3009 38335 3043
rect 1593 2941 1627 2975
rect 1869 2941 1903 2975
rect 28733 2941 28767 2975
rect 30481 2941 30515 2975
rect 31217 2941 31251 2975
rect 33793 2941 33827 2975
rect 34069 2941 34103 2975
rect 5733 2873 5767 2907
rect 20177 2873 20211 2907
rect 35817 2873 35851 2907
rect 3801 2805 3835 2839
rect 17325 2805 17359 2839
rect 18061 2805 18095 2839
rect 25973 2805 26007 2839
rect 32321 2805 32355 2839
rect 4169 2601 4203 2635
rect 14473 2601 14507 2635
rect 27261 2601 27295 2635
rect 29745 2601 29779 2635
rect 33517 2601 33551 2635
rect 35633 2601 35667 2635
rect 9413 2533 9447 2567
rect 36461 2533 36495 2567
rect 1869 2465 1903 2499
rect 11161 2465 11195 2499
rect 11713 2465 11747 2499
rect 18337 2465 18371 2499
rect 22201 2465 22235 2499
rect 22477 2465 22511 2499
rect 24593 2465 24627 2499
rect 26341 2465 26375 2499
rect 28733 2465 28767 2499
rect 29009 2465 29043 2499
rect 31493 2465 31527 2499
rect 37473 2465 37507 2499
rect 37749 2465 37783 2499
rect 1593 2397 1627 2431
rect 3157 2397 3191 2431
rect 5549 2397 5583 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 10885 2397 10919 2431
rect 12633 2397 12667 2431
rect 16865 2397 16899 2431
rect 18061 2397 18095 2431
rect 19717 2397 19751 2431
rect 21189 2397 21223 2431
rect 32965 2397 32999 2431
rect 33609 2397 33643 2431
rect 34253 2397 34287 2431
rect 35081 2397 35115 2431
rect 36277 2397 36311 2431
rect 4077 2329 4111 2363
rect 8585 2329 8619 2363
rect 9229 2329 9263 2363
rect 13737 2329 13771 2363
rect 14381 2329 14415 2363
rect 20177 2329 20211 2363
rect 24869 2329 24903 2363
rect 31217 2329 31251 2363
rect 34161 2329 34195 2363
rect 2973 2261 3007 2295
rect 5365 2261 5399 2295
rect 7297 2261 7331 2295
rect 12449 2261 12483 2295
rect 17049 2261 17083 2295
rect 19533 2261 19567 2295
rect 21373 2261 21407 2295
rect 23949 2261 23983 2295
rect 32873 2261 32907 2295
rect 34989 2261 35023 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 16114 37408 16120 37460
rect 16172 37448 16178 37460
rect 16209 37451 16267 37457
rect 16209 37448 16221 37451
rect 16172 37420 16221 37448
rect 16172 37408 16178 37420
rect 16209 37417 16221 37420
rect 16255 37448 16267 37451
rect 26605 37451 26663 37457
rect 16255 37420 16574 37448
rect 16255 37417 16267 37420
rect 16209 37411 16267 37417
rect 9769 37315 9827 37321
rect 9769 37312 9781 37315
rect 9140 37284 9781 37312
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37213 1915 37247
rect 2314 37244 2320 37256
rect 2275 37216 2320 37244
rect 1857 37207 1915 37213
rect 1872 37176 1900 37207
rect 2314 37204 2320 37216
rect 2372 37204 2378 37256
rect 3418 37204 3424 37256
rect 3476 37244 3482 37256
rect 3973 37247 4031 37253
rect 3973 37244 3985 37247
rect 3476 37216 3985 37244
rect 3476 37204 3482 37216
rect 3973 37213 3985 37216
rect 4019 37213 4031 37247
rect 5534 37244 5540 37256
rect 5495 37216 5540 37244
rect 3973 37207 4031 37213
rect 5534 37204 5540 37216
rect 5592 37204 5598 37256
rect 7469 37247 7527 37253
rect 7469 37213 7481 37247
rect 7515 37244 7527 37247
rect 7515 37216 8064 37244
rect 7515 37213 7527 37216
rect 7469 37207 7527 37213
rect 2406 37176 2412 37188
rect 1872 37148 2412 37176
rect 2406 37136 2412 37148
rect 2464 37176 2470 37188
rect 3053 37179 3111 37185
rect 3053 37176 3065 37179
rect 2464 37148 3065 37176
rect 2464 37136 2470 37148
rect 3053 37145 3065 37148
rect 3099 37145 3111 37179
rect 3053 37139 3111 37145
rect 8036 37120 8064 37216
rect 9030 37204 9036 37256
rect 9088 37244 9094 37256
rect 9140 37253 9168 37284
rect 9769 37281 9781 37284
rect 9815 37281 9827 37315
rect 9769 37275 9827 37281
rect 10318 37272 10324 37324
rect 10376 37312 10382 37324
rect 11149 37315 11207 37321
rect 11149 37312 11161 37315
rect 10376 37284 11161 37312
rect 10376 37272 10382 37284
rect 11149 37281 11161 37284
rect 11195 37312 11207 37315
rect 11698 37312 11704 37324
rect 11195 37284 11704 37312
rect 11195 37281 11207 37284
rect 11149 37275 11207 37281
rect 11698 37272 11704 37284
rect 11756 37272 11762 37324
rect 11885 37315 11943 37321
rect 11885 37281 11897 37315
rect 11931 37312 11943 37315
rect 12250 37312 12256 37324
rect 11931 37284 12256 37312
rect 11931 37281 11943 37284
rect 11885 37275 11943 37281
rect 12250 37272 12256 37284
rect 12308 37312 12314 37324
rect 12345 37315 12403 37321
rect 12345 37312 12357 37315
rect 12308 37284 12357 37312
rect 12308 37272 12314 37284
rect 12345 37281 12357 37284
rect 12391 37281 12403 37315
rect 16546 37312 16574 37420
rect 26605 37417 26617 37451
rect 26651 37448 26663 37451
rect 27062 37448 27068 37460
rect 26651 37420 27068 37448
rect 26651 37417 26663 37420
rect 26605 37411 26663 37417
rect 27062 37408 27068 37420
rect 27120 37408 27126 37460
rect 34146 37408 34152 37460
rect 34204 37448 34210 37460
rect 34241 37451 34299 37457
rect 34241 37448 34253 37451
rect 34204 37420 34253 37448
rect 34204 37408 34210 37420
rect 34241 37417 34253 37420
rect 34287 37417 34299 37451
rect 34241 37411 34299 37417
rect 16853 37315 16911 37321
rect 16853 37312 16865 37315
rect 16546 37284 16865 37312
rect 12345 37275 12403 37281
rect 16853 37281 16865 37284
rect 16899 37281 16911 37315
rect 16853 37275 16911 37281
rect 19613 37315 19671 37321
rect 19613 37281 19625 37315
rect 19659 37312 19671 37315
rect 19978 37312 19984 37324
rect 19659 37284 19984 37312
rect 19659 37281 19671 37284
rect 19613 37275 19671 37281
rect 19978 37272 19984 37284
rect 20036 37312 20042 37324
rect 20073 37315 20131 37321
rect 20073 37312 20085 37315
rect 20036 37284 20085 37312
rect 20036 37272 20042 37284
rect 20073 37281 20085 37284
rect 20119 37281 20131 37315
rect 20073 37275 20131 37281
rect 23198 37272 23204 37324
rect 23256 37312 23262 37324
rect 24029 37315 24087 37321
rect 24029 37312 24041 37315
rect 23256 37284 24041 37312
rect 23256 37272 23262 37284
rect 24029 37281 24041 37284
rect 24075 37312 24087 37315
rect 24581 37315 24639 37321
rect 24581 37312 24593 37315
rect 24075 37284 24593 37312
rect 24075 37281 24087 37284
rect 24029 37275 24087 37281
rect 24581 37281 24593 37284
rect 24627 37281 24639 37315
rect 24581 37275 24639 37281
rect 26786 37272 26792 37324
rect 26844 37312 26850 37324
rect 27157 37315 27215 37321
rect 27157 37312 27169 37315
rect 26844 37284 27169 37312
rect 26844 37272 26850 37284
rect 27157 37281 27169 37284
rect 27203 37281 27215 37315
rect 34256 37312 34284 37411
rect 34256 37284 34560 37312
rect 27157 37275 27215 37281
rect 9125 37247 9183 37253
rect 9125 37244 9137 37247
rect 9088 37216 9137 37244
rect 9088 37204 9094 37216
rect 9125 37213 9137 37216
rect 9171 37213 9183 37247
rect 10870 37244 10876 37256
rect 10831 37216 10876 37244
rect 9125 37207 9183 37213
rect 10870 37204 10876 37216
rect 10928 37204 10934 37256
rect 12621 37247 12679 37253
rect 12621 37213 12633 37247
rect 12667 37213 12679 37247
rect 14274 37244 14280 37256
rect 14235 37216 14280 37244
rect 12621 37207 12679 37213
rect 12636 37176 12664 37207
rect 14274 37204 14280 37216
rect 14332 37204 14338 37256
rect 17126 37244 17132 37256
rect 17087 37216 17132 37244
rect 17126 37204 17132 37216
rect 17184 37204 17190 37256
rect 17862 37204 17868 37256
rect 17920 37244 17926 37256
rect 18141 37247 18199 37253
rect 18141 37244 18153 37247
rect 17920 37216 18153 37244
rect 17920 37204 17926 37216
rect 18141 37213 18153 37216
rect 18187 37213 18199 37247
rect 18141 37207 18199 37213
rect 20349 37247 20407 37253
rect 20349 37213 20361 37247
rect 20395 37244 20407 37247
rect 20395 37216 21312 37244
rect 20395 37213 20407 37216
rect 20349 37207 20407 37213
rect 20714 37176 20720 37188
rect 12636 37148 20720 37176
rect 20714 37136 20720 37148
rect 20772 37136 20778 37188
rect 21284 37176 21312 37216
rect 21358 37204 21364 37256
rect 21416 37244 21422 37256
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 21416 37216 22017 37244
rect 21416 37204 21422 37216
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 23753 37247 23811 37253
rect 23753 37213 23765 37247
rect 23799 37244 23811 37247
rect 25225 37247 25283 37253
rect 25225 37244 25237 37247
rect 23799 37216 24624 37244
rect 23799 37213 23811 37216
rect 23753 37207 23811 37213
rect 24596 37188 24624 37216
rect 24688 37216 25237 37244
rect 23382 37176 23388 37188
rect 21284 37148 23388 37176
rect 23382 37136 23388 37148
rect 23440 37136 23446 37188
rect 24578 37136 24584 37188
rect 24636 37136 24642 37188
rect 1302 37068 1308 37120
rect 1360 37108 1366 37120
rect 1673 37111 1731 37117
rect 1673 37108 1685 37111
rect 1360 37080 1685 37108
rect 1360 37068 1366 37080
rect 1673 37077 1685 37080
rect 1719 37077 1731 37111
rect 1673 37071 1731 37077
rect 2501 37111 2559 37117
rect 2501 37077 2513 37111
rect 2547 37108 2559 37111
rect 2774 37108 2780 37120
rect 2547 37080 2780 37108
rect 2547 37077 2559 37080
rect 2501 37071 2559 37077
rect 2774 37068 2780 37080
rect 2832 37068 2838 37120
rect 3234 37068 3240 37120
rect 3292 37108 3298 37120
rect 4157 37111 4215 37117
rect 4157 37108 4169 37111
rect 3292 37080 4169 37108
rect 3292 37068 3298 37080
rect 4157 37077 4169 37080
rect 4203 37077 4215 37111
rect 4157 37071 4215 37077
rect 5166 37068 5172 37120
rect 5224 37108 5230 37120
rect 5353 37111 5411 37117
rect 5353 37108 5365 37111
rect 5224 37080 5365 37108
rect 5224 37068 5230 37080
rect 5353 37077 5365 37080
rect 5399 37077 5411 37111
rect 5353 37071 5411 37077
rect 7098 37068 7104 37120
rect 7156 37108 7162 37120
rect 7285 37111 7343 37117
rect 7285 37108 7297 37111
rect 7156 37080 7297 37108
rect 7156 37068 7162 37080
rect 7285 37077 7297 37080
rect 7331 37077 7343 37111
rect 8018 37108 8024 37120
rect 7979 37080 8024 37108
rect 7285 37071 7343 37077
rect 8018 37068 8024 37080
rect 8076 37068 8082 37120
rect 9306 37108 9312 37120
rect 9267 37080 9312 37108
rect 9306 37068 9312 37080
rect 9364 37068 9370 37120
rect 14182 37068 14188 37120
rect 14240 37108 14246 37120
rect 14461 37111 14519 37117
rect 14461 37108 14473 37111
rect 14240 37080 14473 37108
rect 14240 37068 14246 37080
rect 14461 37077 14473 37080
rect 14507 37077 14519 37111
rect 14461 37071 14519 37077
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18325 37111 18383 37117
rect 18325 37108 18337 37111
rect 18104 37080 18337 37108
rect 18104 37068 18110 37080
rect 18325 37077 18337 37080
rect 18371 37077 18383 37111
rect 18325 37071 18383 37077
rect 21266 37068 21272 37120
rect 21324 37108 21330 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 21324 37080 22201 37108
rect 21324 37068 21330 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 23842 37068 23848 37120
rect 23900 37108 23906 37120
rect 24688 37108 24716 37216
rect 25225 37213 25237 37216
rect 25271 37213 25283 37247
rect 25225 37207 25283 37213
rect 27062 37204 27068 37256
rect 27120 37244 27126 37256
rect 27341 37247 27399 37253
rect 27341 37244 27353 37247
rect 27120 37216 27353 37244
rect 27120 37204 27126 37216
rect 27341 37213 27353 37216
rect 27387 37213 27399 37247
rect 27341 37207 27399 37213
rect 28718 37204 28724 37256
rect 28776 37244 28782 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 28776 37216 29745 37244
rect 28776 37204 28782 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 30466 37244 30472 37256
rect 30427 37216 30472 37244
rect 29733 37207 29791 37213
rect 30466 37204 30472 37216
rect 30524 37204 30530 37256
rect 32306 37244 32312 37256
rect 32267 37216 32312 37244
rect 32306 37204 32312 37216
rect 32364 37204 32370 37256
rect 34532 37244 34560 37284
rect 34790 37272 34796 37324
rect 34848 37312 34854 37324
rect 34885 37315 34943 37321
rect 34885 37312 34897 37315
rect 34848 37284 34897 37312
rect 34848 37272 34854 37284
rect 34885 37281 34897 37284
rect 34931 37281 34943 37315
rect 34885 37275 34943 37281
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34532 37216 35081 37244
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 36262 37204 36268 37256
rect 36320 37244 36326 37256
rect 36449 37247 36507 37253
rect 36449 37244 36461 37247
rect 36320 37216 36461 37244
rect 36320 37204 36326 37216
rect 36449 37213 36461 37216
rect 36495 37213 36507 37247
rect 36449 37207 36507 37213
rect 36906 37204 36912 37256
rect 36964 37244 36970 37256
rect 38013 37247 38071 37253
rect 38013 37244 38025 37247
rect 36964 37216 38025 37244
rect 36964 37204 36970 37216
rect 38013 37213 38025 37216
rect 38059 37213 38071 37247
rect 38013 37207 38071 37213
rect 23900 37080 24716 37108
rect 23900 37068 23906 37080
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25409 37111 25467 37117
rect 25409 37108 25421 37111
rect 25188 37080 25421 37108
rect 25188 37068 25194 37080
rect 25409 37077 25421 37080
rect 25455 37077 25467 37111
rect 25409 37071 25467 37077
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29052 37080 29929 37108
rect 29052 37068 29058 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 30374 37068 30380 37120
rect 30432 37108 30438 37120
rect 30653 37111 30711 37117
rect 30653 37108 30665 37111
rect 30432 37080 30665 37108
rect 30432 37068 30438 37080
rect 30653 37077 30665 37080
rect 30699 37077 30711 37111
rect 30653 37071 30711 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 36078 37068 36084 37120
rect 36136 37108 36142 37120
rect 36265 37111 36323 37117
rect 36265 37108 36277 37111
rect 36136 37080 36277 37108
rect 36136 37068 36142 37080
rect 36265 37077 36277 37080
rect 36311 37077 36323 37111
rect 36265 37071 36323 37077
rect 38010 37068 38016 37120
rect 38068 37108 38074 37120
rect 38197 37111 38255 37117
rect 38197 37108 38209 37111
rect 38068 37080 38209 37108
rect 38068 37068 38074 37080
rect 38197 37077 38209 37080
rect 38243 37077 38255 37111
rect 38197 37071 38255 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 3418 36904 3424 36916
rect 3379 36876 3424 36904
rect 3418 36864 3424 36876
rect 3476 36864 3482 36916
rect 11698 36904 11704 36916
rect 11659 36876 11704 36904
rect 11698 36864 11704 36876
rect 11756 36864 11762 36916
rect 17862 36904 17868 36916
rect 17823 36876 17868 36904
rect 17862 36864 17868 36876
rect 17920 36864 17926 36916
rect 20714 36904 20720 36916
rect 20675 36876 20720 36904
rect 20714 36864 20720 36876
rect 20772 36864 20778 36916
rect 21358 36904 21364 36916
rect 21319 36876 21364 36904
rect 21358 36864 21364 36876
rect 21416 36864 21422 36916
rect 30101 36907 30159 36913
rect 30101 36873 30113 36907
rect 30147 36904 30159 36907
rect 32306 36904 32312 36916
rect 30147 36876 32312 36904
rect 30147 36873 30159 36876
rect 30101 36867 30159 36873
rect 32306 36864 32312 36876
rect 32364 36864 32370 36916
rect 38197 36907 38255 36913
rect 38197 36873 38209 36907
rect 38243 36904 38255 36907
rect 39298 36904 39304 36916
rect 38243 36876 39304 36904
rect 38243 36873 38255 36876
rect 38197 36867 38255 36873
rect 39298 36864 39304 36876
rect 39356 36864 39362 36916
rect 14 36796 20 36848
rect 72 36836 78 36848
rect 1670 36836 1676 36848
rect 72 36808 1676 36836
rect 72 36796 78 36808
rect 1670 36796 1676 36808
rect 1728 36796 1734 36848
rect 3605 36771 3663 36777
rect 3605 36737 3617 36771
rect 3651 36768 3663 36771
rect 3651 36740 4200 36768
rect 3651 36737 3663 36740
rect 3605 36731 3663 36737
rect 1857 36635 1915 36641
rect 1857 36601 1869 36635
rect 1903 36632 1915 36635
rect 2222 36632 2228 36644
rect 1903 36604 2228 36632
rect 1903 36601 1915 36604
rect 1857 36595 1915 36601
rect 2222 36592 2228 36604
rect 2280 36592 2286 36644
rect 1486 36524 1492 36576
rect 1544 36564 1550 36576
rect 2314 36564 2320 36576
rect 1544 36536 2320 36564
rect 1544 36524 1550 36536
rect 2314 36524 2320 36536
rect 2372 36524 2378 36576
rect 4172 36573 4200 36740
rect 10870 36728 10876 36780
rect 10928 36768 10934 36780
rect 17678 36768 17684 36780
rect 10928 36740 17684 36768
rect 10928 36728 10934 36740
rect 17678 36728 17684 36740
rect 17736 36728 17742 36780
rect 20732 36768 20760 36864
rect 23382 36796 23388 36848
rect 23440 36836 23446 36848
rect 23440 36808 26234 36836
rect 23440 36796 23446 36808
rect 21177 36771 21235 36777
rect 21177 36768 21189 36771
rect 20732 36740 21189 36768
rect 21177 36737 21189 36740
rect 21223 36768 21235 36771
rect 22738 36768 22744 36780
rect 21223 36740 22744 36768
rect 21223 36737 21235 36740
rect 21177 36731 21235 36737
rect 22738 36728 22744 36740
rect 22796 36728 22802 36780
rect 24026 36768 24032 36780
rect 23939 36740 24032 36768
rect 24026 36728 24032 36740
rect 24084 36768 24090 36780
rect 24673 36771 24731 36777
rect 24673 36768 24685 36771
rect 24084 36740 24685 36768
rect 24084 36728 24090 36740
rect 24673 36737 24685 36740
rect 24719 36737 24731 36771
rect 24673 36731 24731 36737
rect 25961 36771 26019 36777
rect 25961 36737 25973 36771
rect 26007 36737 26019 36771
rect 26206 36768 26234 36808
rect 26418 36796 26424 36848
rect 26476 36836 26482 36848
rect 26476 36808 30052 36836
rect 26476 36796 26482 36808
rect 30024 36777 30052 36808
rect 27157 36771 27215 36777
rect 27157 36768 27169 36771
rect 26206 36740 27169 36768
rect 25961 36731 26019 36737
rect 27157 36737 27169 36740
rect 27203 36737 27215 36771
rect 27157 36731 27215 36737
rect 30009 36771 30067 36777
rect 30009 36737 30021 36771
rect 30055 36768 30067 36771
rect 30653 36771 30711 36777
rect 30653 36768 30665 36771
rect 30055 36740 30665 36768
rect 30055 36737 30067 36740
rect 30009 36731 30067 36737
rect 30653 36737 30665 36740
rect 30699 36737 30711 36771
rect 30653 36731 30711 36737
rect 38013 36771 38071 36777
rect 38013 36737 38025 36771
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 17126 36660 17132 36712
rect 17184 36700 17190 36712
rect 25409 36703 25467 36709
rect 25409 36700 25421 36703
rect 17184 36672 25421 36700
rect 17184 36660 17190 36672
rect 25409 36669 25421 36672
rect 25455 36700 25467 36703
rect 25976 36700 26004 36731
rect 26050 36700 26056 36712
rect 25455 36672 26056 36700
rect 25455 36669 25467 36672
rect 25409 36663 25467 36669
rect 26050 36660 26056 36672
rect 26108 36660 26114 36712
rect 36906 36700 36912 36712
rect 26160 36672 36912 36700
rect 26160 36641 26188 36672
rect 36906 36660 36912 36672
rect 36964 36660 36970 36712
rect 26145 36635 26203 36641
rect 26145 36601 26157 36635
rect 26191 36601 26203 36635
rect 26145 36595 26203 36601
rect 27341 36635 27399 36641
rect 27341 36601 27353 36635
rect 27387 36632 27399 36635
rect 38028 36632 38056 36731
rect 27387 36604 38056 36632
rect 27387 36601 27399 36604
rect 27341 36595 27399 36601
rect 4157 36567 4215 36573
rect 4157 36533 4169 36567
rect 4203 36564 4215 36567
rect 4798 36564 4804 36576
rect 4203 36536 4804 36564
rect 4203 36533 4215 36536
rect 4157 36527 4215 36533
rect 4798 36524 4804 36536
rect 4856 36524 4862 36576
rect 24210 36564 24216 36576
rect 24171 36536 24216 36564
rect 24210 36524 24216 36536
rect 24268 36524 24274 36576
rect 36262 36524 36268 36576
rect 36320 36564 36326 36576
rect 36541 36567 36599 36573
rect 36541 36564 36553 36567
rect 36320 36536 36553 36564
rect 36320 36524 36326 36536
rect 36541 36533 36553 36536
rect 36587 36533 36599 36567
rect 36541 36527 36599 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1670 36320 1676 36372
rect 1728 36360 1734 36372
rect 2317 36363 2375 36369
rect 2317 36360 2329 36363
rect 1728 36332 2329 36360
rect 1728 36320 1734 36332
rect 2317 36329 2329 36332
rect 2363 36329 2375 36363
rect 2317 36323 2375 36329
rect 24210 36320 24216 36372
rect 24268 36360 24274 36372
rect 30466 36360 30472 36372
rect 24268 36332 30472 36360
rect 24268 36320 24274 36332
rect 30466 36320 30472 36332
rect 30524 36320 30530 36372
rect 1854 36156 1860 36168
rect 1815 36128 1860 36156
rect 1854 36116 1860 36128
rect 1912 36116 1918 36168
rect 37734 36116 37740 36168
rect 37792 36156 37798 36168
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 37792 36128 38025 36156
rect 37792 36116 37798 36128
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 1670 36020 1676 36032
rect 1631 35992 1676 36020
rect 1670 35980 1676 35992
rect 1728 35980 1734 36032
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1854 35776 1860 35828
rect 1912 35816 1918 35828
rect 1949 35819 2007 35825
rect 1949 35816 1961 35819
rect 1912 35788 1961 35816
rect 1912 35776 1918 35788
rect 1949 35785 1961 35788
rect 1995 35785 2007 35819
rect 1949 35779 2007 35785
rect 38197 35819 38255 35825
rect 38197 35785 38209 35819
rect 38243 35816 38255 35819
rect 38286 35816 38292 35828
rect 38243 35788 38292 35816
rect 38243 35785 38255 35788
rect 38197 35779 38255 35785
rect 38286 35776 38292 35788
rect 38344 35776 38350 35828
rect 2041 35683 2099 35689
rect 2041 35649 2053 35683
rect 2087 35680 2099 35683
rect 2498 35680 2504 35692
rect 2087 35652 2504 35680
rect 2087 35649 2099 35652
rect 2041 35643 2099 35649
rect 2498 35640 2504 35652
rect 2556 35640 2562 35692
rect 37918 35640 37924 35692
rect 37976 35680 37982 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 37976 35652 38025 35680
rect 37976 35640 37982 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 2498 35476 2504 35488
rect 2459 35448 2504 35476
rect 2498 35436 2504 35448
rect 2556 35436 2562 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34592 1915 34595
rect 38013 34595 38071 34601
rect 38013 34592 38025 34595
rect 1903 34564 2176 34592
rect 1903 34561 1915 34564
rect 1857 34555 1915 34561
rect 2148 34536 2176 34564
rect 37476 34564 38025 34592
rect 37476 34536 37504 34564
rect 38013 34561 38025 34564
rect 38059 34561 38071 34595
rect 38013 34555 38071 34561
rect 2130 34484 2136 34536
rect 2188 34524 2194 34536
rect 2317 34527 2375 34533
rect 2317 34524 2329 34527
rect 2188 34496 2329 34524
rect 2188 34484 2194 34496
rect 2317 34493 2329 34496
rect 2363 34493 2375 34527
rect 37458 34524 37464 34536
rect 37419 34496 37464 34524
rect 2317 34487 2375 34493
rect 37458 34484 37464 34496
rect 37516 34484 37522 34536
rect 1670 34388 1676 34400
rect 1631 34360 1676 34388
rect 1670 34348 1676 34360
rect 1728 34348 1734 34400
rect 38194 34388 38200 34400
rect 38155 34360 38200 34388
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 1578 32376 1584 32428
rect 1636 32416 1642 32428
rect 1673 32419 1731 32425
rect 1673 32416 1685 32419
rect 1636 32388 1685 32416
rect 1636 32376 1642 32388
rect 1673 32385 1685 32388
rect 1719 32385 1731 32419
rect 25498 32416 25504 32428
rect 25459 32388 25504 32416
rect 1673 32379 1731 32385
rect 25498 32376 25504 32388
rect 25556 32416 25562 32428
rect 38013 32419 38071 32425
rect 38013 32416 38025 32419
rect 25556 32388 38025 32416
rect 25556 32376 25562 32388
rect 38013 32385 38025 32388
rect 38059 32385 38071 32419
rect 38013 32379 38071 32385
rect 38286 32348 38292 32360
rect 38247 32320 38292 32348
rect 38286 32308 38292 32320
rect 38344 32308 38350 32360
rect 1857 32283 1915 32289
rect 1857 32249 1869 32283
rect 1903 32280 1915 32283
rect 2682 32280 2688 32292
rect 1903 32252 2688 32280
rect 1903 32249 1915 32252
rect 1857 32243 1915 32249
rect 2682 32240 2688 32252
rect 2740 32240 2746 32292
rect 8018 32172 8024 32224
rect 8076 32212 8082 32224
rect 25409 32215 25467 32221
rect 25409 32212 25421 32215
rect 8076 32184 25421 32212
rect 8076 32172 8082 32184
rect 25409 32181 25421 32184
rect 25455 32181 25467 32215
rect 25409 32175 25467 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1578 32008 1584 32020
rect 1539 31980 1584 32008
rect 1578 31968 1584 31980
rect 1636 31968 1642 32020
rect 38286 32008 38292 32020
rect 38247 31980 38292 32008
rect 38286 31968 38292 31980
rect 38344 31968 38350 32020
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 23842 31464 23848 31476
rect 23803 31436 23848 31464
rect 23842 31424 23848 31436
rect 23900 31424 23906 31476
rect 23661 31331 23719 31337
rect 23661 31297 23673 31331
rect 23707 31328 23719 31331
rect 24302 31328 24308 31340
rect 23707 31300 24308 31328
rect 23707 31297 23719 31300
rect 23661 31291 23719 31297
rect 24302 31288 24308 31300
rect 24360 31288 24366 31340
rect 25498 31328 25504 31340
rect 25459 31300 25504 31328
rect 25498 31288 25504 31300
rect 25556 31288 25562 31340
rect 24302 31124 24308 31136
rect 24263 31096 24308 31124
rect 24302 31084 24308 31096
rect 24360 31084 24366 31136
rect 25130 31084 25136 31136
rect 25188 31124 25194 31136
rect 25409 31127 25467 31133
rect 25409 31124 25421 31127
rect 25188 31096 25421 31124
rect 25188 31084 25194 31096
rect 25409 31093 25421 31096
rect 25455 31093 25467 31127
rect 25409 31087 25467 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1857 30719 1915 30725
rect 1857 30685 1869 30719
rect 1903 30716 1915 30719
rect 1903 30688 2360 30716
rect 1903 30685 1915 30688
rect 1857 30679 1915 30685
rect 2332 30592 2360 30688
rect 9306 30676 9312 30728
rect 9364 30716 9370 30728
rect 10965 30719 11023 30725
rect 10965 30716 10977 30719
rect 9364 30688 10977 30716
rect 9364 30676 9370 30688
rect 10965 30685 10977 30688
rect 11011 30685 11023 30719
rect 10965 30679 11023 30685
rect 22925 30719 22983 30725
rect 22925 30685 22937 30719
rect 22971 30716 22983 30719
rect 23382 30716 23388 30728
rect 22971 30688 23388 30716
rect 22971 30685 22983 30688
rect 22925 30679 22983 30685
rect 23382 30676 23388 30688
rect 23440 30676 23446 30728
rect 11241 30651 11299 30657
rect 11241 30617 11253 30651
rect 11287 30648 11299 30651
rect 33686 30648 33692 30660
rect 11287 30620 33692 30648
rect 11287 30617 11299 30620
rect 11241 30611 11299 30617
rect 33686 30608 33692 30620
rect 33744 30608 33750 30660
rect 1670 30580 1676 30592
rect 1631 30552 1676 30580
rect 1670 30540 1676 30552
rect 1728 30540 1734 30592
rect 2314 30580 2320 30592
rect 2275 30552 2320 30580
rect 2314 30540 2320 30552
rect 2372 30540 2378 30592
rect 22922 30540 22928 30592
rect 22980 30580 22986 30592
rect 23017 30583 23075 30589
rect 23017 30580 23029 30583
rect 22980 30552 23029 30580
rect 22980 30540 22986 30552
rect 23017 30549 23029 30552
rect 23063 30549 23075 30583
rect 23017 30543 23075 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 17678 30200 17684 30252
rect 17736 30240 17742 30252
rect 18785 30243 18843 30249
rect 18785 30240 18797 30243
rect 17736 30212 18797 30240
rect 17736 30200 17742 30212
rect 18785 30209 18797 30212
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 25774 30132 25780 30184
rect 25832 30172 25838 30184
rect 38013 30175 38071 30181
rect 38013 30172 38025 30175
rect 25832 30144 38025 30172
rect 25832 30132 25838 30144
rect 38013 30141 38025 30144
rect 38059 30141 38071 30175
rect 38286 30172 38292 30184
rect 38247 30144 38292 30172
rect 38013 30135 38071 30141
rect 38286 30132 38292 30144
rect 38344 30132 38350 30184
rect 18877 30039 18935 30045
rect 18877 30005 18889 30039
rect 18923 30036 18935 30039
rect 20070 30036 20076 30048
rect 18923 30008 20076 30036
rect 18923 30005 18935 30008
rect 18877 29999 18935 30005
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 38286 29832 38292 29844
rect 38247 29804 38292 29832
rect 38286 29792 38292 29804
rect 38344 29792 38350 29844
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 14185 29291 14243 29297
rect 14185 29257 14197 29291
rect 14231 29288 14243 29291
rect 14274 29288 14280 29300
rect 14231 29260 14280 29288
rect 14231 29257 14243 29260
rect 14185 29251 14243 29257
rect 14274 29248 14280 29260
rect 14332 29248 14338 29300
rect 1854 29152 1860 29164
rect 1815 29124 1860 29152
rect 1854 29112 1860 29124
rect 1912 29112 1918 29164
rect 14001 29155 14059 29161
rect 14001 29121 14013 29155
rect 14047 29152 14059 29155
rect 22738 29152 22744 29164
rect 14047 29124 14780 29152
rect 22699 29124 22744 29152
rect 14047 29121 14059 29124
rect 14001 29115 14059 29121
rect 1670 29016 1676 29028
rect 1631 28988 1676 29016
rect 1670 28976 1676 28988
rect 1728 28976 1734 29028
rect 14752 29025 14780 29124
rect 22738 29112 22744 29124
rect 22796 29152 22802 29164
rect 23385 29155 23443 29161
rect 23385 29152 23397 29155
rect 22796 29124 23397 29152
rect 22796 29112 22802 29124
rect 23385 29121 23397 29124
rect 23431 29121 23443 29155
rect 38010 29152 38016 29164
rect 37971 29124 38016 29152
rect 23385 29115 23443 29121
rect 38010 29112 38016 29124
rect 38068 29112 38074 29164
rect 14737 29019 14795 29025
rect 14737 28985 14749 29019
rect 14783 29016 14795 29019
rect 16574 29016 16580 29028
rect 14783 28988 16580 29016
rect 14783 28985 14795 28988
rect 14737 28979 14795 28985
rect 16574 28976 16580 28988
rect 16632 28976 16638 29028
rect 22833 29019 22891 29025
rect 22833 28985 22845 29019
rect 22879 29016 22891 29019
rect 23198 29016 23204 29028
rect 22879 28988 23204 29016
rect 22879 28985 22891 28988
rect 22833 28979 22891 28985
rect 23198 28976 23204 28988
rect 23256 28976 23262 29028
rect 38194 29016 38200 29028
rect 38155 28988 38200 29016
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 2222 28500 2228 28552
rect 2280 28540 2286 28552
rect 23017 28543 23075 28549
rect 23017 28540 23029 28543
rect 2280 28512 23029 28540
rect 2280 28500 2286 28512
rect 23017 28509 23029 28512
rect 23063 28540 23075 28543
rect 23106 28540 23112 28552
rect 23063 28512 23112 28540
rect 23063 28509 23075 28512
rect 23017 28503 23075 28509
rect 23106 28500 23112 28512
rect 23164 28540 23170 28552
rect 23661 28543 23719 28549
rect 23661 28540 23673 28543
rect 23164 28512 23673 28540
rect 23164 28500 23170 28512
rect 23661 28509 23673 28512
rect 23707 28509 23719 28543
rect 23661 28503 23719 28509
rect 23216 28444 26234 28472
rect 23216 28413 23244 28444
rect 23201 28407 23259 28413
rect 23201 28373 23213 28407
rect 23247 28373 23259 28407
rect 26206 28404 26234 28444
rect 38010 28404 38016 28416
rect 26206 28376 38016 28404
rect 23201 28367 23259 28373
rect 38010 28364 38016 28376
rect 38068 28364 38074 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 23109 28203 23167 28209
rect 23109 28169 23121 28203
rect 23155 28200 23167 28203
rect 24026 28200 24032 28212
rect 23155 28172 24032 28200
rect 23155 28169 23167 28172
rect 23109 28163 23167 28169
rect 22557 28067 22615 28073
rect 22557 28064 22569 28067
rect 6886 28036 22569 28064
rect 2682 27820 2688 27872
rect 2740 27860 2746 27872
rect 6886 27860 6914 28036
rect 22557 28033 22569 28036
rect 22603 28064 22615 28067
rect 23124 28064 23152 28163
rect 24026 28160 24032 28172
rect 24084 28160 24090 28212
rect 26050 28160 26056 28212
rect 26108 28200 26114 28212
rect 26145 28203 26203 28209
rect 26145 28200 26157 28203
rect 26108 28172 26157 28200
rect 26108 28160 26114 28172
rect 26145 28169 26157 28172
rect 26191 28169 26203 28203
rect 26145 28163 26203 28169
rect 22603 28036 23152 28064
rect 25501 28067 25559 28073
rect 22603 28033 22615 28036
rect 22557 28027 22615 28033
rect 25501 28033 25513 28067
rect 25547 28064 25559 28067
rect 26068 28064 26096 28160
rect 25547 28036 26096 28064
rect 25547 28033 25559 28036
rect 25501 28027 25559 28033
rect 22462 27860 22468 27872
rect 2740 27832 6914 27860
rect 22423 27832 22468 27860
rect 2740 27820 2746 27832
rect 22462 27820 22468 27832
rect 22520 27820 22526 27872
rect 25593 27863 25651 27869
rect 25593 27829 25605 27863
rect 25639 27860 25651 27863
rect 25682 27860 25688 27872
rect 25639 27832 25688 27860
rect 25639 27829 25651 27832
rect 25593 27823 25651 27829
rect 25682 27820 25688 27832
rect 25740 27820 25746 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1578 26908 1584 26920
rect 1539 26880 1584 26908
rect 1578 26868 1584 26880
rect 1636 26868 1642 26920
rect 1857 26911 1915 26917
rect 1857 26877 1869 26911
rect 1903 26908 1915 26911
rect 2222 26908 2228 26920
rect 1903 26880 2228 26908
rect 1903 26877 1915 26880
rect 1857 26871 1915 26877
rect 2222 26868 2228 26880
rect 2280 26868 2286 26920
rect 38010 26908 38016 26920
rect 37971 26880 38016 26908
rect 38010 26868 38016 26880
rect 38068 26868 38074 26920
rect 38286 26908 38292 26920
rect 38247 26880 38292 26908
rect 38286 26868 38292 26880
rect 38344 26868 38350 26920
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1578 26568 1584 26580
rect 1539 26540 1584 26568
rect 1578 26528 1584 26540
rect 1636 26528 1642 26580
rect 23106 26568 23112 26580
rect 23067 26540 23112 26568
rect 23106 26528 23112 26540
rect 23164 26528 23170 26580
rect 38286 26568 38292 26580
rect 38247 26540 38292 26568
rect 38286 26528 38292 26540
rect 38344 26528 38350 26580
rect 16025 26503 16083 26509
rect 16025 26500 16037 26503
rect 6886 26472 16037 26500
rect 1854 26392 1860 26444
rect 1912 26432 1918 26444
rect 6886 26432 6914 26472
rect 16025 26469 16037 26472
rect 16071 26469 16083 26503
rect 16025 26463 16083 26469
rect 16761 26435 16819 26441
rect 16761 26432 16773 26435
rect 1912 26404 6914 26432
rect 16546 26404 16773 26432
rect 1912 26392 1918 26404
rect 16209 26367 16267 26373
rect 16209 26333 16221 26367
rect 16255 26364 16267 26367
rect 16546 26364 16574 26404
rect 16761 26401 16773 26404
rect 16807 26432 16819 26435
rect 24118 26432 24124 26444
rect 16807 26404 24124 26432
rect 16807 26401 16819 26404
rect 16761 26395 16819 26401
rect 24118 26392 24124 26404
rect 24176 26392 24182 26444
rect 16255 26336 16574 26364
rect 22465 26367 22523 26373
rect 16255 26333 16267 26336
rect 16209 26327 16267 26333
rect 22465 26333 22477 26367
rect 22511 26364 22523 26367
rect 23106 26364 23112 26376
rect 22511 26336 23112 26364
rect 22511 26333 22523 26336
rect 22465 26327 22523 26333
rect 23106 26324 23112 26336
rect 23164 26324 23170 26376
rect 22557 26299 22615 26305
rect 22557 26265 22569 26299
rect 22603 26296 22615 26299
rect 22646 26296 22652 26308
rect 22603 26268 22652 26296
rect 22603 26265 22615 26268
rect 22557 26259 22615 26265
rect 22646 26256 22652 26268
rect 22704 26256 22710 26308
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24800 1915 24803
rect 2038 24800 2044 24812
rect 1903 24772 2044 24800
rect 1903 24769 1915 24772
rect 1857 24763 1915 24769
rect 2038 24760 2044 24772
rect 2096 24760 2102 24812
rect 37553 24803 37611 24809
rect 37553 24769 37565 24803
rect 37599 24800 37611 24803
rect 38194 24800 38200 24812
rect 37599 24772 38200 24800
rect 37599 24769 37611 24772
rect 37553 24763 37611 24769
rect 38194 24760 38200 24772
rect 38252 24760 38258 24812
rect 38013 24667 38071 24673
rect 38013 24664 38025 24667
rect 26206 24636 38025 24664
rect 1670 24596 1676 24608
rect 1631 24568 1676 24596
rect 1670 24556 1676 24568
rect 1728 24556 1734 24608
rect 24118 24556 24124 24608
rect 24176 24596 24182 24608
rect 24762 24596 24768 24608
rect 24176 24568 24768 24596
rect 24176 24556 24182 24568
rect 24762 24556 24768 24568
rect 24820 24596 24826 24608
rect 26206 24596 26234 24636
rect 38013 24633 38025 24636
rect 38059 24633 38071 24667
rect 38013 24627 38071 24633
rect 24820 24568 26234 24596
rect 24820 24556 24826 24568
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 25774 24392 25780 24404
rect 25735 24364 25780 24392
rect 25774 24352 25780 24364
rect 25832 24352 25838 24404
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 4798 23808 4804 23860
rect 4856 23848 4862 23860
rect 28718 23848 28724 23860
rect 4856 23820 23888 23848
rect 28679 23820 28724 23848
rect 4856 23808 4862 23820
rect 23860 23789 23888 23820
rect 28718 23808 28724 23820
rect 28776 23808 28782 23860
rect 37458 23848 37464 23860
rect 35866 23820 37464 23848
rect 23845 23783 23903 23789
rect 23845 23749 23857 23783
rect 23891 23780 23903 23783
rect 24210 23780 24216 23792
rect 23891 23752 24216 23780
rect 23891 23749 23903 23752
rect 23845 23743 23903 23749
rect 24210 23740 24216 23752
rect 24268 23740 24274 23792
rect 24765 23783 24823 23789
rect 24765 23749 24777 23783
rect 24811 23780 24823 23783
rect 26237 23783 26295 23789
rect 26237 23780 26249 23783
rect 24811 23752 26249 23780
rect 24811 23749 24823 23752
rect 24765 23743 24823 23749
rect 26237 23749 26249 23752
rect 26283 23749 26295 23783
rect 35866 23780 35894 23820
rect 37458 23808 37464 23820
rect 37516 23808 37522 23860
rect 26237 23743 26295 23749
rect 27172 23752 35894 23780
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23712 22431 23715
rect 22462 23712 22468 23724
rect 22419 23684 22468 23712
rect 22419 23681 22431 23684
rect 22373 23675 22431 23681
rect 22462 23672 22468 23684
rect 22520 23672 22526 23724
rect 23017 23715 23075 23721
rect 23017 23681 23029 23715
rect 23063 23712 23075 23715
rect 23290 23712 23296 23724
rect 23063 23684 23296 23712
rect 23063 23681 23075 23684
rect 23017 23675 23075 23681
rect 23290 23672 23296 23684
rect 23348 23712 23354 23724
rect 25593 23715 25651 23721
rect 23348 23684 23980 23712
rect 23348 23672 23354 23684
rect 22554 23644 22560 23656
rect 22515 23616 22560 23644
rect 22554 23604 22560 23616
rect 22612 23604 22618 23656
rect 23952 23644 23980 23684
rect 25593 23681 25605 23715
rect 25639 23712 25651 23715
rect 25774 23712 25780 23724
rect 25639 23684 25780 23712
rect 25639 23681 25651 23684
rect 25593 23675 25651 23681
rect 25774 23672 25780 23684
rect 25832 23672 25838 23724
rect 26326 23712 26332 23724
rect 26287 23684 26332 23712
rect 26326 23672 26332 23684
rect 26384 23712 26390 23724
rect 27172 23721 27200 23752
rect 27157 23715 27215 23721
rect 27157 23712 27169 23715
rect 26384 23684 27169 23712
rect 26384 23672 26390 23684
rect 27157 23681 27169 23684
rect 27203 23681 27215 23715
rect 27157 23675 27215 23681
rect 28074 23672 28080 23724
rect 28132 23712 28138 23724
rect 28537 23715 28595 23721
rect 28537 23712 28549 23715
rect 28132 23684 28549 23712
rect 28132 23672 28138 23684
rect 28537 23681 28549 23684
rect 28583 23712 28595 23715
rect 29181 23715 29239 23721
rect 29181 23712 29193 23715
rect 28583 23684 29193 23712
rect 28583 23681 28595 23684
rect 28537 23675 28595 23681
rect 29181 23681 29193 23684
rect 29227 23681 29239 23715
rect 29181 23675 29239 23681
rect 24857 23647 24915 23653
rect 24857 23644 24869 23647
rect 23952 23616 24869 23644
rect 24857 23613 24869 23616
rect 24903 23613 24915 23647
rect 24857 23607 24915 23613
rect 7466 23536 7472 23588
rect 7524 23576 7530 23588
rect 25409 23579 25467 23585
rect 25409 23576 25421 23579
rect 7524 23548 25421 23576
rect 7524 23536 7530 23548
rect 25409 23545 25421 23548
rect 25455 23545 25467 23579
rect 25409 23539 25467 23545
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 5534 23264 5540 23316
rect 5592 23304 5598 23316
rect 7285 23307 7343 23313
rect 7285 23304 7297 23307
rect 5592 23276 7297 23304
rect 5592 23264 5598 23276
rect 7285 23273 7297 23276
rect 7331 23273 7343 23307
rect 23290 23304 23296 23316
rect 23251 23276 23296 23304
rect 7285 23267 7343 23273
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 25774 23264 25780 23316
rect 25832 23304 25838 23316
rect 25961 23307 26019 23313
rect 25961 23304 25973 23307
rect 25832 23276 25973 23304
rect 25832 23264 25838 23276
rect 25961 23273 25973 23276
rect 26007 23273 26019 23307
rect 25961 23267 26019 23273
rect 22646 23168 22652 23180
rect 22607 23140 22652 23168
rect 22646 23128 22652 23140
rect 22704 23128 22710 23180
rect 7469 23103 7527 23109
rect 7469 23069 7481 23103
rect 7515 23100 7527 23103
rect 22830 23100 22836 23112
rect 7515 23072 8064 23100
rect 22791 23072 22836 23100
rect 7515 23069 7527 23072
rect 7469 23063 7527 23069
rect 1670 22964 1676 22976
rect 1631 22936 1676 22964
rect 1670 22924 1676 22936
rect 1728 22924 1734 22976
rect 8036 22973 8064 23072
rect 22830 23060 22836 23072
rect 22888 23060 22894 23112
rect 25501 23103 25559 23109
rect 25501 23069 25513 23103
rect 25547 23100 25559 23103
rect 25774 23100 25780 23112
rect 25547 23072 25780 23100
rect 25547 23069 25559 23072
rect 25501 23063 25559 23069
rect 25774 23060 25780 23072
rect 25832 23060 25838 23112
rect 8021 22967 8079 22973
rect 8021 22933 8033 22967
rect 8067 22964 8079 22967
rect 12066 22964 12072 22976
rect 8067 22936 12072 22964
rect 8067 22933 8079 22936
rect 8021 22927 8079 22933
rect 12066 22924 12072 22936
rect 12124 22924 12130 22976
rect 25409 22967 25467 22973
rect 25409 22933 25421 22967
rect 25455 22964 25467 22967
rect 25498 22964 25504 22976
rect 25455 22936 25504 22964
rect 25455 22933 25467 22936
rect 25409 22927 25467 22933
rect 25498 22924 25504 22936
rect 25556 22924 25562 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 25406 22692 25412 22704
rect 25367 22664 25412 22692
rect 25406 22652 25412 22664
rect 25464 22652 25470 22704
rect 25498 22652 25504 22704
rect 25556 22692 25562 22704
rect 25556 22664 25601 22692
rect 25556 22652 25562 22664
rect 1670 22624 1676 22636
rect 1631 22596 1676 22624
rect 1670 22584 1676 22596
rect 1728 22584 1734 22636
rect 35710 22584 35716 22636
rect 35768 22624 35774 22636
rect 38013 22627 38071 22633
rect 38013 22624 38025 22627
rect 35768 22596 38025 22624
rect 35768 22584 35774 22596
rect 38013 22593 38025 22596
rect 38059 22593 38071 22627
rect 38013 22587 38071 22593
rect 23014 22556 23020 22568
rect 22975 22528 23020 22556
rect 23014 22516 23020 22528
rect 23072 22516 23078 22568
rect 1854 22488 1860 22500
rect 1815 22460 1860 22488
rect 1854 22448 1860 22460
rect 1912 22448 1918 22500
rect 24946 22488 24952 22500
rect 24907 22460 24952 22488
rect 24946 22448 24952 22460
rect 25004 22448 25010 22500
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 22373 22219 22431 22225
rect 22373 22185 22385 22219
rect 22419 22216 22431 22219
rect 22830 22216 22836 22228
rect 22419 22188 22836 22216
rect 22419 22185 22431 22188
rect 22373 22179 22431 22185
rect 22830 22176 22836 22188
rect 22888 22176 22894 22228
rect 23290 22216 23296 22228
rect 23251 22188 23296 22216
rect 23290 22176 23296 22188
rect 23348 22176 23354 22228
rect 25041 22219 25099 22225
rect 25041 22185 25053 22219
rect 25087 22216 25099 22219
rect 25406 22216 25412 22228
rect 25087 22188 25412 22216
rect 25087 22185 25099 22188
rect 25041 22179 25099 22185
rect 25406 22176 25412 22188
rect 25464 22176 25470 22228
rect 22925 22083 22983 22089
rect 22925 22049 22937 22083
rect 22971 22080 22983 22083
rect 23014 22080 23020 22092
rect 22971 22052 23020 22080
rect 22971 22049 22983 22052
rect 22925 22043 22983 22049
rect 23014 22040 23020 22052
rect 23072 22040 23078 22092
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 22012 2283 22015
rect 21821 22015 21879 22021
rect 2271 21984 2820 22012
rect 2271 21981 2283 21984
rect 2225 21975 2283 21981
rect 2038 21876 2044 21888
rect 1999 21848 2044 21876
rect 2038 21836 2044 21848
rect 2096 21836 2102 21888
rect 2792 21885 2820 21984
rect 21821 21981 21833 22015
rect 21867 22012 21879 22015
rect 22278 22012 22284 22024
rect 21867 21984 22284 22012
rect 21867 21981 21879 21984
rect 21821 21975 21879 21981
rect 22278 21972 22284 21984
rect 22336 21972 22342 22024
rect 23106 22012 23112 22024
rect 23067 21984 23112 22012
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 24026 21972 24032 22024
rect 24084 22012 24090 22024
rect 24949 22015 25007 22021
rect 24949 22012 24961 22015
rect 24084 21984 24961 22012
rect 24084 21972 24090 21984
rect 24949 21981 24961 21984
rect 24995 22012 25007 22015
rect 25593 22015 25651 22021
rect 25593 22012 25605 22015
rect 24995 21984 25605 22012
rect 24995 21981 25007 21984
rect 24949 21975 25007 21981
rect 25593 21981 25605 21984
rect 25639 21981 25651 22015
rect 25593 21975 25651 21981
rect 2777 21879 2835 21885
rect 2777 21845 2789 21879
rect 2823 21876 2835 21879
rect 10134 21876 10140 21888
rect 2823 21848 10140 21876
rect 2823 21845 2835 21848
rect 2777 21839 2835 21845
rect 10134 21836 10140 21848
rect 10192 21836 10198 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 22465 21675 22523 21681
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 22554 21672 22560 21684
rect 22511 21644 22560 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 23106 21672 23112 21684
rect 23067 21644 23112 21672
rect 23106 21632 23112 21644
rect 23164 21632 23170 21684
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21536 22431 21539
rect 22738 21536 22744 21548
rect 22419 21508 22744 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 22738 21496 22744 21508
rect 22796 21496 22802 21548
rect 23201 21539 23259 21545
rect 23201 21505 23213 21539
rect 23247 21536 23259 21539
rect 24026 21536 24032 21548
rect 23247 21508 24032 21536
rect 23247 21505 23259 21508
rect 23201 21499 23259 21505
rect 24026 21496 24032 21508
rect 24084 21496 24090 21548
rect 24121 21539 24179 21545
rect 24121 21505 24133 21539
rect 24167 21536 24179 21539
rect 24780 21536 24808 21632
rect 24167 21508 24808 21536
rect 24167 21505 24179 21508
rect 24121 21499 24179 21505
rect 24213 21335 24271 21341
rect 24213 21301 24225 21335
rect 24259 21332 24271 21335
rect 24578 21332 24584 21344
rect 24259 21304 24584 21332
rect 24259 21301 24271 21304
rect 24213 21295 24271 21301
rect 24578 21292 24584 21304
rect 24636 21292 24642 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 30285 21063 30343 21069
rect 30285 21029 30297 21063
rect 30331 21060 30343 21063
rect 30331 21032 35894 21060
rect 30331 21029 30343 21032
rect 30285 21023 30343 21029
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20924 23535 20927
rect 24486 20924 24492 20936
rect 23523 20896 24492 20924
rect 23523 20893 23535 20896
rect 23477 20887 23535 20893
rect 24486 20884 24492 20896
rect 24544 20924 24550 20936
rect 24673 20927 24731 20933
rect 24673 20924 24685 20927
rect 24544 20896 24685 20924
rect 24544 20884 24550 20896
rect 24673 20893 24685 20896
rect 24719 20924 24731 20927
rect 30101 20927 30159 20933
rect 30101 20924 30113 20927
rect 24719 20896 30113 20924
rect 24719 20893 24731 20896
rect 24673 20887 24731 20893
rect 30101 20893 30113 20896
rect 30147 20924 30159 20927
rect 30745 20927 30803 20933
rect 30745 20924 30757 20927
rect 30147 20896 30757 20924
rect 30147 20893 30159 20896
rect 30101 20887 30159 20893
rect 30745 20893 30757 20896
rect 30791 20893 30803 20927
rect 35866 20924 35894 21032
rect 38013 20927 38071 20933
rect 38013 20924 38025 20927
rect 35866 20896 38025 20924
rect 30745 20887 30803 20893
rect 38013 20893 38025 20896
rect 38059 20893 38071 20927
rect 38013 20887 38071 20893
rect 1578 20816 1584 20868
rect 1636 20856 1642 20868
rect 1673 20859 1731 20865
rect 1673 20856 1685 20859
rect 1636 20828 1685 20856
rect 1636 20816 1642 20828
rect 1673 20825 1685 20828
rect 1719 20825 1731 20859
rect 1673 20819 1731 20825
rect 1857 20859 1915 20865
rect 1857 20825 1869 20859
rect 1903 20856 1915 20859
rect 16574 20856 16580 20868
rect 1903 20828 16580 20856
rect 1903 20825 1915 20828
rect 1857 20819 1915 20825
rect 16574 20816 16580 20828
rect 16632 20816 16638 20868
rect 19797 20859 19855 20865
rect 19797 20825 19809 20859
rect 19843 20856 19855 20859
rect 19978 20856 19984 20868
rect 19843 20828 19984 20856
rect 19843 20825 19855 20828
rect 19797 20819 19855 20825
rect 19978 20816 19984 20828
rect 20036 20856 20042 20868
rect 20349 20859 20407 20865
rect 20349 20856 20361 20859
rect 20036 20828 20361 20856
rect 20036 20816 20042 20828
rect 20349 20825 20361 20828
rect 20395 20825 20407 20859
rect 20349 20819 20407 20825
rect 2314 20748 2320 20800
rect 2372 20788 2378 20800
rect 19705 20791 19763 20797
rect 19705 20788 19717 20791
rect 2372 20760 19717 20788
rect 2372 20748 2378 20760
rect 19705 20757 19717 20760
rect 19751 20757 19763 20791
rect 22738 20788 22744 20800
rect 22699 20760 22744 20788
rect 19705 20751 19763 20757
rect 22738 20748 22744 20760
rect 22796 20748 22802 20800
rect 23382 20788 23388 20800
rect 23343 20760 23388 20788
rect 23382 20748 23388 20760
rect 23440 20748 23446 20800
rect 24026 20788 24032 20800
rect 23939 20760 24032 20788
rect 24026 20748 24032 20760
rect 24084 20788 24090 20800
rect 24394 20788 24400 20800
rect 24084 20760 24400 20788
rect 24084 20748 24090 20760
rect 24394 20748 24400 20760
rect 24452 20748 24458 20800
rect 38194 20788 38200 20800
rect 38155 20760 38200 20788
rect 38194 20748 38200 20760
rect 38252 20748 38258 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 22189 20587 22247 20593
rect 22189 20584 22201 20587
rect 6886 20556 22201 20584
rect 1578 20516 1584 20528
rect 1539 20488 1584 20516
rect 1578 20476 1584 20488
rect 1636 20476 1642 20528
rect 1854 20204 1860 20256
rect 1912 20244 1918 20256
rect 6886 20244 6914 20556
rect 22189 20553 22201 20556
rect 22235 20584 22247 20587
rect 24302 20584 24308 20596
rect 22235 20556 24308 20584
rect 22235 20553 22247 20556
rect 22189 20547 22247 20553
rect 22664 20457 22692 20556
rect 24302 20544 24308 20556
rect 24360 20544 24366 20596
rect 37918 20544 37924 20596
rect 37976 20584 37982 20596
rect 38013 20587 38071 20593
rect 38013 20584 38025 20587
rect 37976 20556 38025 20584
rect 37976 20544 37982 20556
rect 38013 20553 38025 20556
rect 38059 20553 38071 20587
rect 38013 20547 38071 20553
rect 23477 20519 23535 20525
rect 23477 20485 23489 20519
rect 23523 20516 23535 20519
rect 23658 20516 23664 20528
rect 23523 20488 23664 20516
rect 23523 20485 23535 20488
rect 23477 20479 23535 20485
rect 23658 20476 23664 20488
rect 23716 20476 23722 20528
rect 25314 20516 25320 20528
rect 25275 20488 25320 20516
rect 25314 20476 25320 20488
rect 25372 20476 25378 20528
rect 22649 20451 22707 20457
rect 22649 20417 22661 20451
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 27341 20451 27399 20457
rect 27341 20417 27353 20451
rect 27387 20448 27399 20451
rect 37826 20448 37832 20460
rect 27387 20420 27936 20448
rect 37787 20420 37832 20448
rect 27387 20417 27399 20420
rect 27341 20411 27399 20417
rect 23382 20380 23388 20392
rect 23343 20352 23388 20380
rect 23382 20340 23388 20352
rect 23440 20340 23446 20392
rect 24029 20383 24087 20389
rect 24029 20349 24041 20383
rect 24075 20380 24087 20383
rect 24946 20380 24952 20392
rect 24075 20352 24952 20380
rect 24075 20349 24087 20352
rect 24029 20343 24087 20349
rect 24946 20340 24952 20352
rect 25004 20380 25010 20392
rect 25222 20380 25228 20392
rect 25004 20352 25228 20380
rect 25004 20340 25010 20352
rect 25222 20340 25228 20352
rect 25280 20340 25286 20392
rect 25409 20383 25467 20389
rect 25409 20349 25421 20383
rect 25455 20380 25467 20383
rect 25455 20352 26464 20380
rect 25455 20349 25467 20352
rect 25409 20343 25467 20349
rect 26436 20256 26464 20352
rect 1912 20216 6914 20244
rect 22741 20247 22799 20253
rect 1912 20204 1918 20216
rect 22741 20213 22753 20247
rect 22787 20244 22799 20247
rect 23750 20244 23756 20256
rect 22787 20216 23756 20244
rect 22787 20213 22799 20216
rect 22741 20207 22799 20213
rect 23750 20204 23756 20216
rect 23808 20204 23814 20256
rect 26418 20204 26424 20256
rect 26476 20244 26482 20256
rect 27908 20253 27936 20420
rect 37826 20408 37832 20420
rect 37884 20408 37890 20460
rect 27249 20247 27307 20253
rect 27249 20244 27261 20247
rect 26476 20216 27261 20244
rect 26476 20204 26482 20216
rect 27249 20213 27261 20216
rect 27295 20213 27307 20247
rect 27249 20207 27307 20213
rect 27893 20247 27951 20253
rect 27893 20213 27905 20247
rect 27939 20244 27951 20247
rect 28074 20244 28080 20256
rect 27939 20216 28080 20244
rect 27939 20213 27951 20216
rect 27893 20207 27951 20213
rect 28074 20204 28080 20216
rect 28132 20204 28138 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 23658 20040 23664 20052
rect 23619 20012 23664 20040
rect 23658 20000 23664 20012
rect 23716 20000 23722 20052
rect 24857 20043 24915 20049
rect 24857 20009 24869 20043
rect 24903 20040 24915 20043
rect 25314 20040 25320 20052
rect 24903 20012 25320 20040
rect 24903 20009 24915 20012
rect 24857 20003 24915 20009
rect 25314 20000 25320 20012
rect 25372 20000 25378 20052
rect 2130 19932 2136 19984
rect 2188 19972 2194 19984
rect 9125 19975 9183 19981
rect 9125 19972 9137 19975
rect 2188 19944 9137 19972
rect 2188 19932 2194 19944
rect 9125 19941 9137 19944
rect 9171 19941 9183 19975
rect 9125 19935 9183 19941
rect 22278 19864 22284 19916
rect 22336 19904 22342 19916
rect 22336 19876 24808 19904
rect 22336 19864 22342 19876
rect 16574 19796 16580 19848
rect 16632 19836 16638 19848
rect 17221 19839 17279 19845
rect 17221 19836 17233 19839
rect 16632 19808 17233 19836
rect 16632 19796 16638 19808
rect 17221 19805 17233 19808
rect 17267 19805 17279 19839
rect 22462 19836 22468 19848
rect 22423 19808 22468 19836
rect 17221 19799 17279 19805
rect 22462 19796 22468 19808
rect 22520 19796 22526 19848
rect 22649 19839 22707 19845
rect 22649 19805 22661 19839
rect 22695 19836 22707 19839
rect 23290 19836 23296 19848
rect 22695 19808 23296 19836
rect 22695 19805 22707 19808
rect 22649 19799 22707 19805
rect 23290 19796 23296 19808
rect 23348 19796 23354 19848
rect 23658 19796 23664 19848
rect 23716 19836 23722 19848
rect 24780 19845 24808 19876
rect 23753 19839 23811 19845
rect 23753 19836 23765 19839
rect 23716 19808 23765 19836
rect 23716 19796 23722 19808
rect 23753 19805 23765 19808
rect 23799 19805 23811 19839
rect 23753 19799 23811 19805
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19836 24823 19839
rect 24811 19808 25544 19836
rect 24811 19805 24823 19808
rect 24765 19799 24823 19805
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19737 9367 19771
rect 9309 19731 9367 19737
rect 16669 19771 16727 19777
rect 16669 19737 16681 19771
rect 16715 19768 16727 19771
rect 19242 19768 19248 19780
rect 16715 19740 19248 19768
rect 16715 19737 16727 19740
rect 16669 19731 16727 19737
rect 9324 19700 9352 19731
rect 19242 19728 19248 19740
rect 19300 19728 19306 19780
rect 22005 19771 22063 19777
rect 22005 19737 22017 19771
rect 22051 19768 22063 19771
rect 22738 19768 22744 19780
rect 22051 19740 22744 19768
rect 22051 19737 22063 19740
rect 22005 19731 22063 19737
rect 22738 19728 22744 19740
rect 22796 19768 22802 19780
rect 23676 19768 23704 19796
rect 25409 19771 25467 19777
rect 25409 19768 25421 19771
rect 22796 19740 25421 19768
rect 22796 19728 22802 19740
rect 25409 19737 25421 19740
rect 25455 19737 25467 19771
rect 25409 19731 25467 19737
rect 25516 19712 25544 19808
rect 9858 19700 9864 19712
rect 9324 19672 9864 19700
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 23109 19703 23167 19709
rect 23109 19669 23121 19703
rect 23155 19700 23167 19703
rect 23474 19700 23480 19712
rect 23155 19672 23480 19700
rect 23155 19669 23167 19672
rect 23109 19663 23167 19669
rect 23474 19660 23480 19672
rect 23532 19660 23538 19712
rect 25498 19660 25504 19712
rect 25556 19700 25562 19712
rect 25961 19703 26019 19709
rect 25961 19700 25973 19703
rect 25556 19672 25973 19700
rect 25556 19660 25562 19672
rect 25961 19669 25973 19672
rect 26007 19669 26019 19703
rect 25961 19663 26019 19669
rect 37274 19660 37280 19712
rect 37332 19700 37338 19712
rect 37645 19703 37703 19709
rect 37645 19700 37657 19703
rect 37332 19672 37657 19700
rect 37332 19660 37338 19672
rect 37645 19669 37657 19672
rect 37691 19700 37703 19703
rect 37826 19700 37832 19712
rect 37691 19672 37832 19700
rect 37691 19669 37703 19672
rect 37645 19663 37703 19669
rect 37826 19660 37832 19672
rect 37884 19660 37890 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 23290 19496 23296 19508
rect 23251 19468 23296 19496
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 26878 19496 26884 19508
rect 25148 19468 26884 19496
rect 22186 19428 22192 19440
rect 22147 19400 22192 19428
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 24210 19428 24216 19440
rect 24171 19400 24216 19428
rect 24210 19388 24216 19400
rect 24268 19388 24274 19440
rect 25148 19437 25176 19468
rect 26878 19456 26884 19468
rect 26936 19456 26942 19508
rect 25133 19431 25191 19437
rect 25133 19397 25145 19431
rect 25179 19397 25191 19431
rect 25133 19391 25191 19397
rect 25222 19388 25228 19440
rect 25280 19428 25286 19440
rect 26326 19428 26332 19440
rect 25280 19400 25325 19428
rect 26287 19400 26332 19428
rect 25280 19388 25286 19400
rect 26326 19388 26332 19400
rect 26384 19388 26390 19440
rect 26418 19388 26424 19440
rect 26476 19428 26482 19440
rect 26476 19400 26521 19428
rect 26476 19388 26482 19400
rect 1857 19363 1915 19369
rect 1857 19329 1869 19363
rect 1903 19360 1915 19363
rect 15746 19360 15752 19372
rect 1903 19332 15752 19360
rect 1903 19329 1915 19332
rect 1857 19323 1915 19329
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 23385 19363 23443 19369
rect 20128 19332 21956 19360
rect 20128 19320 20134 19332
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 21928 19292 21956 19332
rect 23385 19329 23397 19363
rect 23431 19360 23443 19363
rect 23658 19360 23664 19372
rect 23431 19332 23664 19360
rect 23431 19329 23443 19332
rect 23385 19323 23443 19329
rect 23658 19320 23664 19332
rect 23716 19320 23722 19372
rect 33134 19320 33140 19372
rect 33192 19360 33198 19372
rect 38013 19363 38071 19369
rect 38013 19360 38025 19363
rect 33192 19332 38025 19360
rect 33192 19320 33198 19332
rect 38013 19329 38025 19332
rect 38059 19329 38071 19363
rect 38013 19323 38071 19329
rect 22097 19295 22155 19301
rect 22097 19292 22109 19295
rect 21928 19264 22109 19292
rect 22097 19261 22109 19264
rect 22143 19261 22155 19295
rect 22097 19255 22155 19261
rect 22278 19184 22284 19236
rect 22336 19224 22342 19236
rect 22649 19227 22707 19233
rect 22649 19224 22661 19227
rect 22336 19196 22661 19224
rect 22336 19184 22342 19196
rect 22649 19193 22661 19196
rect 22695 19224 22707 19227
rect 25406 19224 25412 19236
rect 22695 19196 25412 19224
rect 22695 19193 22707 19196
rect 22649 19187 22707 19193
rect 25406 19184 25412 19196
rect 25464 19224 25470 19236
rect 25869 19227 25927 19233
rect 25869 19224 25881 19227
rect 25464 19196 25881 19224
rect 25464 19184 25470 19196
rect 25869 19193 25881 19196
rect 25915 19193 25927 19227
rect 25869 19187 25927 19193
rect 38194 19156 38200 19168
rect 38155 19128 38200 19156
rect 38194 19116 38200 19128
rect 38252 19116 38258 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 25961 18955 26019 18961
rect 25961 18921 25973 18955
rect 26007 18952 26019 18955
rect 26326 18952 26332 18964
rect 26007 18924 26332 18952
rect 26007 18921 26019 18924
rect 25961 18915 26019 18921
rect 26326 18912 26332 18924
rect 26384 18912 26390 18964
rect 37734 18912 37740 18964
rect 37792 18952 37798 18964
rect 38013 18955 38071 18961
rect 38013 18952 38025 18955
rect 37792 18924 38025 18952
rect 37792 18912 37798 18924
rect 38013 18921 38025 18924
rect 38059 18921 38071 18955
rect 38013 18915 38071 18921
rect 10321 18887 10379 18893
rect 10321 18853 10333 18887
rect 10367 18884 10379 18887
rect 22462 18884 22468 18896
rect 10367 18856 22468 18884
rect 10367 18853 10379 18856
rect 10321 18847 10379 18853
rect 22462 18844 22468 18856
rect 22520 18844 22526 18896
rect 22554 18844 22560 18896
rect 22612 18884 22618 18896
rect 22612 18856 24808 18884
rect 22612 18844 22618 18856
rect 19242 18776 19248 18828
rect 19300 18816 19306 18828
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 19300 18788 21649 18816
rect 19300 18776 19306 18788
rect 21637 18785 21649 18788
rect 21683 18785 21695 18819
rect 22278 18816 22284 18828
rect 22239 18788 22284 18816
rect 21637 18779 21695 18785
rect 22278 18776 22284 18788
rect 22336 18776 22342 18828
rect 22922 18776 22928 18828
rect 22980 18816 22986 18828
rect 23109 18819 23167 18825
rect 23109 18816 23121 18819
rect 22980 18788 23121 18816
rect 22980 18776 22986 18788
rect 23109 18785 23121 18788
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 23198 18776 23204 18828
rect 23256 18816 23262 18828
rect 23385 18819 23443 18825
rect 23385 18816 23397 18819
rect 23256 18788 23397 18816
rect 23256 18776 23262 18788
rect 23385 18785 23397 18788
rect 23431 18785 23443 18819
rect 23385 18779 23443 18785
rect 24780 18816 24808 18856
rect 24780 18788 25912 18816
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 24780 18757 24808 18788
rect 10229 18751 10287 18757
rect 10229 18748 10241 18751
rect 2280 18720 10241 18748
rect 2280 18708 2286 18720
rect 10229 18717 10241 18720
rect 10275 18748 10287 18751
rect 10873 18751 10931 18757
rect 10873 18748 10885 18751
rect 10275 18720 10885 18748
rect 10275 18717 10287 18720
rect 10229 18711 10287 18717
rect 10873 18717 10885 18720
rect 10919 18717 10931 18751
rect 10873 18711 10931 18717
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 25409 18751 25467 18757
rect 25409 18717 25421 18751
rect 25455 18748 25467 18751
rect 25498 18748 25504 18760
rect 25455 18720 25504 18748
rect 25455 18717 25467 18720
rect 25409 18711 25467 18717
rect 25498 18708 25504 18720
rect 25556 18708 25562 18760
rect 25884 18757 25912 18788
rect 25869 18751 25927 18757
rect 25869 18717 25881 18751
rect 25915 18748 25927 18751
rect 26513 18751 26571 18757
rect 26513 18748 26525 18751
rect 25915 18720 26525 18748
rect 25915 18717 25927 18720
rect 25869 18711 25927 18717
rect 26513 18717 26525 18720
rect 26559 18748 26571 18751
rect 27617 18751 27675 18757
rect 27617 18748 27629 18751
rect 26559 18720 27629 18748
rect 26559 18717 26571 18720
rect 26513 18711 26571 18717
rect 27617 18717 27629 18720
rect 27663 18717 27675 18751
rect 27617 18711 27675 18717
rect 37829 18751 37887 18757
rect 37829 18717 37841 18751
rect 37875 18748 37887 18751
rect 38102 18748 38108 18760
rect 37875 18720 38108 18748
rect 37875 18717 37887 18720
rect 37829 18711 37887 18717
rect 38102 18708 38108 18720
rect 38160 18708 38166 18760
rect 21726 18640 21732 18692
rect 21784 18680 21790 18692
rect 23201 18683 23259 18689
rect 21784 18652 21829 18680
rect 21784 18640 21790 18652
rect 23201 18649 23213 18683
rect 23247 18649 23259 18683
rect 25516 18680 25544 18708
rect 27065 18683 27123 18689
rect 27065 18680 27077 18683
rect 25516 18652 27077 18680
rect 23201 18643 23259 18649
rect 27065 18649 27077 18652
rect 27111 18649 27123 18683
rect 27065 18643 27123 18649
rect 21085 18615 21143 18621
rect 21085 18581 21097 18615
rect 21131 18612 21143 18615
rect 22646 18612 22652 18624
rect 21131 18584 22652 18612
rect 21131 18581 21143 18584
rect 21085 18575 21143 18581
rect 22646 18572 22652 18584
rect 22704 18572 22710 18624
rect 23216 18612 23244 18643
rect 24673 18615 24731 18621
rect 24673 18612 24685 18615
rect 23216 18584 24685 18612
rect 24673 18581 24685 18584
rect 24719 18581 24731 18615
rect 24673 18575 24731 18581
rect 24762 18572 24768 18624
rect 24820 18612 24826 18624
rect 25317 18615 25375 18621
rect 25317 18612 25329 18615
rect 24820 18584 25329 18612
rect 24820 18572 24826 18584
rect 25317 18581 25329 18584
rect 25363 18581 25375 18615
rect 25317 18575 25375 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 21361 18411 21419 18417
rect 21361 18377 21373 18411
rect 21407 18408 21419 18411
rect 21407 18380 22094 18408
rect 21407 18377 21419 18380
rect 21361 18371 21419 18377
rect 22066 18340 22094 18380
rect 22741 18343 22799 18349
rect 22741 18340 22753 18343
rect 22066 18312 22753 18340
rect 22741 18309 22753 18312
rect 22787 18309 22799 18343
rect 25406 18340 25412 18352
rect 25367 18312 25412 18340
rect 22741 18303 22799 18309
rect 25406 18300 25412 18312
rect 25464 18300 25470 18352
rect 25501 18343 25559 18349
rect 25501 18309 25513 18343
rect 25547 18340 25559 18343
rect 26326 18340 26332 18352
rect 25547 18312 26332 18340
rect 25547 18309 25559 18312
rect 25501 18303 25559 18309
rect 26326 18300 26332 18312
rect 26384 18300 26390 18352
rect 26421 18343 26479 18349
rect 26421 18309 26433 18343
rect 26467 18340 26479 18343
rect 26510 18340 26516 18352
rect 26467 18312 26516 18340
rect 26467 18309 26479 18312
rect 26421 18303 26479 18309
rect 26510 18300 26516 18312
rect 26568 18300 26574 18352
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18272 21327 18275
rect 22094 18272 22100 18284
rect 21315 18244 22100 18272
rect 21315 18241 21327 18244
rect 21269 18235 21327 18241
rect 22094 18232 22100 18244
rect 22152 18232 22158 18284
rect 23750 18272 23756 18284
rect 23711 18244 23756 18272
rect 23750 18232 23756 18244
rect 23808 18232 23814 18284
rect 23937 18275 23995 18281
rect 23937 18241 23949 18275
rect 23983 18272 23995 18275
rect 24762 18272 24768 18284
rect 23983 18244 24768 18272
rect 23983 18241 23995 18244
rect 23937 18235 23995 18241
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 22646 18204 22652 18216
rect 22607 18176 22652 18204
rect 22646 18164 22652 18176
rect 22704 18164 22710 18216
rect 23106 18204 23112 18216
rect 23067 18176 23112 18204
rect 23106 18164 23112 18176
rect 23164 18164 23170 18216
rect 23474 18096 23480 18148
rect 23532 18136 23538 18148
rect 24121 18139 24179 18145
rect 24121 18136 24133 18139
rect 23532 18108 24133 18136
rect 23532 18096 23538 18108
rect 24121 18105 24133 18108
rect 24167 18105 24179 18139
rect 24121 18099 24179 18105
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 27154 18068 27160 18080
rect 22152 18040 22197 18068
rect 27115 18040 27160 18068
rect 22152 18028 22158 18040
rect 27154 18028 27160 18040
rect 27212 18028 27218 18080
rect 38102 18068 38108 18080
rect 38063 18040 38108 18068
rect 38102 18028 38108 18040
rect 38160 18028 38166 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 21726 17864 21732 17876
rect 21687 17836 21732 17864
rect 21726 17824 21732 17836
rect 21784 17824 21790 17876
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22373 17867 22431 17873
rect 22373 17864 22385 17867
rect 22244 17836 22385 17864
rect 22244 17824 22250 17836
rect 22373 17833 22385 17836
rect 22419 17833 22431 17867
rect 22373 17827 22431 17833
rect 26326 17824 26332 17876
rect 26384 17864 26390 17876
rect 27525 17867 27583 17873
rect 27525 17864 27537 17867
rect 26384 17836 27537 17864
rect 26384 17824 26390 17836
rect 27525 17833 27537 17836
rect 27571 17833 27583 17867
rect 27525 17827 27583 17833
rect 29825 17867 29883 17873
rect 29825 17833 29837 17867
rect 29871 17864 29883 17867
rect 33134 17864 33140 17876
rect 29871 17836 33140 17864
rect 29871 17833 29883 17836
rect 29825 17827 29883 17833
rect 33134 17824 33140 17836
rect 33192 17824 33198 17876
rect 24949 17799 25007 17805
rect 24949 17796 24961 17799
rect 23492 17768 24961 17796
rect 23492 17740 23520 17768
rect 24949 17765 24961 17768
rect 24995 17765 25007 17799
rect 26878 17796 26884 17808
rect 26839 17768 26884 17796
rect 24949 17759 25007 17765
rect 26878 17756 26884 17768
rect 26936 17756 26942 17808
rect 20625 17731 20683 17737
rect 20625 17697 20637 17731
rect 20671 17728 20683 17731
rect 22094 17728 22100 17740
rect 20671 17700 22100 17728
rect 20671 17697 20683 17700
rect 20625 17691 20683 17697
rect 22066 17688 22100 17700
rect 22152 17688 22158 17740
rect 23017 17731 23075 17737
rect 23017 17697 23029 17731
rect 23063 17728 23075 17731
rect 23474 17728 23480 17740
rect 23063 17700 23480 17728
rect 23063 17697 23075 17700
rect 23017 17691 23075 17697
rect 23474 17688 23480 17700
rect 23532 17688 23538 17740
rect 24029 17731 24087 17737
rect 24029 17697 24041 17731
rect 24075 17728 24087 17731
rect 24210 17728 24216 17740
rect 24075 17700 24216 17728
rect 24075 17697 24087 17700
rect 24029 17691 24087 17697
rect 24210 17688 24216 17700
rect 24268 17688 24274 17740
rect 25682 17728 25688 17740
rect 25643 17700 25688 17728
rect 25682 17688 25688 17700
rect 25740 17688 25746 17740
rect 26694 17688 26700 17740
rect 26752 17728 26758 17740
rect 26752 17700 29776 17728
rect 26752 17688 26758 17700
rect 21821 17663 21879 17669
rect 21821 17660 21833 17663
rect 21192 17632 21833 17660
rect 21192 17536 21220 17632
rect 21821 17629 21833 17632
rect 21867 17629 21879 17663
rect 22066 17660 22094 17688
rect 22465 17663 22523 17669
rect 22465 17660 22477 17663
rect 22066 17632 22477 17660
rect 21821 17623 21879 17629
rect 22465 17629 22477 17632
rect 22511 17660 22523 17663
rect 22738 17660 22744 17672
rect 22511 17632 22744 17660
rect 22511 17629 22523 17632
rect 22465 17623 22523 17629
rect 22738 17620 22744 17632
rect 22796 17620 22802 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17629 24639 17663
rect 24762 17660 24768 17672
rect 24723 17632 24768 17660
rect 24581 17623 24639 17629
rect 23109 17595 23167 17601
rect 23109 17561 23121 17595
rect 23155 17561 23167 17595
rect 23109 17555 23167 17561
rect 21174 17524 21180 17536
rect 21135 17496 21180 17524
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 22646 17484 22652 17536
rect 22704 17524 22710 17536
rect 23124 17524 23152 17555
rect 23290 17552 23296 17604
rect 23348 17592 23354 17604
rect 24596 17592 24624 17623
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25866 17660 25872 17672
rect 25827 17632 25872 17660
rect 25866 17620 25872 17632
rect 25924 17620 25930 17672
rect 26602 17620 26608 17672
rect 26660 17660 26666 17672
rect 26973 17663 27031 17669
rect 26973 17660 26985 17663
rect 26660 17632 26985 17660
rect 26660 17620 26666 17632
rect 26973 17629 26985 17632
rect 27019 17660 27031 17663
rect 27154 17660 27160 17672
rect 27019 17632 27160 17660
rect 27019 17629 27031 17632
rect 26973 17623 27031 17629
rect 27154 17620 27160 17632
rect 27212 17620 27218 17672
rect 29748 17669 29776 17700
rect 27617 17663 27675 17669
rect 27617 17629 27629 17663
rect 27663 17660 27675 17663
rect 29733 17663 29791 17669
rect 27663 17632 28212 17660
rect 27663 17629 27675 17632
rect 27617 17623 27675 17629
rect 23348 17564 24624 17592
rect 23348 17552 23354 17564
rect 22704 17496 23152 17524
rect 22704 17484 22710 17496
rect 26234 17484 26240 17536
rect 26292 17524 26298 17536
rect 28184 17533 28212 17632
rect 29733 17629 29745 17663
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 26329 17527 26387 17533
rect 26329 17524 26341 17527
rect 26292 17496 26341 17524
rect 26292 17484 26298 17496
rect 26329 17493 26341 17496
rect 26375 17493 26387 17527
rect 26329 17487 26387 17493
rect 28169 17527 28227 17533
rect 28169 17493 28181 17527
rect 28215 17524 28227 17527
rect 31202 17524 31208 17536
rect 28215 17496 31208 17524
rect 28215 17493 28227 17496
rect 28169 17487 28227 17493
rect 31202 17484 31208 17496
rect 31260 17484 31266 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 23106 17280 23112 17332
rect 23164 17320 23170 17332
rect 24305 17323 24363 17329
rect 23164 17292 23888 17320
rect 23164 17280 23170 17292
rect 22465 17255 22523 17261
rect 22465 17221 22477 17255
rect 22511 17252 22523 17255
rect 23201 17255 23259 17261
rect 23201 17252 23213 17255
rect 22511 17224 23213 17252
rect 22511 17221 22523 17224
rect 22465 17215 22523 17221
rect 23201 17221 23213 17224
rect 23247 17221 23259 17255
rect 23860 17252 23888 17292
rect 24305 17289 24317 17323
rect 24351 17320 24363 17323
rect 24762 17320 24768 17332
rect 24351 17292 24768 17320
rect 24351 17289 24363 17292
rect 24305 17283 24363 17289
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 25866 17280 25872 17332
rect 25924 17320 25930 17332
rect 27893 17323 27951 17329
rect 27893 17320 27905 17323
rect 25924 17292 27905 17320
rect 25924 17280 25930 17292
rect 27893 17289 27905 17292
rect 27939 17289 27951 17323
rect 27893 17283 27951 17289
rect 25225 17255 25283 17261
rect 25225 17252 25237 17255
rect 23860 17224 25237 17252
rect 23201 17215 23259 17221
rect 25225 17221 25237 17224
rect 25271 17221 25283 17255
rect 25225 17215 25283 17221
rect 25317 17255 25375 17261
rect 25317 17221 25329 17255
rect 25363 17252 25375 17255
rect 26237 17255 26295 17261
rect 25363 17224 26188 17252
rect 25363 17221 25375 17224
rect 25317 17215 25375 17221
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 6822 17184 6828 17196
rect 1903 17156 6828 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17184 20959 17187
rect 22373 17187 22431 17193
rect 22373 17184 22385 17187
rect 20947 17156 22385 17184
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 22373 17153 22385 17156
rect 22419 17184 22431 17187
rect 22738 17184 22744 17196
rect 22419 17156 22744 17184
rect 22419 17153 22431 17156
rect 22373 17147 22431 17153
rect 22738 17144 22744 17156
rect 22796 17144 22802 17196
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17184 24271 17187
rect 24394 17184 24400 17196
rect 24259 17156 24400 17184
rect 24259 17153 24271 17156
rect 24213 17147 24271 17153
rect 24394 17144 24400 17156
rect 24452 17144 24458 17196
rect 26160 17184 26188 17224
rect 26237 17221 26249 17255
rect 26283 17252 26295 17255
rect 26510 17252 26516 17264
rect 26283 17224 26516 17252
rect 26283 17221 26295 17224
rect 26237 17215 26295 17221
rect 26510 17212 26516 17224
rect 26568 17212 26574 17264
rect 27430 17184 27436 17196
rect 26160 17156 27436 17184
rect 27430 17144 27436 17156
rect 27488 17144 27494 17196
rect 27522 17144 27528 17196
rect 27580 17184 27586 17196
rect 27801 17187 27859 17193
rect 27801 17184 27813 17187
rect 27580 17156 27813 17184
rect 27580 17144 27586 17156
rect 27801 17153 27813 17156
rect 27847 17153 27859 17187
rect 27801 17147 27859 17153
rect 37645 17187 37703 17193
rect 37645 17153 37657 17187
rect 37691 17184 37703 17187
rect 38286 17184 38292 17196
rect 37691 17156 38292 17184
rect 37691 17153 37703 17156
rect 37645 17147 37703 17153
rect 38286 17144 38292 17156
rect 38344 17144 38350 17196
rect 23109 17119 23167 17125
rect 23109 17085 23121 17119
rect 23155 17116 23167 17119
rect 23382 17116 23388 17128
rect 23155 17088 23388 17116
rect 23155 17085 23167 17088
rect 23109 17079 23167 17085
rect 23382 17076 23388 17088
rect 23440 17076 23446 17128
rect 26326 17076 26332 17128
rect 26384 17116 26390 17128
rect 27157 17119 27215 17125
rect 27157 17116 27169 17119
rect 26384 17088 27169 17116
rect 26384 17076 26390 17088
rect 27157 17085 27169 17088
rect 27203 17085 27215 17119
rect 27157 17079 27215 17085
rect 1670 17048 1676 17060
rect 1631 17020 1676 17048
rect 1670 17008 1676 17020
rect 1728 17008 1734 17060
rect 23198 17008 23204 17060
rect 23256 17048 23262 17060
rect 23661 17051 23719 17057
rect 23661 17048 23673 17051
rect 23256 17020 23673 17048
rect 23256 17008 23262 17020
rect 23661 17017 23673 17020
rect 23707 17017 23719 17051
rect 23661 17011 23719 17017
rect 21174 16940 21180 16992
rect 21232 16980 21238 16992
rect 21361 16983 21419 16989
rect 21361 16980 21373 16983
rect 21232 16952 21373 16980
rect 21232 16940 21238 16952
rect 21361 16949 21373 16952
rect 21407 16949 21419 16983
rect 23676 16980 23704 17011
rect 24394 17008 24400 17060
rect 24452 17048 24458 17060
rect 28445 17051 28503 17057
rect 28445 17048 28457 17051
rect 24452 17020 28457 17048
rect 24452 17008 24458 17020
rect 28445 17017 28457 17020
rect 28491 17017 28503 17051
rect 28445 17011 28503 17017
rect 25038 16980 25044 16992
rect 23676 16952 25044 16980
rect 21361 16943 21419 16949
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 37918 16940 37924 16992
rect 37976 16980 37982 16992
rect 38105 16983 38163 16989
rect 38105 16980 38117 16983
rect 37976 16952 38117 16980
rect 37976 16940 37982 16952
rect 38105 16949 38117 16952
rect 38151 16949 38163 16983
rect 38105 16943 38163 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 2409 16779 2467 16785
rect 2409 16776 2421 16779
rect 2280 16748 2421 16776
rect 2280 16736 2286 16748
rect 2409 16745 2421 16748
rect 2455 16745 2467 16779
rect 23290 16776 23296 16788
rect 2409 16739 2467 16745
rect 22066 16748 23296 16776
rect 10778 16640 10784 16652
rect 10244 16612 10784 16640
rect 1949 16575 2007 16581
rect 1949 16541 1961 16575
rect 1995 16572 2007 16575
rect 2222 16572 2228 16584
rect 1995 16544 2228 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 10134 16572 10140 16584
rect 10047 16544 10140 16572
rect 10134 16532 10140 16544
rect 10192 16572 10198 16584
rect 10244 16572 10272 16612
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 20070 16640 20076 16652
rect 20031 16612 20076 16640
rect 20070 16600 20076 16612
rect 20128 16600 20134 16652
rect 22066 16640 22094 16748
rect 23290 16736 23296 16748
rect 23348 16736 23354 16788
rect 25314 16736 25320 16788
rect 25372 16776 25378 16788
rect 28169 16779 28227 16785
rect 28169 16776 28181 16779
rect 25372 16748 28181 16776
rect 25372 16736 25378 16748
rect 28169 16745 28181 16748
rect 28215 16776 28227 16779
rect 34790 16776 34796 16788
rect 28215 16748 34796 16776
rect 28215 16745 28227 16748
rect 28169 16739 28227 16745
rect 34790 16736 34796 16748
rect 34848 16736 34854 16788
rect 23106 16708 23112 16720
rect 23067 16680 23112 16708
rect 23106 16668 23112 16680
rect 23164 16668 23170 16720
rect 24780 16680 26924 16708
rect 21100 16612 21404 16640
rect 21100 16572 21128 16612
rect 10192 16544 10272 16572
rect 16546 16544 21128 16572
rect 10192 16532 10198 16544
rect 10229 16507 10287 16513
rect 10229 16473 10241 16507
rect 10275 16504 10287 16507
rect 16546 16504 16574 16544
rect 21174 16532 21180 16584
rect 21232 16572 21238 16584
rect 21376 16572 21404 16612
rect 21928 16612 22094 16640
rect 22388 16612 23244 16640
rect 21928 16572 21956 16612
rect 21232 16544 21277 16572
rect 21376 16544 21956 16572
rect 22005 16575 22063 16581
rect 21232 16532 21238 16544
rect 22005 16541 22017 16575
rect 22051 16572 22063 16575
rect 22388 16572 22416 16612
rect 22051 16544 22416 16572
rect 23216 16572 23244 16612
rect 23566 16572 23572 16584
rect 23216 16544 23572 16572
rect 22051 16541 22063 16544
rect 22005 16535 22063 16541
rect 23566 16532 23572 16544
rect 23624 16572 23630 16584
rect 23937 16575 23995 16581
rect 23937 16572 23949 16575
rect 23624 16544 23949 16572
rect 23624 16532 23630 16544
rect 23937 16541 23949 16544
rect 23983 16541 23995 16575
rect 23937 16535 23995 16541
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16572 24639 16575
rect 24780 16572 24808 16680
rect 25038 16600 25044 16652
rect 25096 16640 25102 16652
rect 25317 16643 25375 16649
rect 25317 16640 25329 16643
rect 25096 16612 25329 16640
rect 25096 16600 25102 16612
rect 25317 16609 25329 16612
rect 25363 16609 25375 16643
rect 25317 16603 25375 16609
rect 26145 16643 26203 16649
rect 26145 16609 26157 16643
rect 26191 16640 26203 16643
rect 26510 16640 26516 16652
rect 26191 16612 26516 16640
rect 26191 16609 26203 16612
rect 26145 16603 26203 16609
rect 26510 16600 26516 16612
rect 26568 16600 26574 16652
rect 24627 16544 24808 16572
rect 26896 16572 26924 16680
rect 26970 16572 26976 16584
rect 26896 16544 26976 16572
rect 24627 16541 24639 16544
rect 24581 16535 24639 16541
rect 20254 16504 20260 16516
rect 10275 16476 16574 16504
rect 20215 16476 20260 16504
rect 10275 16473 10287 16476
rect 10229 16467 10287 16473
rect 20254 16464 20260 16476
rect 20312 16464 20318 16516
rect 21269 16507 21327 16513
rect 21269 16473 21281 16507
rect 21315 16504 21327 16507
rect 22554 16504 22560 16516
rect 21315 16476 22094 16504
rect 22515 16476 22560 16504
rect 21315 16473 21327 16476
rect 21269 16467 21327 16473
rect 1762 16436 1768 16448
rect 1723 16408 1768 16436
rect 1762 16396 1768 16408
rect 1820 16396 1826 16448
rect 21818 16436 21824 16448
rect 21779 16408 21824 16436
rect 21818 16396 21824 16408
rect 21876 16396 21882 16448
rect 22066 16436 22094 16476
rect 22554 16464 22560 16476
rect 22612 16464 22618 16516
rect 22649 16507 22707 16513
rect 22649 16473 22661 16507
rect 22695 16473 22707 16507
rect 22649 16467 22707 16473
rect 22664 16436 22692 16467
rect 23474 16464 23480 16516
rect 23532 16504 23538 16516
rect 23661 16507 23719 16513
rect 23661 16504 23673 16507
rect 23532 16476 23673 16504
rect 23532 16464 23538 16476
rect 23661 16473 23673 16476
rect 23707 16473 23719 16507
rect 23952 16504 23980 16535
rect 26970 16532 26976 16544
rect 27028 16532 27034 16584
rect 27154 16532 27160 16584
rect 27212 16572 27218 16584
rect 27522 16572 27528 16584
rect 27212 16544 27528 16572
rect 27212 16532 27218 16544
rect 27522 16532 27528 16544
rect 27580 16572 27586 16584
rect 27617 16575 27675 16581
rect 27617 16572 27629 16575
rect 27580 16544 27629 16572
rect 27580 16532 27586 16544
rect 27617 16541 27629 16544
rect 27663 16541 27675 16575
rect 27617 16535 27675 16541
rect 25314 16504 25320 16516
rect 23952 16476 25320 16504
rect 23661 16467 23719 16473
rect 25314 16464 25320 16476
rect 25372 16464 25378 16516
rect 25409 16507 25467 16513
rect 25409 16473 25421 16507
rect 25455 16504 25467 16507
rect 27338 16504 27344 16516
rect 25455 16476 27344 16504
rect 25455 16473 25467 16476
rect 25409 16467 25467 16473
rect 27338 16464 27344 16476
rect 27396 16464 27402 16516
rect 22066 16408 22692 16436
rect 24673 16439 24731 16445
rect 24673 16405 24685 16439
rect 24719 16436 24731 16439
rect 24762 16436 24768 16448
rect 24719 16408 24768 16436
rect 24719 16405 24731 16408
rect 24673 16399 24731 16405
rect 24762 16396 24768 16408
rect 24820 16396 24826 16448
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 26881 16439 26939 16445
rect 26881 16436 26893 16439
rect 24912 16408 26893 16436
rect 24912 16396 24918 16408
rect 26881 16405 26893 16408
rect 26927 16405 26939 16439
rect 27522 16436 27528 16448
rect 27483 16408 27528 16436
rect 26881 16399 26939 16405
rect 27522 16396 27528 16408
rect 27580 16396 27586 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 21361 16235 21419 16241
rect 21361 16201 21373 16235
rect 21407 16232 21419 16235
rect 22646 16232 22652 16244
rect 21407 16204 22652 16232
rect 21407 16201 21419 16204
rect 21361 16195 21419 16201
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 37826 16232 37832 16244
rect 22848 16204 37832 16232
rect 20254 16124 20260 16176
rect 20312 16164 20318 16176
rect 20533 16167 20591 16173
rect 20533 16164 20545 16167
rect 20312 16136 20545 16164
rect 20312 16124 20318 16136
rect 20533 16133 20545 16136
rect 20579 16164 20591 16167
rect 22848 16164 22876 16204
rect 37826 16192 37832 16204
rect 37884 16192 37890 16244
rect 23474 16164 23480 16176
rect 20579 16136 22876 16164
rect 22940 16136 23480 16164
rect 20579 16133 20591 16136
rect 20533 16127 20591 16133
rect 21450 16096 21456 16108
rect 21411 16068 21456 16096
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 22940 16105 22968 16136
rect 23474 16124 23480 16136
rect 23532 16124 23538 16176
rect 23569 16167 23627 16173
rect 23569 16133 23581 16167
rect 23615 16164 23627 16167
rect 23934 16164 23940 16176
rect 23615 16136 23940 16164
rect 23615 16133 23627 16136
rect 23569 16127 23627 16133
rect 23934 16124 23940 16136
rect 23992 16124 23998 16176
rect 26053 16167 26111 16173
rect 26053 16133 26065 16167
rect 26099 16164 26111 16167
rect 27062 16164 27068 16176
rect 26099 16136 27068 16164
rect 26099 16133 26111 16136
rect 26053 16127 26111 16133
rect 27062 16124 27068 16136
rect 27120 16124 27126 16176
rect 22925 16099 22983 16105
rect 22925 16065 22937 16099
rect 22971 16065 22983 16099
rect 24578 16096 24584 16108
rect 24539 16068 24584 16096
rect 22925 16059 22983 16065
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 24762 16096 24768 16108
rect 24723 16068 24768 16096
rect 24762 16056 24768 16068
rect 24820 16056 24826 16108
rect 26605 16099 26663 16105
rect 26605 16065 26617 16099
rect 26651 16096 26663 16099
rect 26694 16096 26700 16108
rect 26651 16068 26700 16096
rect 26651 16065 26663 16068
rect 26605 16059 26663 16065
rect 26694 16056 26700 16068
rect 26752 16056 26758 16108
rect 27154 16096 27160 16108
rect 27115 16068 27160 16096
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 22741 16031 22799 16037
rect 22741 15997 22753 16031
rect 22787 15997 22799 16031
rect 22741 15991 22799 15997
rect 23477 16031 23535 16037
rect 23477 15997 23489 16031
rect 23523 16028 23535 16031
rect 23750 16028 23756 16040
rect 23523 16000 23756 16028
rect 23523 15997 23535 16000
rect 23477 15991 23535 15997
rect 22756 15960 22784 15991
rect 23750 15988 23756 16000
rect 23808 15988 23814 16040
rect 25961 16031 26019 16037
rect 25961 15997 25973 16031
rect 26007 16028 26019 16031
rect 26234 16028 26240 16040
rect 26007 16000 26240 16028
rect 26007 15997 26019 16000
rect 25961 15991 26019 15997
rect 23842 15960 23848 15972
rect 22756 15932 23848 15960
rect 23842 15920 23848 15932
rect 23900 15920 23906 15972
rect 24026 15960 24032 15972
rect 23987 15932 24032 15960
rect 24026 15920 24032 15932
rect 24084 15920 24090 15972
rect 25976 15960 26004 15991
rect 26234 15988 26240 16000
rect 26292 15988 26298 16040
rect 24964 15932 26004 15960
rect 22557 15895 22615 15901
rect 22557 15861 22569 15895
rect 22603 15892 22615 15895
rect 24964 15892 24992 15932
rect 22603 15864 24992 15892
rect 25225 15895 25283 15901
rect 22603 15861 22615 15864
rect 22557 15855 22615 15861
rect 25225 15861 25237 15895
rect 25271 15892 25283 15895
rect 25682 15892 25688 15904
rect 25271 15864 25688 15892
rect 25271 15861 25283 15864
rect 25225 15855 25283 15861
rect 25682 15852 25688 15864
rect 25740 15852 25746 15904
rect 27246 15892 27252 15904
rect 27207 15864 27252 15892
rect 27246 15852 27252 15864
rect 27304 15852 27310 15904
rect 27890 15892 27896 15904
rect 27851 15864 27896 15892
rect 27890 15852 27896 15864
rect 27948 15852 27954 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6880 15660 6929 15688
rect 6880 15648 6886 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 22189 15691 22247 15697
rect 22189 15657 22201 15691
rect 22235 15688 22247 15691
rect 22554 15688 22560 15700
rect 22235 15660 22560 15688
rect 22235 15657 22247 15660
rect 22189 15651 22247 15657
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 22940 15660 26372 15688
rect 21450 15580 21456 15632
rect 21508 15620 21514 15632
rect 21545 15623 21603 15629
rect 21545 15620 21557 15623
rect 21508 15592 21557 15620
rect 21508 15580 21514 15592
rect 21545 15589 21557 15592
rect 21591 15620 21603 15623
rect 22940 15620 22968 15660
rect 21591 15592 22968 15620
rect 21591 15589 21603 15592
rect 21545 15583 21603 15589
rect 23014 15580 23020 15632
rect 23072 15620 23078 15632
rect 25225 15623 25283 15629
rect 23072 15592 24624 15620
rect 23072 15580 23078 15592
rect 24596 15564 24624 15592
rect 25225 15589 25237 15623
rect 25271 15620 25283 15623
rect 26234 15620 26240 15632
rect 25271 15592 26240 15620
rect 25271 15589 25283 15592
rect 25225 15583 25283 15589
rect 26234 15580 26240 15592
rect 26292 15580 26298 15632
rect 26344 15620 26372 15660
rect 27430 15648 27436 15700
rect 27488 15688 27494 15700
rect 27525 15691 27583 15697
rect 27525 15688 27537 15691
rect 27488 15660 27537 15688
rect 27488 15648 27494 15660
rect 27525 15657 27537 15660
rect 27571 15657 27583 15691
rect 27525 15651 27583 15657
rect 29362 15620 29368 15632
rect 26344 15592 29368 15620
rect 29362 15580 29368 15592
rect 29420 15580 29426 15632
rect 23106 15552 23112 15564
rect 23067 15524 23112 15552
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 24578 15552 24584 15564
rect 24491 15524 24584 15552
rect 24578 15512 24584 15524
rect 24636 15512 24642 15564
rect 24765 15555 24823 15561
rect 24765 15521 24777 15555
rect 24811 15552 24823 15555
rect 24854 15552 24860 15564
rect 24811 15524 24860 15552
rect 24811 15521 24823 15524
rect 24765 15515 24823 15521
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 25682 15552 25688 15564
rect 25643 15524 25688 15552
rect 25682 15512 25688 15524
rect 25740 15512 25746 15564
rect 26145 15555 26203 15561
rect 26145 15521 26157 15555
rect 26191 15552 26203 15555
rect 27522 15552 27528 15564
rect 26191 15524 27528 15552
rect 26191 15521 26203 15524
rect 26145 15515 26203 15521
rect 27522 15512 27528 15524
rect 27580 15512 27586 15564
rect 27890 15552 27896 15564
rect 27632 15524 27896 15552
rect 1857 15487 1915 15493
rect 1857 15453 1869 15487
rect 1903 15484 1915 15487
rect 7101 15487 7159 15493
rect 1903 15456 6914 15484
rect 1903 15453 1915 15456
rect 1857 15447 1915 15453
rect 1670 15348 1676 15360
rect 1631 15320 1676 15348
rect 1670 15308 1676 15320
rect 1728 15308 1734 15360
rect 6886 15348 6914 15456
rect 7101 15453 7113 15487
rect 7147 15453 7159 15487
rect 22186 15484 22192 15496
rect 22099 15456 22192 15484
rect 7101 15447 7159 15453
rect 7116 15416 7144 15447
rect 22186 15444 22192 15456
rect 22244 15484 22250 15496
rect 26326 15484 26332 15496
rect 22244 15456 22692 15484
rect 26287 15456 26332 15484
rect 22244 15444 22250 15456
rect 7653 15419 7711 15425
rect 7653 15416 7665 15419
rect 7116 15388 7665 15416
rect 7653 15385 7665 15388
rect 7699 15416 7711 15419
rect 19150 15416 19156 15428
rect 7699 15388 19156 15416
rect 7699 15385 7711 15388
rect 7653 15379 7711 15385
rect 19150 15376 19156 15388
rect 19208 15376 19214 15428
rect 12158 15348 12164 15360
rect 6886 15320 12164 15348
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 22664 15348 22692 15456
rect 26326 15444 26332 15456
rect 26384 15444 26390 15496
rect 27632 15493 27660 15524
rect 27890 15512 27896 15524
rect 27948 15552 27954 15564
rect 30466 15552 30472 15564
rect 27948 15524 30472 15552
rect 27948 15512 27954 15524
rect 30466 15512 30472 15524
rect 30524 15512 30530 15564
rect 26789 15487 26847 15493
rect 26789 15453 26801 15487
rect 26835 15453 26847 15487
rect 26789 15447 26847 15453
rect 27617 15487 27675 15493
rect 27617 15453 27629 15487
rect 27663 15453 27675 15487
rect 27617 15447 27675 15453
rect 28261 15487 28319 15493
rect 28261 15453 28273 15487
rect 28307 15453 28319 15487
rect 38010 15484 38016 15496
rect 37971 15456 38016 15484
rect 28261 15447 28319 15453
rect 22830 15416 22836 15428
rect 22791 15388 22836 15416
rect 22830 15376 22836 15388
rect 22888 15376 22894 15428
rect 22922 15376 22928 15428
rect 22980 15416 22986 15428
rect 22980 15388 23025 15416
rect 22980 15376 22986 15388
rect 25866 15376 25872 15428
rect 25924 15416 25930 15428
rect 26804 15416 26832 15447
rect 25924 15388 26832 15416
rect 28276 15416 28304 15447
rect 38010 15444 38016 15456
rect 38068 15444 38074 15496
rect 28813 15419 28871 15425
rect 28813 15416 28825 15419
rect 28276 15388 28825 15416
rect 25924 15376 25930 15388
rect 28813 15385 28825 15388
rect 28859 15416 28871 15419
rect 37274 15416 37280 15428
rect 28859 15388 37280 15416
rect 28859 15385 28871 15388
rect 28813 15379 28871 15385
rect 37274 15376 37280 15388
rect 37332 15376 37338 15428
rect 23198 15348 23204 15360
rect 22664 15320 23204 15348
rect 23198 15308 23204 15320
rect 23256 15348 23262 15360
rect 23937 15351 23995 15357
rect 23937 15348 23949 15351
rect 23256 15320 23949 15348
rect 23256 15308 23262 15320
rect 23937 15317 23949 15320
rect 23983 15317 23995 15351
rect 23937 15311 23995 15317
rect 26326 15308 26332 15360
rect 26384 15348 26390 15360
rect 26881 15351 26939 15357
rect 26881 15348 26893 15351
rect 26384 15320 26893 15348
rect 26384 15308 26390 15320
rect 26881 15317 26893 15320
rect 26927 15317 26939 15351
rect 28166 15348 28172 15360
rect 28127 15320 28172 15348
rect 26881 15311 26939 15317
rect 28166 15308 28172 15320
rect 28224 15308 28230 15360
rect 38194 15348 38200 15360
rect 38155 15320 38200 15348
rect 38194 15308 38200 15320
rect 38252 15308 38258 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 12158 15144 12164 15156
rect 12119 15116 12164 15144
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 22741 15147 22799 15153
rect 22741 15113 22753 15147
rect 22787 15144 22799 15147
rect 22922 15144 22928 15156
rect 22787 15116 22928 15144
rect 22787 15113 22799 15116
rect 22741 15107 22799 15113
rect 22922 15104 22928 15116
rect 22980 15104 22986 15156
rect 23566 15144 23572 15156
rect 23308 15116 23572 15144
rect 22189 15079 22247 15085
rect 22189 15045 22201 15079
rect 22235 15076 22247 15079
rect 23308 15076 23336 15116
rect 23566 15104 23572 15116
rect 23624 15104 23630 15156
rect 23842 15104 23848 15156
rect 23900 15144 23906 15156
rect 25777 15147 25835 15153
rect 25777 15144 25789 15147
rect 23900 15116 25789 15144
rect 23900 15104 23906 15116
rect 25777 15113 25789 15116
rect 25823 15113 25835 15147
rect 25777 15107 25835 15113
rect 27338 15104 27344 15156
rect 27396 15144 27402 15156
rect 28353 15147 28411 15153
rect 28353 15144 28365 15147
rect 27396 15116 28365 15144
rect 27396 15104 27402 15116
rect 28353 15113 28365 15116
rect 28399 15113 28411 15147
rect 28353 15107 28411 15113
rect 23474 15076 23480 15088
rect 22235 15048 23336 15076
rect 23435 15048 23480 15076
rect 22235 15045 22247 15048
rect 22189 15039 22247 15045
rect 23474 15036 23480 15048
rect 23532 15036 23538 15088
rect 24026 15076 24032 15088
rect 23987 15048 24032 15076
rect 24026 15036 24032 15048
rect 24084 15036 24090 15088
rect 24578 15076 24584 15088
rect 24539 15048 24584 15076
rect 24578 15036 24584 15048
rect 24636 15036 24642 15088
rect 24673 15079 24731 15085
rect 24673 15045 24685 15079
rect 24719 15076 24731 15079
rect 26421 15079 26479 15085
rect 26421 15076 26433 15079
rect 24719 15048 26433 15076
rect 24719 15045 24731 15048
rect 24673 15039 24731 15045
rect 26421 15045 26433 15048
rect 26467 15045 26479 15079
rect 26421 15039 26479 15045
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 15008 12403 15011
rect 21453 15011 21511 15017
rect 12391 14980 12940 15008
rect 12391 14977 12403 14980
rect 12345 14971 12403 14977
rect 12912 14881 12940 14980
rect 21453 14977 21465 15011
rect 21499 15008 21511 15011
rect 22554 15008 22560 15020
rect 21499 14980 22560 15008
rect 21499 14977 21511 14980
rect 21453 14971 21511 14977
rect 22554 14968 22560 14980
rect 22612 15008 22618 15020
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 22612 14980 22661 15008
rect 22612 14968 22618 14980
rect 22649 14977 22661 14980
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 25590 14968 25596 15020
rect 25648 15008 25654 15020
rect 25866 15008 25872 15020
rect 25648 14980 25872 15008
rect 25648 14968 25654 14980
rect 25866 14968 25872 14980
rect 25924 14968 25930 15020
rect 26234 14968 26240 15020
rect 26292 15008 26298 15020
rect 26513 15011 26571 15017
rect 26513 15008 26525 15011
rect 26292 14980 26525 15008
rect 26292 14968 26298 14980
rect 26513 14977 26525 14980
rect 26559 14977 26571 15011
rect 26513 14971 26571 14977
rect 27246 14968 27252 15020
rect 27304 15008 27310 15020
rect 27341 15011 27399 15017
rect 27341 15008 27353 15011
rect 27304 14980 27353 15008
rect 27304 14968 27310 14980
rect 27341 14977 27353 14980
rect 27387 14977 27399 15011
rect 27341 14971 27399 14977
rect 28445 15011 28503 15017
rect 28445 14977 28457 15011
rect 28491 15008 28503 15011
rect 28534 15008 28540 15020
rect 28491 14980 28540 15008
rect 28491 14977 28503 14980
rect 28445 14971 28503 14977
rect 28534 14968 28540 14980
rect 28592 14968 28598 15020
rect 23382 14940 23388 14952
rect 23343 14912 23388 14940
rect 23382 14900 23388 14912
rect 23440 14900 23446 14952
rect 25225 14943 25283 14949
rect 25225 14909 25237 14943
rect 25271 14940 25283 14943
rect 26418 14940 26424 14952
rect 25271 14912 26424 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 27157 14943 27215 14949
rect 27157 14909 27169 14943
rect 27203 14940 27215 14943
rect 27614 14940 27620 14952
rect 27203 14912 27620 14940
rect 27203 14909 27215 14912
rect 27157 14903 27215 14909
rect 27614 14900 27620 14912
rect 27672 14940 27678 14952
rect 28166 14940 28172 14952
rect 27672 14912 28172 14940
rect 27672 14900 27678 14912
rect 28166 14900 28172 14912
rect 28224 14900 28230 14952
rect 12897 14875 12955 14881
rect 12897 14841 12909 14875
rect 12943 14872 12955 14875
rect 22186 14872 22192 14884
rect 12943 14844 22192 14872
rect 12943 14841 12955 14844
rect 12897 14835 12955 14841
rect 22186 14832 22192 14844
rect 22244 14832 22250 14884
rect 27706 14804 27712 14816
rect 27667 14776 27712 14804
rect 27706 14764 27712 14776
rect 27764 14764 27770 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 1949 14603 2007 14609
rect 1949 14600 1961 14603
rect 1912 14572 1961 14600
rect 1912 14560 1918 14572
rect 1949 14569 1961 14572
rect 1995 14569 2007 14603
rect 35710 14600 35716 14612
rect 35671 14572 35716 14600
rect 1949 14563 2007 14569
rect 35710 14560 35716 14572
rect 35768 14560 35774 14612
rect 27706 14532 27712 14544
rect 24780 14504 27712 14532
rect 22094 14424 22100 14476
rect 22152 14464 22158 14476
rect 22741 14467 22799 14473
rect 22152 14436 22197 14464
rect 22152 14424 22158 14436
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 23106 14464 23112 14476
rect 22787 14436 23112 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 23106 14424 23112 14436
rect 23164 14424 23170 14476
rect 12066 14396 12072 14408
rect 12027 14368 12072 14396
rect 12066 14356 12072 14368
rect 12124 14396 12130 14408
rect 12713 14399 12771 14405
rect 12713 14396 12725 14399
rect 12124 14368 12725 14396
rect 12124 14356 12130 14368
rect 12713 14365 12725 14368
rect 12759 14365 12771 14399
rect 23382 14396 23388 14408
rect 23343 14368 23388 14396
rect 12713 14359 12771 14365
rect 23382 14356 23388 14368
rect 23440 14356 23446 14408
rect 23566 14396 23572 14408
rect 23527 14368 23572 14396
rect 23566 14356 23572 14368
rect 23624 14356 23630 14408
rect 24780 14405 24808 14504
rect 27706 14492 27712 14504
rect 27764 14532 27770 14544
rect 27764 14504 28028 14532
rect 27764 14492 27770 14504
rect 25225 14467 25283 14473
rect 25225 14433 25237 14467
rect 25271 14464 25283 14467
rect 26326 14464 26332 14476
rect 25271 14436 26332 14464
rect 25271 14433 25283 14436
rect 25225 14427 25283 14433
rect 26326 14424 26332 14436
rect 26384 14424 26390 14476
rect 26418 14424 26424 14476
rect 26476 14464 26482 14476
rect 26789 14467 26847 14473
rect 26476 14436 26521 14464
rect 26476 14424 26482 14436
rect 26789 14433 26801 14467
rect 26835 14464 26847 14467
rect 27614 14464 27620 14476
rect 26835 14436 27620 14464
rect 26835 14433 26847 14436
rect 26789 14427 26847 14433
rect 27614 14424 27620 14436
rect 27672 14424 27678 14476
rect 28000 14473 28028 14504
rect 27985 14467 28043 14473
rect 27985 14433 27997 14467
rect 28031 14433 28043 14467
rect 27985 14427 28043 14433
rect 24029 14399 24087 14405
rect 24029 14365 24041 14399
rect 24075 14396 24087 14399
rect 24765 14399 24823 14405
rect 24765 14396 24777 14399
rect 24075 14368 24777 14396
rect 24075 14365 24087 14368
rect 24029 14359 24087 14365
rect 24765 14365 24777 14368
rect 24811 14365 24823 14399
rect 24765 14359 24823 14365
rect 25130 14356 25136 14408
rect 25188 14396 25194 14408
rect 25409 14399 25467 14405
rect 25409 14396 25421 14399
rect 25188 14368 25421 14396
rect 25188 14356 25194 14368
rect 25409 14365 25421 14368
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 35342 14356 35348 14408
rect 35400 14396 35406 14408
rect 35529 14399 35587 14405
rect 35529 14396 35541 14399
rect 35400 14368 35541 14396
rect 35400 14356 35406 14368
rect 35529 14365 35541 14368
rect 35575 14365 35587 14399
rect 35529 14359 35587 14365
rect 1857 14331 1915 14337
rect 1857 14297 1869 14331
rect 1903 14328 1915 14331
rect 1946 14328 1952 14340
rect 1903 14300 1952 14328
rect 1903 14297 1915 14300
rect 1857 14291 1915 14297
rect 1946 14288 1952 14300
rect 2004 14328 2010 14340
rect 2501 14331 2559 14337
rect 2501 14328 2513 14331
rect 2004 14300 2513 14328
rect 2004 14288 2010 14300
rect 2501 14297 2513 14300
rect 2547 14297 2559 14331
rect 2501 14291 2559 14297
rect 12161 14331 12219 14337
rect 12161 14297 12173 14331
rect 12207 14328 12219 14331
rect 12207 14300 16574 14328
rect 12207 14297 12219 14300
rect 12161 14291 12219 14297
rect 16546 14260 16574 14300
rect 22186 14288 22192 14340
rect 22244 14328 22250 14340
rect 26694 14328 26700 14340
rect 22244 14300 22289 14328
rect 26655 14300 26700 14328
rect 22244 14288 22250 14300
rect 26694 14288 26700 14300
rect 26752 14288 26758 14340
rect 26786 14288 26792 14340
rect 26844 14328 26850 14340
rect 27341 14331 27399 14337
rect 27341 14328 27353 14331
rect 26844 14300 27353 14328
rect 26844 14288 26850 14300
rect 27341 14297 27353 14300
rect 27387 14297 27399 14331
rect 27890 14328 27896 14340
rect 27851 14300 27896 14328
rect 27341 14291 27399 14297
rect 27890 14288 27896 14300
rect 27948 14288 27954 14340
rect 22646 14260 22652 14272
rect 16546 14232 22652 14260
rect 22646 14220 22652 14232
rect 22704 14260 22710 14272
rect 22830 14260 22836 14272
rect 22704 14232 22836 14260
rect 22704 14220 22710 14232
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 23658 14220 23664 14272
rect 23716 14260 23722 14272
rect 26970 14260 26976 14272
rect 23716 14232 26976 14260
rect 23716 14220 23722 14232
rect 26970 14220 26976 14232
rect 27028 14220 27034 14272
rect 37734 14220 37740 14272
rect 37792 14260 37798 14272
rect 38105 14263 38163 14269
rect 38105 14260 38117 14263
rect 37792 14232 38117 14260
rect 37792 14220 37798 14232
rect 38105 14229 38117 14232
rect 38151 14229 38163 14263
rect 38105 14223 38163 14229
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 22186 14056 22192 14068
rect 22147 14028 22192 14056
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 23293 14059 23351 14065
rect 23293 14025 23305 14059
rect 23339 14056 23351 14059
rect 23566 14056 23572 14068
rect 23339 14028 23572 14056
rect 23339 14025 23351 14028
rect 23293 14019 23351 14025
rect 23566 14016 23572 14028
rect 23624 14016 23630 14068
rect 23934 14056 23940 14068
rect 23895 14028 23940 14056
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 26326 14056 26332 14068
rect 25056 14028 26332 14056
rect 25056 13997 25084 14028
rect 26326 14016 26332 14028
rect 26384 14016 26390 14068
rect 27062 14016 27068 14068
rect 27120 14056 27126 14068
rect 27249 14059 27307 14065
rect 27249 14056 27261 14059
rect 27120 14028 27261 14056
rect 27120 14016 27126 14028
rect 27249 14025 27261 14028
rect 27295 14025 27307 14059
rect 38010 14056 38016 14068
rect 37971 14028 38016 14056
rect 27249 14019 27307 14025
rect 38010 14016 38016 14028
rect 38068 14016 38074 14068
rect 25041 13991 25099 13997
rect 25041 13957 25053 13991
rect 25087 13957 25099 13991
rect 25041 13951 25099 13957
rect 25130 13948 25136 14000
rect 25188 13988 25194 14000
rect 25188 13960 25233 13988
rect 25188 13948 25194 13960
rect 25682 13948 25688 14000
rect 25740 13988 25746 14000
rect 25869 13991 25927 13997
rect 25869 13988 25881 13991
rect 25740 13960 25881 13988
rect 25740 13948 25746 13960
rect 25869 13957 25881 13960
rect 25915 13957 25927 13991
rect 25869 13951 25927 13957
rect 25961 13991 26019 13997
rect 25961 13957 25973 13991
rect 26007 13988 26019 13991
rect 28442 13988 28448 14000
rect 26007 13960 28448 13988
rect 26007 13957 26019 13960
rect 25961 13951 26019 13957
rect 28442 13948 28448 13960
rect 28500 13948 28506 14000
rect 19150 13920 19156 13932
rect 19111 13892 19156 13920
rect 19150 13880 19156 13892
rect 19208 13920 19214 13932
rect 19797 13923 19855 13929
rect 19797 13920 19809 13923
rect 19208 13892 19809 13920
rect 19208 13880 19214 13892
rect 19797 13889 19809 13892
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 21174 13880 21180 13932
rect 21232 13920 21238 13932
rect 21453 13923 21511 13929
rect 21453 13920 21465 13923
rect 21232 13892 21465 13920
rect 21232 13880 21238 13892
rect 21453 13889 21465 13892
rect 21499 13920 21511 13923
rect 22281 13923 22339 13929
rect 22281 13920 22293 13923
rect 21499 13892 22293 13920
rect 21499 13889 21511 13892
rect 21453 13883 21511 13889
rect 22281 13889 22293 13892
rect 22327 13920 22339 13923
rect 23198 13920 23204 13932
rect 22327 13892 23204 13920
rect 22327 13889 22339 13892
rect 22281 13883 22339 13889
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 23385 13923 23443 13929
rect 23385 13889 23397 13923
rect 23431 13920 23443 13923
rect 23658 13920 23664 13932
rect 23431 13892 23664 13920
rect 23431 13889 23443 13892
rect 23385 13883 23443 13889
rect 23658 13880 23664 13892
rect 23716 13880 23722 13932
rect 24029 13923 24087 13929
rect 24029 13889 24041 13923
rect 24075 13920 24087 13923
rect 26513 13923 26571 13929
rect 24075 13892 24348 13920
rect 24075 13889 24087 13892
rect 24029 13883 24087 13889
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 22370 13852 22376 13864
rect 19291 13824 22376 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 22370 13812 22376 13824
rect 22428 13812 22434 13864
rect 24320 13784 24348 13892
rect 26513 13889 26525 13923
rect 26559 13920 26571 13923
rect 26786 13920 26792 13932
rect 26559 13892 26792 13920
rect 26559 13889 26571 13892
rect 26513 13883 26571 13889
rect 26786 13880 26792 13892
rect 26844 13880 26850 13932
rect 27341 13923 27399 13929
rect 27341 13889 27353 13923
rect 27387 13920 27399 13923
rect 27522 13920 27528 13932
rect 27387 13892 27528 13920
rect 27387 13889 27399 13892
rect 27341 13883 27399 13889
rect 27522 13880 27528 13892
rect 27580 13880 27586 13932
rect 37734 13880 37740 13932
rect 37792 13920 37798 13932
rect 37829 13923 37887 13929
rect 37829 13920 37841 13923
rect 37792 13892 37841 13920
rect 37792 13880 37798 13892
rect 37829 13889 37841 13892
rect 37875 13889 37887 13923
rect 37829 13883 37887 13889
rect 24486 13852 24492 13864
rect 24447 13824 24492 13852
rect 24486 13812 24492 13824
rect 24544 13812 24550 13864
rect 26234 13852 26240 13864
rect 24596 13824 26240 13852
rect 24596 13784 24624 13824
rect 26234 13812 26240 13824
rect 26292 13812 26298 13864
rect 24320 13756 24624 13784
rect 22830 13676 22836 13728
rect 22888 13716 22894 13728
rect 26878 13716 26884 13728
rect 22888 13688 26884 13716
rect 22888 13676 22894 13688
rect 26878 13676 26884 13688
rect 26936 13676 26942 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 23474 13472 23480 13524
rect 23532 13512 23538 13524
rect 23937 13515 23995 13521
rect 23937 13512 23949 13515
rect 23532 13484 23949 13512
rect 23532 13472 23538 13484
rect 23937 13481 23949 13484
rect 23983 13481 23995 13515
rect 23937 13475 23995 13481
rect 25682 13472 25688 13524
rect 25740 13512 25746 13524
rect 26237 13515 26295 13521
rect 26237 13512 26249 13515
rect 25740 13484 26249 13512
rect 25740 13472 25746 13484
rect 26237 13481 26249 13484
rect 26283 13481 26295 13515
rect 26237 13475 26295 13481
rect 26694 13472 26700 13524
rect 26752 13512 26758 13524
rect 26973 13515 27031 13521
rect 26973 13512 26985 13515
rect 26752 13484 26985 13512
rect 26752 13472 26758 13484
rect 26973 13481 26985 13484
rect 27019 13481 27031 13515
rect 26973 13475 27031 13481
rect 22925 13447 22983 13453
rect 22925 13413 22937 13447
rect 22971 13444 22983 13447
rect 24302 13444 24308 13456
rect 22971 13416 24308 13444
rect 22971 13413 22983 13416
rect 22925 13407 22983 13413
rect 24302 13404 24308 13416
rect 24360 13444 24366 13456
rect 24486 13444 24492 13456
rect 24360 13416 24492 13444
rect 24360 13404 24366 13416
rect 24486 13404 24492 13416
rect 24544 13404 24550 13456
rect 22370 13376 22376 13388
rect 22283 13348 22376 13376
rect 22370 13336 22376 13348
rect 22428 13376 22434 13388
rect 23382 13376 23388 13388
rect 22428 13348 23388 13376
rect 22428 13336 22434 13348
rect 23382 13336 23388 13348
rect 23440 13336 23446 13388
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13308 1915 13311
rect 4614 13308 4620 13320
rect 1903 13280 4620 13308
rect 1903 13277 1915 13280
rect 1857 13271 1915 13277
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 10505 13311 10563 13317
rect 10505 13308 10517 13311
rect 6886 13280 10517 13308
rect 1946 13200 1952 13252
rect 2004 13240 2010 13252
rect 6886 13240 6914 13280
rect 10505 13277 10517 13280
rect 10551 13308 10563 13311
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 10551 13280 11161 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 21637 13311 21695 13317
rect 21637 13308 21649 13311
rect 11149 13271 11207 13277
rect 21100 13280 21649 13308
rect 2004 13212 6914 13240
rect 2004 13200 2010 13212
rect 1670 13172 1676 13184
rect 1631 13144 1676 13172
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 10594 13172 10600 13184
rect 10555 13144 10600 13172
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 20898 13132 20904 13184
rect 20956 13172 20962 13184
rect 21100 13181 21128 13280
rect 21637 13277 21649 13280
rect 21683 13277 21695 13311
rect 21637 13271 21695 13277
rect 24029 13311 24087 13317
rect 24029 13277 24041 13311
rect 24075 13277 24087 13311
rect 25774 13308 25780 13320
rect 25735 13280 25780 13308
rect 24029 13271 24087 13277
rect 22465 13243 22523 13249
rect 22465 13209 22477 13243
rect 22511 13209 22523 13243
rect 22465 13203 22523 13209
rect 21085 13175 21143 13181
rect 21085 13172 21097 13175
rect 20956 13144 21097 13172
rect 20956 13132 20962 13144
rect 21085 13141 21097 13144
rect 21131 13141 21143 13175
rect 21085 13135 21143 13141
rect 21729 13175 21787 13181
rect 21729 13141 21741 13175
rect 21775 13172 21787 13175
rect 22480 13172 22508 13203
rect 21775 13144 22508 13172
rect 24044 13172 24072 13271
rect 25774 13268 25780 13280
rect 25832 13268 25838 13320
rect 25958 13308 25964 13320
rect 25919 13280 25964 13308
rect 25958 13268 25964 13280
rect 26016 13268 26022 13320
rect 27065 13311 27123 13317
rect 27065 13277 27077 13311
rect 27111 13308 27123 13311
rect 27246 13308 27252 13320
rect 27111 13280 27252 13308
rect 27111 13277 27123 13280
rect 27065 13271 27123 13277
rect 27246 13268 27252 13280
rect 27304 13268 27310 13320
rect 38010 13308 38016 13320
rect 37971 13280 38016 13308
rect 38010 13268 38016 13280
rect 38068 13268 38074 13320
rect 24578 13240 24584 13252
rect 24539 13212 24584 13240
rect 24578 13200 24584 13212
rect 24636 13200 24642 13252
rect 24762 13200 24768 13252
rect 24820 13240 24826 13252
rect 25133 13243 25191 13249
rect 25133 13240 25145 13243
rect 24820 13212 25145 13240
rect 24820 13200 24826 13212
rect 25133 13209 25145 13212
rect 25179 13209 25191 13243
rect 25133 13203 25191 13209
rect 25222 13200 25228 13252
rect 25280 13240 25286 13252
rect 25280 13212 25325 13240
rect 25280 13200 25286 13212
rect 25866 13172 25872 13184
rect 24044 13144 25872 13172
rect 21775 13141 21787 13144
rect 21729 13135 21787 13141
rect 25866 13132 25872 13144
rect 25924 13132 25930 13184
rect 38194 13172 38200 13184
rect 38155 13144 38200 13172
rect 38194 13132 38200 13144
rect 38252 13132 38258 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 10594 12928 10600 12980
rect 10652 12968 10658 12980
rect 22094 12968 22100 12980
rect 10652 12940 22100 12968
rect 10652 12928 10658 12940
rect 22094 12928 22100 12940
rect 22152 12928 22158 12980
rect 25685 12971 25743 12977
rect 25685 12937 25697 12971
rect 25731 12968 25743 12971
rect 25958 12968 25964 12980
rect 25731 12940 25964 12968
rect 25731 12937 25743 12940
rect 25685 12931 25743 12937
rect 25958 12928 25964 12940
rect 26016 12928 26022 12980
rect 26326 12968 26332 12980
rect 26287 12940 26332 12968
rect 26326 12928 26332 12940
rect 26384 12928 26390 12980
rect 27249 12971 27307 12977
rect 27249 12937 27261 12971
rect 27295 12937 27307 12971
rect 27890 12968 27896 12980
rect 27851 12940 27896 12968
rect 27249 12931 27307 12937
rect 20806 12900 20812 12912
rect 20767 12872 20812 12900
rect 20806 12860 20812 12872
rect 20864 12860 20870 12912
rect 23750 12900 23756 12912
rect 23711 12872 23756 12900
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 24026 12860 24032 12912
rect 24084 12900 24090 12912
rect 24397 12903 24455 12909
rect 24397 12900 24409 12903
rect 24084 12872 24409 12900
rect 24084 12860 24090 12872
rect 24397 12869 24409 12872
rect 24443 12869 24455 12903
rect 24397 12863 24455 12869
rect 24949 12903 25007 12909
rect 24949 12869 24961 12903
rect 24995 12900 25007 12903
rect 27264 12900 27292 12931
rect 27890 12928 27896 12940
rect 27948 12928 27954 12980
rect 29178 12900 29184 12912
rect 24995 12872 27292 12900
rect 28000 12872 29184 12900
rect 24995 12869 25007 12872
rect 24949 12863 25007 12869
rect 22649 12835 22707 12841
rect 22649 12801 22661 12835
rect 22695 12832 22707 12835
rect 22830 12832 22836 12844
rect 22695 12804 22836 12832
rect 22695 12801 22707 12804
rect 22649 12795 22707 12801
rect 20714 12764 20720 12776
rect 20675 12736 20720 12764
rect 20714 12724 20720 12736
rect 20772 12724 20778 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 22278 12764 22284 12776
rect 21407 12736 22284 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 22278 12724 22284 12736
rect 22336 12724 22342 12776
rect 22664 12764 22692 12795
rect 22830 12792 22836 12804
rect 22888 12792 22894 12844
rect 25590 12832 25596 12844
rect 25551 12804 25596 12832
rect 25590 12792 25596 12804
rect 25648 12792 25654 12844
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12801 26479 12835
rect 26421 12795 26479 12801
rect 22572 12736 22692 12764
rect 20165 12631 20223 12637
rect 20165 12597 20177 12631
rect 20211 12628 20223 12631
rect 22094 12628 22100 12640
rect 20211 12600 22100 12628
rect 20211 12597 20223 12600
rect 20165 12591 20223 12597
rect 22094 12588 22100 12600
rect 22152 12628 22158 12640
rect 22572 12628 22600 12736
rect 22922 12724 22928 12776
rect 22980 12764 22986 12776
rect 23201 12767 23259 12773
rect 23201 12764 23213 12767
rect 22980 12736 23213 12764
rect 22980 12724 22986 12736
rect 23201 12733 23213 12736
rect 23247 12733 23259 12767
rect 23201 12727 23259 12733
rect 23845 12767 23903 12773
rect 23845 12733 23857 12767
rect 23891 12733 23903 12767
rect 23845 12727 23903 12733
rect 25041 12767 25099 12773
rect 25041 12733 25053 12767
rect 25087 12733 25099 12767
rect 26436 12764 26464 12795
rect 27246 12792 27252 12844
rect 27304 12832 27310 12844
rect 28000 12841 28028 12872
rect 29178 12860 29184 12872
rect 29236 12860 29242 12912
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 27304 12804 27353 12832
rect 27304 12792 27310 12804
rect 27341 12801 27353 12804
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 27985 12835 28043 12841
rect 27985 12801 27997 12835
rect 28031 12801 28043 12835
rect 27985 12795 28043 12801
rect 28629 12835 28687 12841
rect 28629 12801 28641 12835
rect 28675 12832 28687 12835
rect 28675 12804 29224 12832
rect 28675 12801 28687 12804
rect 28629 12795 28687 12801
rect 27890 12764 27896 12776
rect 26436 12736 27896 12764
rect 25041 12727 25099 12733
rect 22649 12699 22707 12705
rect 22649 12665 22661 12699
rect 22695 12696 22707 12699
rect 23860 12696 23888 12727
rect 22695 12668 23888 12696
rect 25056 12696 25084 12727
rect 27890 12724 27896 12736
rect 27948 12724 27954 12776
rect 25222 12696 25228 12708
rect 25056 12668 25228 12696
rect 22695 12665 22707 12668
rect 22649 12659 22707 12665
rect 25222 12656 25228 12668
rect 25280 12696 25286 12708
rect 26510 12696 26516 12708
rect 25280 12668 26516 12696
rect 25280 12656 25286 12668
rect 26510 12656 26516 12668
rect 26568 12656 26574 12708
rect 22152 12600 22600 12628
rect 22152 12588 22158 12600
rect 27614 12588 27620 12640
rect 27672 12628 27678 12640
rect 29196 12637 29224 12804
rect 28537 12631 28595 12637
rect 28537 12628 28549 12631
rect 27672 12600 28549 12628
rect 27672 12588 27678 12600
rect 28537 12597 28549 12600
rect 28583 12597 28595 12631
rect 28537 12591 28595 12597
rect 29181 12631 29239 12637
rect 29181 12597 29193 12631
rect 29227 12628 29239 12631
rect 37734 12628 37740 12640
rect 29227 12600 37740 12628
rect 29227 12597 29239 12600
rect 29181 12591 29239 12597
rect 37734 12588 37740 12600
rect 37792 12588 37798 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 4341 12427 4399 12433
rect 4341 12393 4353 12427
rect 4387 12424 4399 12427
rect 4614 12424 4620 12436
rect 4387 12396 4620 12424
rect 4387 12393 4399 12396
rect 4341 12387 4399 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 20806 12424 20812 12436
rect 20763 12396 20812 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 22278 12384 22284 12436
rect 22336 12424 22342 12436
rect 28442 12424 28448 12436
rect 22336 12396 26004 12424
rect 28403 12396 28448 12424
rect 22336 12384 22342 12396
rect 6886 12328 23060 12356
rect 2498 12248 2504 12300
rect 2556 12288 2562 12300
rect 6886 12288 6914 12328
rect 2556 12260 6914 12288
rect 17221 12291 17279 12297
rect 2556 12248 2562 12260
rect 17221 12257 17233 12291
rect 17267 12288 17279 12291
rect 20714 12288 20720 12300
rect 17267 12260 20720 12288
rect 17267 12257 17279 12260
rect 17221 12251 17279 12257
rect 20714 12248 20720 12260
rect 20772 12248 20778 12300
rect 22278 12288 22284 12300
rect 22239 12260 22284 12288
rect 22278 12248 22284 12260
rect 22336 12248 22342 12300
rect 23032 12288 23060 12328
rect 23106 12316 23112 12368
rect 23164 12356 23170 12368
rect 23290 12356 23296 12368
rect 23164 12328 23296 12356
rect 23164 12316 23170 12328
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 24946 12288 24952 12300
rect 23032 12260 24952 12288
rect 24946 12248 24952 12260
rect 25004 12248 25010 12300
rect 25976 12297 26004 12396
rect 28442 12384 28448 12396
rect 28500 12384 28506 12436
rect 25961 12291 26019 12297
rect 25961 12257 25973 12291
rect 26007 12288 26019 12291
rect 26513 12291 26571 12297
rect 26513 12288 26525 12291
rect 26007 12260 26525 12288
rect 26007 12257 26019 12260
rect 25961 12251 26019 12257
rect 26513 12257 26525 12260
rect 26559 12257 26571 12291
rect 26513 12251 26571 12257
rect 27157 12291 27215 12297
rect 27157 12257 27169 12291
rect 27203 12288 27215 12291
rect 27614 12288 27620 12300
rect 27203 12260 27620 12288
rect 27203 12257 27215 12260
rect 27157 12251 27215 12257
rect 27614 12248 27620 12260
rect 27672 12248 27678 12300
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4479 12192 5028 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 5000 12096 5028 12192
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 16390 12220 16396 12232
rect 15804 12192 16396 12220
rect 15804 12180 15810 12192
rect 16390 12180 16396 12192
rect 16448 12220 16454 12232
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 16448 12192 17141 12220
rect 16448 12180 16454 12192
rect 17129 12189 17141 12192
rect 17175 12220 17187 12223
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 17175 12192 17785 12220
rect 17175 12189 17187 12192
rect 17129 12183 17187 12189
rect 17773 12189 17785 12192
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12220 20223 12223
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 20211 12192 20637 12220
rect 20211 12189 20223 12192
rect 20165 12183 20223 12189
rect 20625 12189 20637 12192
rect 20671 12220 20683 12223
rect 20806 12220 20812 12232
rect 20671 12192 20812 12220
rect 20671 12189 20683 12192
rect 20625 12183 20683 12189
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 27890 12220 27896 12232
rect 27803 12192 27896 12220
rect 27890 12180 27896 12192
rect 27948 12180 27954 12232
rect 28537 12223 28595 12229
rect 28537 12189 28549 12223
rect 28583 12220 28595 12223
rect 29454 12220 29460 12232
rect 28583 12192 29460 12220
rect 28583 12189 28595 12192
rect 28537 12183 28595 12189
rect 29454 12180 29460 12192
rect 29512 12180 29518 12232
rect 21453 12155 21511 12161
rect 21453 12121 21465 12155
rect 21499 12152 21511 12155
rect 22005 12155 22063 12161
rect 22005 12152 22017 12155
rect 21499 12124 22017 12152
rect 21499 12121 21511 12124
rect 21453 12115 21511 12121
rect 22005 12121 22017 12124
rect 22051 12121 22063 12155
rect 22005 12115 22063 12121
rect 22097 12155 22155 12161
rect 22097 12121 22109 12155
rect 22143 12152 22155 12155
rect 22370 12152 22376 12164
rect 22143 12124 22376 12152
rect 22143 12121 22155 12124
rect 22097 12115 22155 12121
rect 22370 12112 22376 12124
rect 22428 12112 22434 12164
rect 23201 12155 23259 12161
rect 23201 12121 23213 12155
rect 23247 12121 23259 12155
rect 23201 12115 23259 12121
rect 4982 12084 4988 12096
rect 4943 12056 4988 12084
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 22646 12044 22652 12096
rect 22704 12084 22710 12096
rect 23216 12084 23244 12115
rect 23290 12112 23296 12164
rect 23348 12152 23354 12164
rect 23845 12155 23903 12161
rect 23348 12124 23393 12152
rect 23348 12112 23354 12124
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 24118 12152 24124 12164
rect 23891 12124 24124 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 24118 12112 24124 12124
rect 24176 12152 24182 12164
rect 24578 12152 24584 12164
rect 24176 12124 24584 12152
rect 24176 12112 24182 12124
rect 24578 12112 24584 12124
rect 24636 12112 24642 12164
rect 25682 12112 25688 12164
rect 25740 12152 25746 12164
rect 25869 12155 25927 12161
rect 25869 12152 25881 12155
rect 25740 12124 25881 12152
rect 25740 12112 25746 12124
rect 25869 12121 25881 12124
rect 25915 12121 25927 12155
rect 25869 12115 25927 12121
rect 27065 12155 27123 12161
rect 27065 12121 27077 12155
rect 27111 12121 27123 12155
rect 27908 12152 27936 12180
rect 29086 12152 29092 12164
rect 27908 12124 29092 12152
rect 27065 12115 27123 12121
rect 22704 12056 23244 12084
rect 27080 12084 27108 12115
rect 29086 12112 29092 12124
rect 29144 12112 29150 12164
rect 27801 12087 27859 12093
rect 27801 12084 27813 12087
rect 27080 12056 27813 12084
rect 22704 12044 22710 12056
rect 27801 12053 27813 12056
rect 27847 12053 27859 12087
rect 27801 12047 27859 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 22094 11880 22100 11892
rect 22020 11852 22100 11880
rect 20809 11747 20867 11753
rect 20809 11713 20821 11747
rect 20855 11744 20867 11747
rect 21453 11747 21511 11753
rect 21453 11744 21465 11747
rect 20855 11716 21465 11744
rect 20855 11713 20867 11716
rect 20809 11707 20867 11713
rect 21453 11713 21465 11716
rect 21499 11744 21511 11747
rect 22020 11744 22048 11852
rect 22094 11840 22100 11852
rect 22152 11840 22158 11892
rect 25774 11840 25780 11892
rect 25832 11880 25838 11892
rect 26053 11883 26111 11889
rect 26053 11880 26065 11883
rect 25832 11852 26065 11880
rect 25832 11840 25838 11852
rect 26053 11849 26065 11852
rect 26099 11849 26111 11883
rect 26053 11843 26111 11849
rect 26510 11840 26516 11892
rect 26568 11880 26574 11892
rect 27249 11883 27307 11889
rect 27249 11880 27261 11883
rect 26568 11852 27261 11880
rect 26568 11840 26574 11852
rect 27249 11849 27261 11852
rect 27295 11849 27307 11883
rect 27249 11843 27307 11849
rect 22186 11812 22192 11824
rect 22147 11784 22192 11812
rect 22186 11772 22192 11784
rect 22244 11772 22250 11824
rect 22281 11815 22339 11821
rect 22281 11781 22293 11815
rect 22327 11812 22339 11815
rect 23014 11812 23020 11824
rect 22327 11784 23020 11812
rect 22327 11781 22339 11784
rect 22281 11775 22339 11781
rect 23014 11772 23020 11784
rect 23072 11772 23078 11824
rect 24026 11772 24032 11824
rect 24084 11812 24090 11824
rect 24489 11815 24547 11821
rect 24489 11812 24501 11815
rect 24084 11784 24501 11812
rect 24084 11772 24090 11784
rect 24489 11781 24501 11784
rect 24535 11781 24547 11815
rect 24489 11775 24547 11781
rect 24578 11772 24584 11824
rect 24636 11812 24642 11824
rect 24636 11784 24681 11812
rect 24636 11772 24642 11784
rect 25866 11772 25872 11824
rect 25924 11812 25930 11824
rect 25924 11784 27844 11812
rect 25924 11772 25930 11784
rect 21499 11716 22048 11744
rect 23293 11747 23351 11753
rect 21499 11713 21511 11716
rect 21453 11707 21511 11713
rect 23293 11713 23305 11747
rect 23339 11713 23351 11747
rect 23293 11707 23351 11713
rect 26145 11747 26203 11753
rect 26145 11713 26157 11747
rect 26191 11744 26203 11747
rect 27062 11744 27068 11756
rect 26191 11716 27068 11744
rect 26191 11713 26203 11716
rect 26145 11707 26203 11713
rect 23308 11676 23336 11707
rect 24854 11676 24860 11688
rect 22066 11648 23336 11676
rect 24815 11648 24860 11676
rect 19978 11568 19984 11620
rect 20036 11608 20042 11620
rect 20036 11580 21404 11608
rect 20036 11568 20042 11580
rect 21174 11500 21180 11552
rect 21232 11540 21238 11552
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 21232 11512 21281 11540
rect 21232 11500 21238 11512
rect 21269 11509 21281 11512
rect 21315 11509 21327 11543
rect 21376 11540 21404 11580
rect 21542 11568 21548 11620
rect 21600 11608 21606 11620
rect 22066 11608 22094 11648
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 25130 11636 25136 11688
rect 25188 11676 25194 11688
rect 26160 11676 26188 11707
rect 27062 11704 27068 11716
rect 27120 11704 27126 11756
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11744 27399 11747
rect 27430 11744 27436 11756
rect 27387 11716 27436 11744
rect 27387 11713 27399 11716
rect 27341 11707 27399 11713
rect 27430 11704 27436 11716
rect 27488 11704 27494 11756
rect 27816 11753 27844 11784
rect 27801 11747 27859 11753
rect 27801 11713 27813 11747
rect 27847 11713 27859 11747
rect 27801 11707 27859 11713
rect 25188 11648 26188 11676
rect 26620 11648 31754 11676
rect 25188 11636 25194 11648
rect 21600 11580 22094 11608
rect 21600 11568 21606 11580
rect 22646 11568 22652 11620
rect 22704 11608 22710 11620
rect 22741 11611 22799 11617
rect 22741 11608 22753 11611
rect 22704 11580 22753 11608
rect 22704 11568 22710 11580
rect 22741 11577 22753 11580
rect 22787 11608 22799 11611
rect 22922 11608 22928 11620
rect 22787 11580 22928 11608
rect 22787 11577 22799 11580
rect 22741 11571 22799 11577
rect 22922 11568 22928 11580
rect 22980 11568 22986 11620
rect 23477 11611 23535 11617
rect 23477 11577 23489 11611
rect 23523 11608 23535 11611
rect 26620 11608 26648 11648
rect 23523 11580 26648 11608
rect 23523 11577 23535 11580
rect 23477 11571 23535 11577
rect 26694 11568 26700 11620
rect 26752 11608 26758 11620
rect 27893 11611 27951 11617
rect 27893 11608 27905 11611
rect 26752 11580 27905 11608
rect 26752 11568 26758 11580
rect 27893 11577 27905 11580
rect 27939 11577 27951 11611
rect 31726 11608 31754 11648
rect 38010 11608 38016 11620
rect 31726 11580 38016 11608
rect 27893 11571 27951 11577
rect 38010 11568 38016 11580
rect 38068 11568 38074 11620
rect 26786 11540 26792 11552
rect 21376 11512 26792 11540
rect 21269 11503 21327 11509
rect 26786 11500 26792 11512
rect 26844 11500 26850 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 16390 11336 16396 11348
rect 5040 11308 6914 11336
rect 16351 11308 16396 11336
rect 5040 11296 5046 11308
rect 6886 11268 6914 11308
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 22370 11336 22376 11348
rect 22331 11308 22376 11336
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 23014 11336 23020 11348
rect 22975 11308 23020 11336
rect 23014 11296 23020 11308
rect 23072 11296 23078 11348
rect 23661 11339 23719 11345
rect 23661 11305 23673 11339
rect 23707 11336 23719 11339
rect 23750 11336 23756 11348
rect 23707 11308 23756 11336
rect 23707 11305 23719 11308
rect 23661 11299 23719 11305
rect 23750 11296 23756 11308
rect 23808 11296 23814 11348
rect 24854 11268 24860 11280
rect 6886 11240 24860 11268
rect 24854 11228 24860 11240
rect 24912 11228 24918 11280
rect 24946 11200 24952 11212
rect 24907 11172 24952 11200
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 26418 11200 26424 11212
rect 26379 11172 26424 11200
rect 26418 11160 26424 11172
rect 26476 11160 26482 11212
rect 26786 11160 26792 11212
rect 26844 11200 26850 11212
rect 38013 11203 38071 11209
rect 38013 11200 38025 11203
rect 26844 11172 38025 11200
rect 26844 11160 26850 11172
rect 38013 11169 38025 11172
rect 38059 11169 38071 11203
rect 38013 11163 38071 11169
rect 1762 11092 1768 11144
rect 1820 11132 1826 11144
rect 1857 11135 1915 11141
rect 1857 11132 1869 11135
rect 1820 11104 1869 11132
rect 1820 11092 1826 11104
rect 1857 11101 1869 11104
rect 1903 11101 1915 11135
rect 1857 11095 1915 11101
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11132 15807 11135
rect 16390 11132 16396 11144
rect 15795 11104 16396 11132
rect 15795 11101 15807 11104
rect 15749 11095 15807 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 21085 11135 21143 11141
rect 21085 11101 21097 11135
rect 21131 11132 21143 11135
rect 21542 11132 21548 11144
rect 21131 11104 21548 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 21542 11092 21548 11104
rect 21600 11092 21606 11144
rect 22094 11092 22100 11144
rect 22152 11132 22158 11144
rect 22465 11135 22523 11141
rect 22465 11132 22477 11135
rect 22152 11104 22477 11132
rect 22152 11092 22158 11104
rect 22465 11101 22477 11104
rect 22511 11101 22523 11135
rect 22465 11095 22523 11101
rect 23109 11135 23167 11141
rect 23109 11101 23121 11135
rect 23155 11132 23167 11135
rect 23474 11132 23480 11144
rect 23155 11104 23480 11132
rect 23155 11101 23167 11104
rect 23109 11095 23167 11101
rect 23474 11092 23480 11104
rect 23532 11092 23538 11144
rect 23753 11135 23811 11141
rect 23753 11101 23765 11135
rect 23799 11132 23811 11135
rect 24210 11132 24216 11144
rect 23799 11104 24216 11132
rect 23799 11101 23811 11104
rect 23753 11095 23811 11101
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 27062 11092 27068 11144
rect 27120 11132 27126 11144
rect 27341 11135 27399 11141
rect 27341 11132 27353 11135
rect 27120 11104 27353 11132
rect 27120 11092 27126 11104
rect 27341 11101 27353 11104
rect 27387 11132 27399 11135
rect 31478 11132 31484 11144
rect 27387 11104 31484 11132
rect 27387 11101 27399 11104
rect 27341 11095 27399 11101
rect 31478 11092 31484 11104
rect 31536 11092 31542 11144
rect 38286 11132 38292 11144
rect 38247 11104 38292 11132
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 21821 11067 21879 11073
rect 21821 11033 21833 11067
rect 21867 11064 21879 11067
rect 21910 11064 21916 11076
rect 21867 11036 21916 11064
rect 21867 11033 21879 11036
rect 21821 11027 21879 11033
rect 21910 11024 21916 11036
rect 21968 11024 21974 11076
rect 24302 11024 24308 11076
rect 24360 11064 24366 11076
rect 24670 11064 24676 11076
rect 24360 11036 24676 11064
rect 24360 11024 24366 11036
rect 24670 11024 24676 11036
rect 24728 11024 24734 11076
rect 24765 11067 24823 11073
rect 24765 11033 24777 11067
rect 24811 11033 24823 11067
rect 26694 11064 26700 11076
rect 26655 11036 26700 11064
rect 24765 11027 24823 11033
rect 1670 10996 1676 11008
rect 1631 10968 1676 10996
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 15930 10996 15936 11008
rect 15891 10968 15936 10996
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 24486 10956 24492 11008
rect 24544 10996 24550 11008
rect 24780 10996 24808 11027
rect 26694 11024 26700 11036
rect 26752 11024 26758 11076
rect 26786 11024 26792 11076
rect 26844 11064 26850 11076
rect 26844 11036 26889 11064
rect 26844 11024 26850 11036
rect 27430 11024 27436 11076
rect 27488 11064 27494 11076
rect 27985 11067 28043 11073
rect 27985 11064 27997 11067
rect 27488 11036 27997 11064
rect 27488 11024 27494 11036
rect 27985 11033 27997 11036
rect 28031 11064 28043 11067
rect 38102 11064 38108 11076
rect 28031 11036 38108 11064
rect 28031 11033 28043 11036
rect 27985 11027 28043 11033
rect 38102 11024 38108 11036
rect 38160 11024 38166 11076
rect 24544 10968 24808 10996
rect 24544 10956 24550 10968
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 23290 10792 23296 10804
rect 23251 10764 23296 10792
rect 23290 10752 23296 10764
rect 23348 10752 23354 10804
rect 24213 10795 24271 10801
rect 24213 10761 24225 10795
rect 24259 10792 24271 10795
rect 24762 10792 24768 10804
rect 24259 10764 24768 10792
rect 24259 10761 24271 10764
rect 24213 10755 24271 10761
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 24854 10752 24860 10804
rect 24912 10792 24918 10804
rect 25314 10792 25320 10804
rect 24912 10764 25320 10792
rect 24912 10752 24918 10764
rect 25314 10752 25320 10764
rect 25372 10792 25378 10804
rect 36262 10792 36268 10804
rect 25372 10764 26188 10792
rect 36223 10764 36268 10792
rect 25372 10752 25378 10764
rect 2041 10727 2099 10733
rect 2041 10693 2053 10727
rect 2087 10724 2099 10727
rect 2406 10724 2412 10736
rect 2087 10696 2412 10724
rect 2087 10693 2099 10696
rect 2041 10687 2099 10693
rect 2406 10684 2412 10696
rect 2464 10684 2470 10736
rect 15749 10727 15807 10733
rect 15749 10693 15761 10727
rect 15795 10724 15807 10727
rect 17218 10724 17224 10736
rect 15795 10696 17224 10724
rect 15795 10693 15807 10696
rect 15749 10687 15807 10693
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 21910 10684 21916 10736
rect 21968 10724 21974 10736
rect 22086 10727 22144 10733
rect 22086 10724 22098 10727
rect 21968 10696 22098 10724
rect 21968 10684 21974 10696
rect 22086 10693 22098 10696
rect 22132 10693 22144 10727
rect 22086 10687 22144 10693
rect 22186 10684 22192 10736
rect 22244 10724 22250 10736
rect 25406 10724 25412 10736
rect 22244 10696 22289 10724
rect 25367 10696 25412 10724
rect 22244 10684 22250 10696
rect 25406 10684 25412 10696
rect 25464 10684 25470 10736
rect 26160 10724 26188 10764
rect 36262 10752 36268 10764
rect 36320 10752 36326 10804
rect 38286 10792 38292 10804
rect 38247 10764 38292 10792
rect 38286 10752 38292 10764
rect 38344 10752 38350 10804
rect 26329 10727 26387 10733
rect 26329 10724 26341 10727
rect 26160 10696 26341 10724
rect 26329 10693 26341 10696
rect 26375 10693 26387 10727
rect 26329 10687 26387 10693
rect 29181 10727 29239 10733
rect 29181 10693 29193 10727
rect 29227 10724 29239 10727
rect 31205 10727 31263 10733
rect 31205 10724 31217 10727
rect 29227 10696 31217 10724
rect 29227 10693 29239 10696
rect 29181 10687 29239 10693
rect 31205 10693 31217 10696
rect 31251 10693 31263 10727
rect 31205 10687 31263 10693
rect 1854 10656 1860 10668
rect 1767 10628 1860 10656
rect 1854 10616 1860 10628
rect 1912 10656 1918 10668
rect 14274 10656 14280 10668
rect 1912 10628 14280 10656
rect 1912 10616 1918 10628
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 21358 10656 21364 10668
rect 21319 10628 21364 10656
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10625 21511 10659
rect 21453 10619 21511 10625
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 15657 10591 15715 10597
rect 15657 10588 15669 10591
rect 14424 10560 15669 10588
rect 14424 10548 14430 10560
rect 15657 10557 15669 10560
rect 15703 10557 15715 10591
rect 21468 10588 21496 10619
rect 22738 10616 22744 10668
rect 22796 10656 22802 10668
rect 23385 10659 23443 10665
rect 23385 10656 23397 10659
rect 22796 10628 23397 10656
rect 22796 10616 22802 10628
rect 23385 10625 23397 10628
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10656 24179 10659
rect 24210 10656 24216 10668
rect 24167 10628 24216 10656
rect 24167 10625 24179 10628
rect 24121 10619 24179 10625
rect 24210 10616 24216 10628
rect 24268 10616 24274 10668
rect 26418 10656 26424 10668
rect 26160 10628 26424 10656
rect 22094 10588 22100 10600
rect 21468 10560 22100 10588
rect 15657 10551 15715 10557
rect 22094 10548 22100 10560
rect 22152 10548 22158 10600
rect 25317 10591 25375 10597
rect 25317 10557 25329 10591
rect 25363 10588 25375 10591
rect 26160 10588 26188 10628
rect 26418 10616 26424 10628
rect 26476 10616 26482 10668
rect 29086 10656 29092 10668
rect 28999 10628 29092 10656
rect 29086 10616 29092 10628
rect 29144 10656 29150 10668
rect 29546 10656 29552 10668
rect 29144 10628 29552 10656
rect 29144 10616 29150 10628
rect 29546 10616 29552 10628
rect 29604 10616 29610 10668
rect 36170 10656 36176 10668
rect 36131 10628 36176 10656
rect 36170 10616 36176 10628
rect 36228 10616 36234 10668
rect 25363 10560 26188 10588
rect 31297 10591 31355 10597
rect 25363 10557 25375 10560
rect 25317 10551 25375 10557
rect 31297 10557 31309 10591
rect 31343 10588 31355 10591
rect 33594 10588 33600 10600
rect 31343 10560 33600 10588
rect 31343 10557 31355 10560
rect 31297 10551 31355 10557
rect 33594 10548 33600 10560
rect 33652 10548 33658 10600
rect 16209 10523 16267 10529
rect 16209 10489 16221 10523
rect 16255 10520 16267 10523
rect 22649 10523 22707 10529
rect 22649 10520 22661 10523
rect 16255 10492 22661 10520
rect 16255 10489 16267 10492
rect 16209 10483 16267 10489
rect 22649 10489 22661 10492
rect 22695 10520 22707 10523
rect 26602 10520 26608 10532
rect 22695 10492 26608 10520
rect 22695 10489 22707 10492
rect 22649 10483 22707 10489
rect 26602 10480 26608 10492
rect 26660 10520 26666 10532
rect 30745 10523 30803 10529
rect 30745 10520 30757 10523
rect 26660 10492 30757 10520
rect 26660 10480 26666 10492
rect 30745 10489 30757 10492
rect 30791 10489 30803 10523
rect 30745 10483 30803 10489
rect 20806 10412 20812 10464
rect 20864 10452 20870 10464
rect 27798 10452 27804 10464
rect 20864 10424 27804 10452
rect 20864 10412 20870 10424
rect 27798 10412 27804 10424
rect 27856 10412 27862 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 17218 10248 17224 10260
rect 17179 10220 17224 10248
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 17865 10251 17923 10257
rect 17865 10217 17877 10251
rect 17911 10248 17923 10251
rect 20806 10248 20812 10260
rect 17911 10220 20812 10248
rect 17911 10217 17923 10220
rect 17865 10211 17923 10217
rect 1854 10112 1860 10124
rect 1815 10084 1860 10112
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 14274 10044 14280 10056
rect 14235 10016 14280 10044
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 17880 10044 17908 10211
rect 20806 10208 20812 10220
rect 20864 10208 20870 10260
rect 33594 10248 33600 10260
rect 33555 10220 33600 10248
rect 33594 10208 33600 10220
rect 33652 10208 33658 10260
rect 21542 10140 21548 10192
rect 21600 10180 21606 10192
rect 23385 10183 23443 10189
rect 23385 10180 23397 10183
rect 21600 10152 23397 10180
rect 21600 10140 21606 10152
rect 23385 10149 23397 10152
rect 23431 10149 23443 10183
rect 27062 10180 27068 10192
rect 23385 10143 23443 10149
rect 24780 10152 27068 10180
rect 22925 10115 22983 10121
rect 22925 10081 22937 10115
rect 22971 10112 22983 10115
rect 24670 10112 24676 10124
rect 22971 10084 24676 10112
rect 22971 10081 22983 10084
rect 22925 10075 22983 10081
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 17359 10016 17908 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 23474 10004 23480 10056
rect 23532 10044 23538 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 23532 10016 24593 10044
rect 23532 10004 23538 10016
rect 24581 10013 24593 10016
rect 24627 10044 24639 10047
rect 24780 10044 24808 10152
rect 27062 10140 27068 10152
rect 27120 10140 27126 10192
rect 24946 10072 24952 10124
rect 25004 10112 25010 10124
rect 25593 10115 25651 10121
rect 25593 10112 25605 10115
rect 25004 10084 25605 10112
rect 25004 10072 25010 10084
rect 25593 10081 25605 10084
rect 25639 10081 25651 10115
rect 26602 10112 26608 10124
rect 26563 10084 26608 10112
rect 25593 10075 25651 10081
rect 26602 10072 26608 10084
rect 26660 10072 26666 10124
rect 24627 10016 24808 10044
rect 27341 10047 27399 10053
rect 24627 10013 24639 10016
rect 24581 10007 24639 10013
rect 27341 10013 27353 10047
rect 27387 10044 27399 10047
rect 29086 10044 29092 10056
rect 27387 10016 29092 10044
rect 27387 10013 27399 10016
rect 27341 10007 27399 10013
rect 29086 10004 29092 10016
rect 29144 10004 29150 10056
rect 33689 10047 33747 10053
rect 33689 10013 33701 10047
rect 33735 10044 33747 10047
rect 36170 10044 36176 10056
rect 33735 10016 36176 10044
rect 33735 10013 33747 10016
rect 33689 10007 33747 10013
rect 36170 10004 36176 10016
rect 36228 10004 36234 10056
rect 22278 9976 22284 9988
rect 22239 9948 22284 9976
rect 22278 9936 22284 9948
rect 22336 9936 22342 9988
rect 22370 9936 22376 9988
rect 22428 9976 22434 9988
rect 26510 9976 26516 9988
rect 22428 9948 22473 9976
rect 26471 9948 26516 9976
rect 22428 9936 22434 9948
rect 26510 9936 26516 9948
rect 26568 9936 26574 9988
rect 24670 9908 24676 9920
rect 24631 9880 24676 9908
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 26234 9868 26240 9920
rect 26292 9908 26298 9920
rect 27249 9911 27307 9917
rect 27249 9908 27261 9911
rect 26292 9880 27261 9908
rect 26292 9868 26298 9880
rect 27249 9877 27261 9880
rect 27295 9877 27307 9911
rect 27249 9871 27307 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 22281 9707 22339 9713
rect 22281 9673 22293 9707
rect 22327 9704 22339 9707
rect 22370 9704 22376 9716
rect 22327 9676 22376 9704
rect 22327 9673 22339 9676
rect 22281 9667 22339 9673
rect 22370 9664 22376 9676
rect 22428 9664 22434 9716
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 24670 9636 24676 9648
rect 24631 9608 24676 9636
rect 24670 9596 24676 9608
rect 24728 9596 24734 9648
rect 25314 9636 25320 9648
rect 25275 9608 25320 9636
rect 25314 9596 25320 9608
rect 25372 9596 25378 9648
rect 26234 9636 26240 9648
rect 26195 9608 26240 9636
rect 26234 9596 26240 9608
rect 26292 9596 26298 9648
rect 22094 9528 22100 9580
rect 22152 9568 22158 9580
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 22152 9540 22201 9568
rect 22152 9528 22158 9540
rect 22189 9537 22201 9540
rect 22235 9568 22247 9571
rect 23290 9568 23296 9580
rect 22235 9540 23296 9568
rect 22235 9537 22247 9540
rect 22189 9531 22247 9537
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 24118 9500 24124 9512
rect 24079 9472 24124 9500
rect 24118 9460 24124 9472
rect 24176 9460 24182 9512
rect 24765 9503 24823 9509
rect 24765 9469 24777 9503
rect 24811 9469 24823 9503
rect 26326 9500 26332 9512
rect 26287 9472 26332 9500
rect 24765 9463 24823 9469
rect 24780 9432 24808 9463
rect 26326 9460 26332 9472
rect 26384 9460 26390 9512
rect 25038 9432 25044 9444
rect 24780 9404 25044 9432
rect 25038 9392 25044 9404
rect 25096 9432 25102 9444
rect 26786 9432 26792 9444
rect 25096 9404 26792 9432
rect 25096 9392 25102 9404
rect 26786 9392 26792 9404
rect 26844 9392 26850 9444
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 20901 9163 20959 9169
rect 20901 9129 20913 9163
rect 20947 9160 20959 9163
rect 22278 9160 22284 9172
rect 20947 9132 22284 9160
rect 20947 9129 20959 9132
rect 20901 9123 20959 9129
rect 22278 9120 22284 9132
rect 22336 9120 22342 9172
rect 23477 9163 23535 9169
rect 23477 9129 23489 9163
rect 23523 9160 23535 9163
rect 24486 9160 24492 9172
rect 23523 9132 24492 9160
rect 23523 9129 23535 9132
rect 23477 9123 23535 9129
rect 24486 9120 24492 9132
rect 24544 9120 24550 9172
rect 25038 9160 25044 9172
rect 24999 9132 25044 9160
rect 25038 9120 25044 9132
rect 25096 9120 25102 9172
rect 37826 9160 37832 9172
rect 25148 9132 37832 9160
rect 22097 9027 22155 9033
rect 22097 8993 22109 9027
rect 22143 9024 22155 9027
rect 24118 9024 24124 9036
rect 22143 8996 24124 9024
rect 22143 8993 22155 8996
rect 22097 8987 22155 8993
rect 24118 8984 24124 8996
rect 24176 8984 24182 9036
rect 20806 8956 20812 8968
rect 20767 8928 20812 8956
rect 20806 8916 20812 8928
rect 20864 8916 20870 8968
rect 23569 8959 23627 8965
rect 23569 8925 23581 8959
rect 23615 8956 23627 8959
rect 24854 8956 24860 8968
rect 23615 8928 24860 8956
rect 23615 8925 23627 8928
rect 23569 8919 23627 8925
rect 24854 8916 24860 8928
rect 24912 8916 24918 8968
rect 25148 8965 25176 9132
rect 37826 9120 37832 9132
rect 37884 9120 37890 9172
rect 38102 9160 38108 9172
rect 38063 9132 38108 9160
rect 38102 9120 38108 9132
rect 38160 9120 38166 9172
rect 25682 9092 25688 9104
rect 25643 9064 25688 9092
rect 25682 9052 25688 9064
rect 25740 9052 25746 9104
rect 26326 8984 26332 9036
rect 26384 9024 26390 9036
rect 26421 9027 26479 9033
rect 26421 9024 26433 9027
rect 26384 8996 26433 9024
rect 26384 8984 26390 8996
rect 26421 8993 26433 8996
rect 26467 8993 26479 9027
rect 26421 8987 26479 8993
rect 25133 8959 25191 8965
rect 25133 8925 25145 8959
rect 25179 8925 25191 8959
rect 25133 8919 25191 8925
rect 25777 8959 25835 8965
rect 25777 8925 25789 8959
rect 25823 8956 25835 8959
rect 28810 8956 28816 8968
rect 25823 8928 28816 8956
rect 25823 8925 25835 8928
rect 25777 8919 25835 8925
rect 28810 8916 28816 8928
rect 28868 8916 28874 8968
rect 29362 8916 29368 8968
rect 29420 8956 29426 8968
rect 30745 8959 30803 8965
rect 30745 8956 30757 8959
rect 29420 8928 30757 8956
rect 29420 8916 29426 8928
rect 30745 8925 30757 8928
rect 30791 8925 30803 8959
rect 30745 8919 30803 8925
rect 21450 8888 21456 8900
rect 21411 8860 21456 8888
rect 21450 8848 21456 8860
rect 21508 8848 21514 8900
rect 22005 8891 22063 8897
rect 22005 8857 22017 8891
rect 22051 8857 22063 8891
rect 22005 8851 22063 8857
rect 22020 8820 22048 8851
rect 28534 8848 28540 8900
rect 28592 8888 28598 8900
rect 30466 8888 30472 8900
rect 28592 8860 30472 8888
rect 28592 8848 28598 8860
rect 30466 8848 30472 8860
rect 30524 8848 30530 8900
rect 37553 8891 37611 8897
rect 37553 8857 37565 8891
rect 37599 8888 37611 8891
rect 38194 8888 38200 8900
rect 37599 8860 38200 8888
rect 37599 8857 37611 8860
rect 37553 8851 37611 8857
rect 38194 8848 38200 8860
rect 38252 8848 38258 8900
rect 22462 8820 22468 8832
rect 22020 8792 22468 8820
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 27246 8820 27252 8832
rect 27207 8792 27252 8820
rect 27246 8780 27252 8792
rect 27304 8780 27310 8832
rect 29270 8780 29276 8832
rect 29328 8820 29334 8832
rect 29825 8823 29883 8829
rect 29825 8820 29837 8823
rect 29328 8792 29837 8820
rect 29328 8780 29334 8792
rect 29825 8789 29837 8792
rect 29871 8820 29883 8823
rect 30926 8820 30932 8832
rect 29871 8792 30932 8820
rect 29871 8789 29883 8792
rect 29825 8783 29883 8789
rect 30926 8780 30932 8792
rect 30984 8780 30990 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 25406 8616 25412 8628
rect 25367 8588 25412 8616
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 26053 8619 26111 8625
rect 26053 8585 26065 8619
rect 26099 8616 26111 8619
rect 26510 8616 26516 8628
rect 26099 8588 26516 8616
rect 26099 8585 26111 8588
rect 26053 8579 26111 8585
rect 26510 8576 26516 8588
rect 26568 8576 26574 8628
rect 27062 8576 27068 8628
rect 27120 8616 27126 8628
rect 27525 8619 27583 8625
rect 27525 8616 27537 8619
rect 27120 8588 27537 8616
rect 27120 8576 27126 8588
rect 27525 8585 27537 8588
rect 27571 8585 27583 8619
rect 27525 8579 27583 8585
rect 27632 8588 29224 8616
rect 22186 8508 22192 8560
rect 22244 8548 22250 8560
rect 22281 8551 22339 8557
rect 22281 8548 22293 8551
rect 22244 8520 22293 8548
rect 22244 8508 22250 8520
rect 22281 8517 22293 8520
rect 22327 8517 22339 8551
rect 22281 8511 22339 8517
rect 23290 8508 23296 8560
rect 23348 8548 23354 8560
rect 23385 8551 23443 8557
rect 23385 8548 23397 8551
rect 23348 8520 23397 8548
rect 23348 8508 23354 8520
rect 23385 8517 23397 8520
rect 23431 8517 23443 8551
rect 27632 8548 27660 8588
rect 23385 8511 23443 8517
rect 26252 8520 27660 8548
rect 22373 8483 22431 8489
rect 22373 8449 22385 8483
rect 22419 8480 22431 8483
rect 22738 8480 22744 8492
rect 22419 8452 22744 8480
rect 22419 8449 22431 8452
rect 22373 8443 22431 8449
rect 22738 8440 22744 8452
rect 22796 8440 22802 8492
rect 25501 8483 25559 8489
rect 22278 8372 22284 8424
rect 22336 8412 22342 8424
rect 23109 8415 23167 8421
rect 23109 8412 23121 8415
rect 22336 8384 23121 8412
rect 22336 8372 22342 8384
rect 23109 8381 23121 8384
rect 23155 8381 23167 8415
rect 23109 8375 23167 8381
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 20806 8344 20812 8356
rect 19300 8316 20812 8344
rect 19300 8304 19306 8316
rect 20806 8304 20812 8316
rect 20864 8344 20870 8356
rect 21085 8347 21143 8353
rect 21085 8344 21097 8347
rect 20864 8316 21097 8344
rect 20864 8304 20870 8316
rect 21085 8313 21097 8316
rect 21131 8313 21143 8347
rect 24504 8344 24532 8466
rect 25501 8449 25513 8483
rect 25547 8480 25559 8483
rect 26050 8480 26056 8492
rect 25547 8452 26056 8480
rect 25547 8449 25559 8452
rect 25501 8443 25559 8449
rect 26050 8440 26056 8452
rect 26108 8440 26114 8492
rect 26145 8483 26203 8489
rect 26145 8449 26157 8483
rect 26191 8480 26203 8483
rect 26252 8480 26280 8520
rect 28534 8508 28540 8560
rect 28592 8508 28598 8560
rect 28997 8551 29055 8557
rect 28997 8517 29009 8551
rect 29043 8548 29055 8551
rect 29086 8548 29092 8560
rect 29043 8520 29092 8548
rect 29043 8517 29055 8520
rect 28997 8511 29055 8517
rect 29086 8508 29092 8520
rect 29144 8508 29150 8560
rect 29196 8548 29224 8588
rect 29196 8520 29684 8548
rect 26191 8452 26280 8480
rect 26191 8449 26203 8452
rect 26145 8443 26203 8449
rect 29270 8440 29276 8492
rect 29328 8480 29334 8492
rect 29328 8452 29373 8480
rect 29328 8440 29334 8452
rect 24854 8412 24860 8424
rect 24767 8384 24860 8412
rect 24854 8372 24860 8384
rect 24912 8412 24918 8424
rect 28902 8412 28908 8424
rect 24912 8384 28908 8412
rect 24912 8372 24918 8384
rect 28902 8372 28908 8384
rect 28960 8372 28966 8424
rect 29656 8412 29684 8520
rect 30926 8508 30932 8560
rect 30984 8548 30990 8560
rect 30984 8520 31524 8548
rect 30984 8508 30990 8520
rect 30098 8440 30104 8492
rect 30156 8440 30162 8492
rect 31496 8489 31524 8520
rect 31481 8483 31539 8489
rect 31481 8449 31493 8483
rect 31527 8449 31539 8483
rect 31481 8443 31539 8449
rect 31202 8412 31208 8424
rect 29656 8384 31208 8412
rect 31202 8372 31208 8384
rect 31260 8372 31266 8424
rect 27430 8344 27436 8356
rect 24504 8316 27436 8344
rect 21085 8307 21143 8313
rect 27430 8304 27436 8316
rect 27488 8304 27494 8356
rect 29733 8347 29791 8353
rect 29733 8344 29745 8347
rect 29196 8316 29745 8344
rect 28810 8236 28816 8288
rect 28868 8276 28874 8288
rect 29196 8276 29224 8316
rect 29733 8313 29745 8316
rect 29779 8313 29791 8347
rect 29733 8307 29791 8313
rect 28868 8248 29224 8276
rect 28868 8236 28874 8248
rect 30006 8236 30012 8288
rect 30064 8276 30070 8288
rect 32122 8276 32128 8288
rect 30064 8248 32128 8276
rect 30064 8236 30070 8248
rect 32122 8236 32128 8248
rect 32180 8236 32186 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 23290 8032 23296 8084
rect 23348 8072 23354 8084
rect 23348 8044 23612 8072
rect 23348 8032 23354 8044
rect 23584 8004 23612 8044
rect 24578 8032 24584 8084
rect 24636 8072 24642 8084
rect 24673 8075 24731 8081
rect 24673 8072 24685 8075
rect 24636 8044 24685 8072
rect 24636 8032 24642 8044
rect 24673 8041 24685 8044
rect 24719 8041 24731 8075
rect 24673 8035 24731 8041
rect 26510 8032 26516 8084
rect 26568 8072 26574 8084
rect 26568 8044 31064 8072
rect 26568 8032 26574 8044
rect 25501 8007 25559 8013
rect 25501 8004 25513 8007
rect 23584 7976 25513 8004
rect 25501 7973 25513 7976
rect 25547 7973 25559 8007
rect 25501 7967 25559 7973
rect 27522 7964 27528 8016
rect 27580 8004 27586 8016
rect 29546 8004 29552 8016
rect 27580 7976 29552 8004
rect 27580 7964 27586 7976
rect 29546 7964 29552 7976
rect 29604 7964 29610 8016
rect 31036 8004 31064 8044
rect 31202 8032 31208 8084
rect 31260 8072 31266 8084
rect 31481 8075 31539 8081
rect 31481 8072 31493 8075
rect 31260 8044 31493 8072
rect 31260 8032 31266 8044
rect 31481 8041 31493 8044
rect 31527 8041 31539 8075
rect 31481 8035 31539 8041
rect 31570 8004 31576 8016
rect 31036 7976 31576 8004
rect 31570 7964 31576 7976
rect 31628 7964 31634 8016
rect 31662 7964 31668 8016
rect 31720 8004 31726 8016
rect 32033 8007 32091 8013
rect 32033 8004 32045 8007
rect 31720 7976 32045 8004
rect 31720 7964 31726 7976
rect 32033 7973 32045 7976
rect 32079 7973 32091 8007
rect 32033 7967 32091 7973
rect 21450 7936 21456 7948
rect 21411 7908 21456 7936
rect 21450 7896 21456 7908
rect 21508 7896 21514 7948
rect 21729 7939 21787 7945
rect 21729 7905 21741 7939
rect 21775 7936 21787 7939
rect 22646 7936 22652 7948
rect 21775 7908 22652 7936
rect 21775 7905 21787 7908
rect 21729 7899 21787 7905
rect 22646 7896 22652 7908
rect 22704 7896 22710 7948
rect 30006 7936 30012 7948
rect 23676 7908 30012 7936
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 14090 7868 14096 7880
rect 1903 7840 14096 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 22278 7868 22284 7880
rect 22239 7840 22284 7868
rect 22278 7828 22284 7840
rect 22336 7828 22342 7880
rect 23676 7854 23704 7908
rect 30006 7896 30012 7908
rect 30064 7896 30070 7948
rect 30742 7896 30748 7948
rect 30800 7936 30806 7948
rect 32677 7939 32735 7945
rect 32677 7936 32689 7939
rect 30800 7908 32689 7936
rect 30800 7896 30806 7908
rect 32677 7905 32689 7908
rect 32723 7905 32735 7939
rect 32677 7899 32735 7905
rect 37826 7896 37832 7948
rect 37884 7936 37890 7948
rect 38013 7939 38071 7945
rect 38013 7936 38025 7939
rect 37884 7908 38025 7936
rect 37884 7896 37890 7908
rect 38013 7905 38025 7908
rect 38059 7905 38071 7939
rect 38013 7899 38071 7905
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7868 24823 7871
rect 25682 7868 25688 7880
rect 24811 7840 25688 7868
rect 24811 7837 24823 7840
rect 24765 7831 24823 7837
rect 25682 7828 25688 7840
rect 25740 7828 25746 7880
rect 27246 7828 27252 7880
rect 27304 7868 27310 7880
rect 29270 7868 29276 7880
rect 27304 7840 27752 7868
rect 27304 7828 27310 7840
rect 21358 7760 21364 7812
rect 21416 7800 21422 7812
rect 21637 7803 21695 7809
rect 21637 7800 21649 7803
rect 21416 7772 21649 7800
rect 21416 7760 21422 7772
rect 21637 7769 21649 7772
rect 21683 7769 21695 7803
rect 21637 7763 21695 7769
rect 22557 7803 22615 7809
rect 22557 7769 22569 7803
rect 22603 7769 22615 7803
rect 22557 7763 22615 7769
rect 23860 7772 25636 7800
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 22370 7692 22376 7744
rect 22428 7732 22434 7744
rect 22572 7732 22600 7763
rect 23860 7732 23888 7772
rect 22428 7704 23888 7732
rect 24029 7735 24087 7741
rect 22428 7692 22434 7704
rect 24029 7701 24041 7735
rect 24075 7732 24087 7735
rect 24118 7732 24124 7744
rect 24075 7704 24124 7732
rect 24075 7701 24087 7704
rect 24029 7695 24087 7701
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 25608 7732 25636 7772
rect 26510 7760 26516 7812
rect 26568 7760 26574 7812
rect 26973 7803 27031 7809
rect 26973 7769 26985 7803
rect 27019 7800 27031 7803
rect 27522 7800 27528 7812
rect 27019 7772 27528 7800
rect 27019 7769 27031 7772
rect 26973 7763 27031 7769
rect 27522 7760 27528 7772
rect 27580 7760 27586 7812
rect 27724 7744 27752 7840
rect 28920 7840 29276 7868
rect 26602 7732 26608 7744
rect 25608 7704 26608 7732
rect 26602 7692 26608 7704
rect 26660 7692 26666 7744
rect 27706 7732 27712 7744
rect 27667 7704 27712 7732
rect 27706 7692 27712 7704
rect 27764 7732 27770 7744
rect 28537 7735 28595 7741
rect 28537 7732 28549 7735
rect 27764 7704 28549 7732
rect 27764 7692 27770 7704
rect 28537 7701 28549 7704
rect 28583 7732 28595 7735
rect 28920 7732 28948 7840
rect 29270 7828 29276 7840
rect 29328 7868 29334 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29328 7840 29745 7868
rect 29328 7828 29334 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 32125 7871 32183 7877
rect 32125 7837 32137 7871
rect 32171 7868 32183 7871
rect 32769 7871 32827 7877
rect 32769 7868 32781 7871
rect 32171 7840 32781 7868
rect 32171 7837 32183 7840
rect 32125 7831 32183 7837
rect 32769 7837 32781 7840
rect 32815 7868 32827 7871
rect 33134 7868 33140 7880
rect 32815 7840 33140 7868
rect 32815 7837 32827 7840
rect 32769 7831 32827 7837
rect 33134 7828 33140 7840
rect 33192 7828 33198 7880
rect 38286 7868 38292 7880
rect 38247 7840 38292 7868
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 28994 7760 29000 7812
rect 29052 7800 29058 7812
rect 30009 7803 30067 7809
rect 30009 7800 30021 7803
rect 29052 7772 30021 7800
rect 29052 7760 29058 7772
rect 30009 7769 30021 7772
rect 30055 7769 30067 7803
rect 32030 7800 32036 7812
rect 31234 7772 32036 7800
rect 30009 7763 30067 7769
rect 32030 7760 32036 7772
rect 32088 7760 32094 7812
rect 29089 7735 29147 7741
rect 29089 7732 29101 7735
rect 28583 7704 29101 7732
rect 28583 7701 28595 7704
rect 28537 7695 28595 7701
rect 29089 7701 29101 7704
rect 29135 7701 29147 7735
rect 29089 7695 29147 7701
rect 29546 7692 29552 7744
rect 29604 7732 29610 7744
rect 30190 7732 30196 7744
rect 29604 7704 30196 7732
rect 29604 7692 29610 7704
rect 30190 7692 30196 7704
rect 30248 7692 30254 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 14090 7528 14096 7540
rect 14051 7500 14096 7528
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 21358 7528 21364 7540
rect 21319 7500 21364 7528
rect 21358 7488 21364 7500
rect 21416 7488 21422 7540
rect 22462 7528 22468 7540
rect 22423 7500 22468 7528
rect 22462 7488 22468 7500
rect 22520 7488 22526 7540
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 23477 7531 23535 7537
rect 23477 7528 23489 7531
rect 22796 7500 23489 7528
rect 22796 7488 22802 7500
rect 23477 7497 23489 7500
rect 23523 7497 23535 7531
rect 23477 7491 23535 7497
rect 26142 7488 26148 7540
rect 26200 7528 26206 7540
rect 33045 7531 33103 7537
rect 33045 7528 33057 7531
rect 26200 7500 33057 7528
rect 26200 7488 26206 7500
rect 33045 7497 33057 7500
rect 33091 7497 33103 7531
rect 33686 7528 33692 7540
rect 33647 7500 33692 7528
rect 33045 7491 33103 7497
rect 33686 7488 33692 7500
rect 33744 7488 33750 7540
rect 38286 7528 38292 7540
rect 38247 7500 38292 7528
rect 38286 7488 38292 7500
rect 38344 7488 38350 7540
rect 22370 7460 22376 7472
rect 21468 7432 22376 7460
rect 21468 7401 21496 7432
rect 22370 7420 22376 7432
rect 22428 7420 22434 7472
rect 27246 7460 27252 7472
rect 24518 7432 27252 7460
rect 27246 7420 27252 7432
rect 27304 7420 27310 7472
rect 27430 7420 27436 7472
rect 27488 7460 27494 7472
rect 28994 7460 29000 7472
rect 27488 7432 29000 7460
rect 27488 7420 27494 7432
rect 28994 7420 29000 7432
rect 29052 7420 29058 7472
rect 30650 7460 30656 7472
rect 30611 7432 30656 7460
rect 30650 7420 30656 7432
rect 30708 7420 30714 7472
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7392 14335 7395
rect 21453 7395 21511 7401
rect 14323 7364 14872 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 14844 7197 14872 7364
rect 21453 7361 21465 7395
rect 21499 7361 21511 7395
rect 21453 7355 21511 7361
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7361 22615 7395
rect 31757 7395 31815 7401
rect 30038 7364 30880 7392
rect 22557 7355 22615 7361
rect 22572 7324 22600 7355
rect 23934 7324 23940 7336
rect 22572 7296 23940 7324
rect 23934 7284 23940 7296
rect 23992 7284 23998 7336
rect 24210 7284 24216 7336
rect 24268 7324 24274 7336
rect 24486 7324 24492 7336
rect 24268 7296 24492 7324
rect 24268 7284 24274 7296
rect 24486 7284 24492 7296
rect 24544 7324 24550 7336
rect 24949 7327 25007 7333
rect 24949 7324 24961 7327
rect 24544 7296 24961 7324
rect 24544 7284 24550 7296
rect 24949 7293 24961 7296
rect 24995 7293 25007 7327
rect 24949 7287 25007 7293
rect 25225 7327 25283 7333
rect 25225 7293 25237 7327
rect 25271 7293 25283 7327
rect 25225 7287 25283 7293
rect 25240 7256 25268 7287
rect 25682 7284 25688 7336
rect 25740 7324 25746 7336
rect 27982 7324 27988 7336
rect 25740 7296 27988 7324
rect 25740 7284 25746 7296
rect 27982 7284 27988 7296
rect 28040 7284 28046 7336
rect 28442 7324 28448 7336
rect 28092 7296 28448 7324
rect 27706 7256 27712 7268
rect 25240 7228 25820 7256
rect 25792 7200 25820 7228
rect 26252 7228 27712 7256
rect 14829 7191 14887 7197
rect 14829 7157 14841 7191
rect 14875 7188 14887 7191
rect 25130 7188 25136 7200
rect 14875 7160 25136 7188
rect 14875 7157 14887 7160
rect 14829 7151 14887 7157
rect 25130 7148 25136 7160
rect 25188 7148 25194 7200
rect 25774 7188 25780 7200
rect 25735 7160 25780 7188
rect 25774 7148 25780 7160
rect 25832 7188 25838 7200
rect 26252 7197 26280 7228
rect 27706 7216 27712 7228
rect 27764 7256 27770 7268
rect 28092 7265 28120 7296
rect 28442 7284 28448 7296
rect 28500 7324 28506 7336
rect 28618 7327 28676 7333
rect 28618 7324 28630 7327
rect 28500 7296 28630 7324
rect 28500 7284 28506 7296
rect 28618 7293 28630 7296
rect 28664 7293 28676 7327
rect 28618 7287 28676 7293
rect 28994 7284 29000 7336
rect 29052 7324 29058 7336
rect 30650 7324 30656 7336
rect 29052 7296 30656 7324
rect 29052 7284 29058 7296
rect 30650 7284 30656 7296
rect 30708 7284 30714 7336
rect 30852 7324 30880 7364
rect 31757 7361 31769 7395
rect 31803 7392 31815 7395
rect 32214 7392 32220 7404
rect 31803 7364 32220 7392
rect 31803 7361 31815 7364
rect 31757 7355 31815 7361
rect 32214 7352 32220 7364
rect 32272 7392 32278 7404
rect 32493 7395 32551 7401
rect 32493 7392 32505 7395
rect 32272 7364 32505 7392
rect 32272 7352 32278 7364
rect 32493 7361 32505 7364
rect 32539 7361 32551 7395
rect 33134 7392 33140 7404
rect 33095 7364 33140 7392
rect 32493 7355 32551 7361
rect 33134 7352 33140 7364
rect 33192 7352 33198 7404
rect 34054 7324 34060 7336
rect 30852 7296 34060 7324
rect 34054 7284 34060 7296
rect 34112 7284 34118 7336
rect 28077 7259 28135 7265
rect 28077 7256 28089 7259
rect 27764 7228 28089 7256
rect 27764 7216 27770 7228
rect 28077 7225 28089 7228
rect 28123 7225 28135 7259
rect 32401 7259 32459 7265
rect 32401 7256 32413 7259
rect 28077 7219 28135 7225
rect 30576 7228 32413 7256
rect 26237 7191 26295 7197
rect 26237 7188 26249 7191
rect 25832 7160 26249 7188
rect 25832 7148 25838 7160
rect 26237 7157 26249 7160
rect 26283 7157 26295 7191
rect 26237 7151 26295 7157
rect 27617 7191 27675 7197
rect 27617 7157 27629 7191
rect 27663 7188 27675 7191
rect 27798 7188 27804 7200
rect 27663 7160 27804 7188
rect 27663 7157 27675 7160
rect 27617 7151 27675 7157
rect 27798 7148 27804 7160
rect 27856 7148 27862 7200
rect 28892 7191 28950 7197
rect 28892 7157 28904 7191
rect 28938 7188 28950 7191
rect 29362 7188 29368 7200
rect 28938 7160 29368 7188
rect 28938 7157 28950 7160
rect 28892 7151 28950 7157
rect 29362 7148 29368 7160
rect 29420 7148 29426 7200
rect 29638 7148 29644 7200
rect 29696 7188 29702 7200
rect 30576 7188 30604 7228
rect 32401 7225 32413 7228
rect 32447 7225 32459 7259
rect 32401 7219 32459 7225
rect 29696 7160 30604 7188
rect 29696 7148 29702 7160
rect 30650 7148 30656 7200
rect 30708 7188 30714 7200
rect 31665 7191 31723 7197
rect 31665 7188 31677 7191
rect 30708 7160 31677 7188
rect 30708 7148 30714 7160
rect 31665 7157 31677 7160
rect 31711 7157 31723 7191
rect 31665 7151 31723 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 22544 6987 22602 6993
rect 22544 6953 22556 6987
rect 22590 6984 22602 6987
rect 22738 6984 22744 6996
rect 22590 6956 22744 6984
rect 22590 6953 22602 6956
rect 22544 6947 22602 6953
rect 22738 6944 22744 6956
rect 22796 6944 22802 6996
rect 24844 6987 24902 6993
rect 24844 6953 24856 6987
rect 24890 6984 24902 6987
rect 25590 6984 25596 6996
rect 24890 6956 25596 6984
rect 24890 6953 24902 6956
rect 24844 6947 24902 6953
rect 25590 6944 25596 6956
rect 25648 6944 25654 6996
rect 28463 6987 28521 6993
rect 28463 6953 28475 6987
rect 28509 6984 28521 6987
rect 28810 6984 28816 6996
rect 28509 6956 28816 6984
rect 28509 6953 28521 6956
rect 28463 6947 28521 6953
rect 28810 6944 28816 6956
rect 28868 6944 28874 6996
rect 28902 6944 28908 6996
rect 28960 6984 28966 6996
rect 31662 6984 31668 6996
rect 28960 6956 31668 6984
rect 28960 6944 28966 6956
rect 31662 6944 31668 6956
rect 31720 6944 31726 6996
rect 20625 6851 20683 6857
rect 20625 6817 20637 6851
rect 20671 6848 20683 6851
rect 20714 6848 20720 6860
rect 20671 6820 20720 6848
rect 20671 6817 20683 6820
rect 20625 6811 20683 6817
rect 20714 6808 20720 6820
rect 20772 6848 20778 6860
rect 21450 6848 21456 6860
rect 20772 6820 21456 6848
rect 20772 6808 20778 6820
rect 21450 6808 21456 6820
rect 21508 6808 21514 6860
rect 22278 6848 22284 6860
rect 22191 6820 22284 6848
rect 22278 6808 22284 6820
rect 22336 6848 22342 6860
rect 23290 6848 23296 6860
rect 22336 6820 23296 6848
rect 22336 6808 22342 6820
rect 23290 6808 23296 6820
rect 23348 6808 23354 6860
rect 26142 6848 26148 6860
rect 23676 6820 26148 6848
rect 23676 6766 23704 6820
rect 26142 6808 26148 6820
rect 26200 6808 26206 6860
rect 26329 6851 26387 6857
rect 26329 6817 26341 6851
rect 26375 6848 26387 6851
rect 27154 6848 27160 6860
rect 26375 6820 27160 6848
rect 26375 6817 26387 6820
rect 26329 6811 26387 6817
rect 27154 6808 27160 6820
rect 27212 6808 27218 6860
rect 28442 6808 28448 6860
rect 28500 6848 28506 6860
rect 28721 6851 28779 6857
rect 28721 6848 28733 6851
rect 28500 6820 28733 6848
rect 28500 6808 28506 6820
rect 28721 6817 28733 6820
rect 28767 6848 28779 6851
rect 28767 6820 28994 6848
rect 28767 6817 28779 6820
rect 28721 6811 28779 6817
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 23952 6752 24593 6780
rect 20806 6712 20812 6724
rect 20767 6684 20812 6712
rect 20806 6672 20812 6684
rect 20864 6672 20870 6724
rect 20898 6672 20904 6724
rect 20956 6712 20962 6724
rect 20956 6684 21001 6712
rect 20956 6672 20962 6684
rect 23382 6604 23388 6656
rect 23440 6644 23446 6656
rect 23952 6644 23980 6752
rect 24581 6749 24593 6752
rect 24627 6749 24639 6783
rect 28966 6780 28994 6820
rect 30098 6808 30104 6860
rect 30156 6848 30162 6860
rect 32769 6851 32827 6857
rect 32769 6848 32781 6851
rect 30156 6820 32781 6848
rect 30156 6808 30162 6820
rect 32769 6817 32781 6820
rect 32815 6817 32827 6851
rect 32769 6811 32827 6817
rect 34057 6851 34115 6857
rect 34057 6817 34069 6851
rect 34103 6848 34115 6851
rect 37918 6848 37924 6860
rect 34103 6820 37924 6848
rect 34103 6817 34115 6820
rect 34057 6811 34115 6817
rect 29730 6780 29736 6792
rect 28966 6752 29736 6780
rect 24581 6743 24639 6749
rect 29730 6740 29736 6752
rect 29788 6740 29794 6792
rect 32030 6740 32036 6792
rect 32088 6780 32094 6792
rect 32125 6783 32183 6789
rect 32125 6780 32137 6783
rect 32088 6752 32137 6780
rect 32088 6740 32094 6752
rect 32125 6749 32137 6752
rect 32171 6749 32183 6783
rect 32125 6743 32183 6749
rect 32214 6740 32220 6792
rect 32272 6780 32278 6792
rect 32861 6783 32919 6789
rect 32861 6780 32873 6783
rect 32272 6752 32873 6780
rect 32272 6740 32278 6752
rect 32861 6749 32873 6752
rect 32907 6780 32919 6783
rect 33505 6783 33563 6789
rect 33505 6780 33517 6783
rect 32907 6752 33517 6780
rect 32907 6749 32919 6752
rect 32861 6743 32919 6749
rect 33505 6749 33517 6752
rect 33551 6749 33563 6783
rect 33505 6743 33563 6749
rect 27154 6712 27160 6724
rect 26082 6684 27160 6712
rect 27154 6672 27160 6684
rect 27212 6672 27218 6724
rect 28014 6684 28396 6712
rect 23440 6616 23980 6644
rect 23440 6604 23446 6616
rect 24026 6604 24032 6656
rect 24084 6644 24090 6656
rect 26970 6644 26976 6656
rect 24084 6616 24129 6644
rect 26931 6616 26976 6644
rect 24084 6604 24090 6616
rect 26970 6604 26976 6616
rect 27028 6604 27034 6656
rect 28368 6644 28396 6684
rect 28442 6672 28448 6724
rect 28500 6712 28506 6724
rect 30009 6715 30067 6721
rect 30009 6712 30021 6715
rect 28500 6684 30021 6712
rect 28500 6672 28506 6684
rect 30009 6681 30021 6684
rect 30055 6681 30067 6715
rect 31938 6712 31944 6724
rect 31234 6684 31944 6712
rect 30009 6675 30067 6681
rect 31938 6672 31944 6684
rect 31996 6672 32002 6724
rect 33413 6715 33471 6721
rect 33413 6712 33425 6715
rect 32048 6684 33425 6712
rect 29914 6644 29920 6656
rect 28368 6616 29920 6644
rect 29914 6604 29920 6616
rect 29972 6604 29978 6656
rect 30190 6604 30196 6656
rect 30248 6644 30254 6656
rect 31481 6647 31539 6653
rect 31481 6644 31493 6647
rect 30248 6616 31493 6644
rect 30248 6604 30254 6616
rect 31481 6613 31493 6616
rect 31527 6613 31539 6647
rect 31481 6607 31539 6613
rect 31570 6604 31576 6656
rect 31628 6644 31634 6656
rect 32048 6644 32076 6684
rect 33413 6681 33425 6684
rect 33459 6681 33471 6715
rect 33413 6675 33471 6681
rect 31628 6616 32076 6644
rect 31628 6604 31634 6616
rect 32398 6604 32404 6656
rect 32456 6644 32462 6656
rect 34072 6644 34100 6811
rect 37918 6808 37924 6820
rect 37976 6808 37982 6860
rect 32456 6616 34100 6644
rect 32456 6604 32462 6616
rect 34698 6604 34704 6656
rect 34756 6644 34762 6656
rect 34885 6647 34943 6653
rect 34885 6644 34897 6647
rect 34756 6616 34897 6644
rect 34756 6604 34762 6616
rect 34885 6613 34897 6616
rect 34931 6613 34943 6647
rect 34885 6607 34943 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 20806 6400 20812 6452
rect 20864 6440 20870 6452
rect 21361 6443 21419 6449
rect 21361 6440 21373 6443
rect 20864 6412 21373 6440
rect 20864 6400 20870 6412
rect 21361 6409 21373 6412
rect 21407 6409 21419 6443
rect 24118 6440 24124 6452
rect 21361 6403 21419 6409
rect 21468 6412 24124 6440
rect 21468 6313 21496 6412
rect 24118 6400 24124 6412
rect 24176 6400 24182 6452
rect 27154 6400 27160 6452
rect 27212 6440 27218 6452
rect 31665 6443 31723 6449
rect 31665 6440 31677 6443
rect 27212 6412 31677 6440
rect 27212 6400 27218 6412
rect 31665 6409 31677 6412
rect 31711 6409 31723 6443
rect 31665 6403 31723 6409
rect 31938 6400 31944 6452
rect 31996 6440 32002 6452
rect 32401 6443 32459 6449
rect 32401 6440 32413 6443
rect 31996 6412 32413 6440
rect 31996 6400 32002 6412
rect 32401 6409 32413 6412
rect 32447 6409 32459 6443
rect 32401 6403 32459 6409
rect 22186 6372 22192 6384
rect 22147 6344 22192 6372
rect 22186 6332 22192 6344
rect 22244 6332 22250 6384
rect 24578 6332 24584 6384
rect 24636 6332 24642 6384
rect 25041 6375 25099 6381
rect 25041 6341 25053 6375
rect 25087 6372 25099 6375
rect 26234 6372 26240 6384
rect 25087 6344 26240 6372
rect 25087 6341 25099 6344
rect 25041 6335 25099 6341
rect 26234 6332 26240 6344
rect 26292 6372 26298 6384
rect 27062 6372 27068 6384
rect 26292 6344 27068 6372
rect 26292 6332 26298 6344
rect 27062 6332 27068 6344
rect 27120 6332 27126 6384
rect 27798 6332 27804 6384
rect 27856 6372 27862 6384
rect 27893 6375 27951 6381
rect 27893 6372 27905 6375
rect 27856 6344 27905 6372
rect 27856 6332 27862 6344
rect 27893 6341 27905 6344
rect 27939 6372 27951 6375
rect 28350 6372 28356 6384
rect 27939 6344 28356 6372
rect 27939 6341 27951 6344
rect 27893 6335 27951 6341
rect 28350 6332 28356 6344
rect 28408 6332 28414 6384
rect 29638 6372 29644 6384
rect 29210 6344 29644 6372
rect 29638 6332 29644 6344
rect 29696 6332 29702 6384
rect 29730 6332 29736 6384
rect 29788 6372 29794 6384
rect 30377 6375 30435 6381
rect 30377 6372 30389 6375
rect 29788 6344 30389 6372
rect 29788 6332 29794 6344
rect 29932 6313 29960 6344
rect 30377 6341 30389 6344
rect 30423 6341 30435 6375
rect 30377 6335 30435 6341
rect 30466 6332 30472 6384
rect 30524 6372 30530 6384
rect 33045 6375 33103 6381
rect 33045 6372 33057 6375
rect 30524 6344 33057 6372
rect 30524 6332 30530 6344
rect 33045 6341 33057 6344
rect 33091 6341 33103 6375
rect 33045 6335 33103 6341
rect 33152 6344 34468 6372
rect 33152 6316 33180 6344
rect 21453 6307 21511 6313
rect 21453 6273 21465 6307
rect 21499 6273 21511 6307
rect 21453 6267 21511 6273
rect 29917 6307 29975 6313
rect 29917 6273 29929 6307
rect 29963 6273 29975 6307
rect 29917 6267 29975 6273
rect 31113 6307 31171 6313
rect 31113 6273 31125 6307
rect 31159 6304 31171 6307
rect 31757 6307 31815 6313
rect 31757 6304 31769 6307
rect 31159 6276 31769 6304
rect 31159 6273 31171 6276
rect 31113 6267 31171 6273
rect 31757 6273 31769 6276
rect 31803 6304 31815 6307
rect 32214 6304 32220 6316
rect 31803 6276 32220 6304
rect 31803 6273 31815 6276
rect 31757 6267 31815 6273
rect 32214 6264 32220 6276
rect 32272 6304 32278 6316
rect 32493 6307 32551 6313
rect 32493 6304 32505 6307
rect 32272 6276 32505 6304
rect 32272 6264 32278 6276
rect 32493 6273 32505 6276
rect 32539 6273 32551 6307
rect 33134 6304 33140 6316
rect 33095 6276 33140 6304
rect 32493 6267 32551 6273
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 25317 6239 25375 6245
rect 22152 6208 22197 6236
rect 22152 6196 22158 6208
rect 25317 6205 25329 6239
rect 25363 6236 25375 6239
rect 29641 6239 29699 6245
rect 25363 6208 25820 6236
rect 25363 6205 25375 6208
rect 25317 6199 25375 6205
rect 22646 6168 22652 6180
rect 22607 6140 22652 6168
rect 22646 6128 22652 6140
rect 22704 6128 22710 6180
rect 25792 6112 25820 6208
rect 29641 6205 29653 6239
rect 29687 6236 29699 6239
rect 32398 6236 32404 6248
rect 29687 6208 32404 6236
rect 29687 6205 29699 6208
rect 29641 6199 29699 6205
rect 32398 6196 32404 6208
rect 32456 6196 32462 6248
rect 32508 6236 32536 6267
rect 33134 6264 33140 6276
rect 33192 6264 33198 6316
rect 34440 6313 34468 6344
rect 33597 6307 33655 6313
rect 33597 6273 33609 6307
rect 33643 6273 33655 6307
rect 33597 6267 33655 6273
rect 34425 6307 34483 6313
rect 34425 6273 34437 6307
rect 34471 6273 34483 6307
rect 34425 6267 34483 6273
rect 33612 6236 33640 6267
rect 32508 6208 33640 6236
rect 29914 6128 29920 6180
rect 29972 6168 29978 6180
rect 34333 6171 34391 6177
rect 34333 6168 34345 6171
rect 29972 6140 34345 6168
rect 29972 6128 29978 6140
rect 34333 6137 34345 6140
rect 34379 6137 34391 6171
rect 34333 6131 34391 6137
rect 23566 6100 23572 6112
rect 23527 6072 23572 6100
rect 23566 6060 23572 6072
rect 23624 6100 23630 6112
rect 24486 6100 24492 6112
rect 23624 6072 24492 6100
rect 23624 6060 23630 6072
rect 24486 6060 24492 6072
rect 24544 6060 24550 6112
rect 25774 6100 25780 6112
rect 25735 6072 25780 6100
rect 25774 6060 25780 6072
rect 25832 6100 25838 6112
rect 26329 6103 26387 6109
rect 26329 6100 26341 6103
rect 25832 6072 26341 6100
rect 25832 6060 25838 6072
rect 26329 6069 26341 6072
rect 26375 6100 26387 6103
rect 27157 6103 27215 6109
rect 27157 6100 27169 6103
rect 26375 6072 27169 6100
rect 26375 6069 26387 6072
rect 26329 6063 26387 6069
rect 27157 6069 27169 6072
rect 27203 6069 27215 6103
rect 27157 6063 27215 6069
rect 27982 6060 27988 6112
rect 28040 6100 28046 6112
rect 30834 6100 30840 6112
rect 28040 6072 30840 6100
rect 28040 6060 28046 6072
rect 30834 6060 30840 6072
rect 30892 6060 30898 6112
rect 31018 6100 31024 6112
rect 30979 6072 31024 6100
rect 31018 6060 31024 6072
rect 31076 6060 31082 6112
rect 31110 6060 31116 6112
rect 31168 6100 31174 6112
rect 31662 6100 31668 6112
rect 31168 6072 31668 6100
rect 31168 6060 31174 6072
rect 31662 6060 31668 6072
rect 31720 6060 31726 6112
rect 32030 6060 32036 6112
rect 32088 6100 32094 6112
rect 33689 6103 33747 6109
rect 33689 6100 33701 6103
rect 32088 6072 33701 6100
rect 32088 6060 32094 6072
rect 33689 6069 33701 6072
rect 33735 6069 33747 6103
rect 33689 6063 33747 6069
rect 34790 6060 34796 6112
rect 34848 6100 34854 6112
rect 34885 6103 34943 6109
rect 34885 6100 34897 6103
rect 34848 6072 34897 6100
rect 34848 6060 34854 6072
rect 34885 6069 34897 6072
rect 34931 6069 34943 6103
rect 35526 6100 35532 6112
rect 35487 6072 35532 6100
rect 34885 6063 34943 6069
rect 35526 6060 35532 6072
rect 35584 6060 35590 6112
rect 36078 6100 36084 6112
rect 36039 6072 36084 6100
rect 36078 6060 36084 6072
rect 36136 6060 36142 6112
rect 37458 6060 37464 6112
rect 37516 6100 37522 6112
rect 37645 6103 37703 6109
rect 37645 6100 37657 6103
rect 37516 6072 37657 6100
rect 37516 6060 37522 6072
rect 37645 6069 37657 6072
rect 37691 6069 37703 6103
rect 38194 6100 38200 6112
rect 38155 6072 38200 6100
rect 37645 6063 37703 6069
rect 38194 6060 38200 6072
rect 38252 6060 38258 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 24578 5856 24584 5908
rect 24636 5896 24642 5908
rect 33873 5899 33931 5905
rect 33873 5896 33885 5899
rect 24636 5868 33885 5896
rect 24636 5856 24642 5868
rect 33873 5865 33885 5868
rect 33919 5865 33931 5899
rect 33873 5859 33931 5865
rect 36170 5856 36176 5908
rect 36228 5896 36234 5908
rect 38105 5899 38163 5905
rect 38105 5896 38117 5899
rect 36228 5868 38117 5896
rect 36228 5856 36234 5868
rect 38105 5865 38117 5868
rect 38151 5865 38163 5899
rect 38105 5859 38163 5865
rect 26602 5788 26608 5840
rect 26660 5828 26666 5840
rect 26973 5831 27031 5837
rect 26973 5828 26985 5831
rect 26660 5800 26985 5828
rect 26660 5788 26666 5800
rect 26973 5797 26985 5800
rect 27019 5797 27031 5831
rect 29178 5828 29184 5840
rect 29139 5800 29184 5828
rect 26973 5791 27031 5797
rect 29178 5788 29184 5800
rect 29236 5788 29242 5840
rect 33686 5828 33692 5840
rect 32876 5800 33692 5828
rect 24026 5720 24032 5772
rect 24084 5760 24090 5772
rect 25501 5763 25559 5769
rect 25501 5760 25513 5763
rect 24084 5732 25513 5760
rect 24084 5720 24090 5732
rect 25501 5729 25513 5732
rect 25547 5729 25559 5763
rect 25501 5723 25559 5729
rect 27246 5720 27252 5772
rect 27304 5760 27310 5772
rect 27709 5763 27767 5769
rect 27709 5760 27721 5763
rect 27304 5732 27721 5760
rect 27304 5720 27310 5732
rect 27709 5729 27721 5732
rect 27755 5729 27767 5763
rect 27709 5723 27767 5729
rect 28828 5732 31616 5760
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 4985 5695 5043 5701
rect 4985 5692 4997 5695
rect 1903 5664 4997 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 4985 5661 4997 5664
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5692 5135 5695
rect 25225 5695 25283 5701
rect 25225 5692 25237 5695
rect 5123 5664 5672 5692
rect 5123 5661 5135 5664
rect 5077 5655 5135 5661
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 5644 5565 5672 5664
rect 24596 5664 25237 5692
rect 24596 5568 24624 5664
rect 25225 5661 25237 5664
rect 25271 5661 25283 5695
rect 27430 5692 27436 5704
rect 27391 5664 27436 5692
rect 25225 5655 25283 5661
rect 27430 5652 27436 5664
rect 27488 5652 27494 5704
rect 28828 5678 28856 5732
rect 31481 5695 31539 5701
rect 31481 5661 31493 5695
rect 31527 5661 31539 5695
rect 31481 5655 31539 5661
rect 31110 5624 31116 5636
rect 26726 5596 27384 5624
rect 30774 5596 31116 5624
rect 5629 5559 5687 5565
rect 5629 5525 5641 5559
rect 5675 5556 5687 5559
rect 20714 5556 20720 5568
rect 5675 5528 20720 5556
rect 5675 5525 5687 5528
rect 5629 5519 5687 5525
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 21821 5559 21879 5565
rect 21821 5525 21833 5559
rect 21867 5556 21879 5559
rect 22186 5556 22192 5568
rect 21867 5528 22192 5556
rect 21867 5525 21879 5528
rect 21821 5519 21879 5525
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 22278 5516 22284 5568
rect 22336 5556 22342 5568
rect 24578 5556 24584 5568
rect 22336 5528 22381 5556
rect 24539 5528 24584 5556
rect 22336 5516 22342 5528
rect 24578 5516 24584 5528
rect 24636 5516 24642 5568
rect 27356 5556 27384 5596
rect 31110 5584 31116 5596
rect 31168 5584 31174 5636
rect 31202 5584 31208 5636
rect 31260 5624 31266 5636
rect 31496 5624 31524 5655
rect 31260 5596 31305 5624
rect 31404 5596 31524 5624
rect 31260 5584 31266 5596
rect 31404 5568 31432 5596
rect 28718 5556 28724 5568
rect 27356 5528 28724 5556
rect 28718 5516 28724 5528
rect 28776 5516 28782 5568
rect 29086 5516 29092 5568
rect 29144 5556 29150 5568
rect 29733 5559 29791 5565
rect 29733 5556 29745 5559
rect 29144 5528 29745 5556
rect 29144 5516 29150 5528
rect 29733 5525 29745 5528
rect 29779 5525 29791 5559
rect 29733 5519 29791 5525
rect 31386 5516 31392 5568
rect 31444 5516 31450 5568
rect 31588 5556 31616 5732
rect 31662 5720 31668 5772
rect 31720 5760 31726 5772
rect 32306 5760 32312 5772
rect 31720 5732 32312 5760
rect 31720 5720 31726 5732
rect 32306 5720 32312 5732
rect 32364 5720 32370 5772
rect 32876 5704 32904 5800
rect 33686 5788 33692 5800
rect 33744 5788 33750 5840
rect 34977 5763 35035 5769
rect 34977 5760 34989 5763
rect 32968 5732 34989 5760
rect 32125 5695 32183 5701
rect 32125 5661 32137 5695
rect 32171 5692 32183 5695
rect 32214 5692 32220 5704
rect 32171 5664 32220 5692
rect 32171 5661 32183 5664
rect 32125 5655 32183 5661
rect 32214 5652 32220 5664
rect 32272 5652 32278 5704
rect 32858 5692 32864 5704
rect 32771 5664 32864 5692
rect 32858 5652 32864 5664
rect 32916 5652 32922 5704
rect 31662 5584 31668 5636
rect 31720 5624 31726 5636
rect 32968 5624 32996 5732
rect 34977 5729 34989 5732
rect 35023 5729 35035 5763
rect 34977 5723 35035 5729
rect 33226 5652 33232 5704
rect 33284 5692 33290 5704
rect 33965 5695 34023 5701
rect 33965 5692 33977 5695
rect 33284 5664 33977 5692
rect 33284 5652 33290 5664
rect 33965 5661 33977 5664
rect 34011 5692 34023 5695
rect 34422 5692 34428 5704
rect 34011 5664 34428 5692
rect 34011 5661 34023 5664
rect 33965 5655 34023 5661
rect 34422 5652 34428 5664
rect 34480 5692 34486 5704
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 34480 5664 34897 5692
rect 34480 5652 34486 5664
rect 34885 5661 34897 5664
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 37645 5695 37703 5701
rect 37645 5661 37657 5695
rect 37691 5692 37703 5695
rect 38286 5692 38292 5704
rect 37691 5664 38292 5692
rect 37691 5661 37703 5664
rect 37645 5655 37703 5661
rect 38286 5652 38292 5664
rect 38344 5652 38350 5704
rect 31720 5596 32996 5624
rect 33137 5627 33195 5633
rect 31720 5584 31726 5596
rect 33137 5593 33149 5627
rect 33183 5593 33195 5627
rect 33137 5587 33195 5593
rect 32033 5559 32091 5565
rect 32033 5556 32045 5559
rect 31588 5528 32045 5556
rect 32033 5525 32045 5528
rect 32079 5525 32091 5559
rect 32033 5519 32091 5525
rect 32214 5516 32220 5568
rect 32272 5556 32278 5568
rect 33152 5556 33180 5587
rect 34790 5584 34796 5636
rect 34848 5624 34854 5636
rect 36633 5627 36691 5633
rect 36633 5624 36645 5627
rect 34848 5596 36645 5624
rect 34848 5584 34854 5596
rect 36633 5593 36645 5596
rect 36679 5593 36691 5627
rect 36633 5587 36691 5593
rect 35526 5556 35532 5568
rect 32272 5528 33180 5556
rect 35487 5528 35532 5556
rect 32272 5516 32278 5528
rect 35526 5516 35532 5528
rect 35584 5556 35590 5568
rect 36081 5559 36139 5565
rect 36081 5556 36093 5559
rect 35584 5528 36093 5556
rect 35584 5516 35590 5528
rect 36081 5525 36093 5528
rect 36127 5525 36139 5559
rect 36081 5519 36139 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22152 5324 22197 5352
rect 22152 5312 22158 5324
rect 24578 5312 24584 5364
rect 24636 5352 24642 5364
rect 25685 5355 25743 5361
rect 25685 5352 25697 5355
rect 24636 5324 25697 5352
rect 24636 5312 24642 5324
rect 25685 5321 25697 5324
rect 25731 5352 25743 5355
rect 25774 5352 25780 5364
rect 25731 5324 25780 5352
rect 25731 5321 25743 5324
rect 25685 5315 25743 5321
rect 25774 5312 25780 5324
rect 25832 5352 25838 5364
rect 26513 5355 26571 5361
rect 26513 5352 26525 5355
rect 25832 5324 26525 5352
rect 25832 5312 25838 5324
rect 26513 5321 26525 5324
rect 26559 5352 26571 5355
rect 26694 5352 26700 5364
rect 26559 5324 26700 5352
rect 26559 5321 26571 5324
rect 26513 5315 26571 5321
rect 26694 5312 26700 5324
rect 26752 5352 26758 5364
rect 27157 5355 27215 5361
rect 27157 5352 27169 5355
rect 26752 5324 27169 5352
rect 26752 5312 26758 5324
rect 27157 5321 27169 5324
rect 27203 5352 27215 5355
rect 27430 5352 27436 5364
rect 27203 5324 27436 5352
rect 27203 5321 27215 5324
rect 27157 5315 27215 5321
rect 27430 5312 27436 5324
rect 27488 5352 27494 5364
rect 27709 5355 27767 5361
rect 27709 5352 27721 5355
rect 27488 5324 27721 5352
rect 27488 5312 27494 5324
rect 27709 5321 27721 5324
rect 27755 5352 27767 5355
rect 28350 5352 28356 5364
rect 27755 5324 28356 5352
rect 27755 5321 27767 5324
rect 27709 5315 27767 5321
rect 28350 5312 28356 5324
rect 28408 5312 28414 5364
rect 29454 5312 29460 5364
rect 29512 5352 29518 5364
rect 29914 5352 29920 5364
rect 29512 5324 29920 5352
rect 29512 5312 29518 5324
rect 29914 5312 29920 5324
rect 29972 5352 29978 5364
rect 30101 5355 30159 5361
rect 30101 5352 30113 5355
rect 29972 5324 30113 5352
rect 29972 5312 29978 5324
rect 30101 5321 30113 5324
rect 30147 5321 30159 5355
rect 30101 5315 30159 5321
rect 23566 5284 23572 5296
rect 21192 5256 23572 5284
rect 21192 5225 21220 5256
rect 23566 5244 23572 5256
rect 23624 5244 23630 5296
rect 27522 5244 27528 5296
rect 27580 5284 27586 5296
rect 28629 5287 28687 5293
rect 28629 5284 28641 5287
rect 27580 5256 28641 5284
rect 27580 5244 27586 5256
rect 28629 5253 28641 5256
rect 28675 5284 28687 5287
rect 28902 5284 28908 5296
rect 28675 5256 28908 5284
rect 28675 5253 28687 5256
rect 28629 5247 28687 5253
rect 28902 5244 28908 5256
rect 28960 5244 28966 5296
rect 31018 5284 31024 5296
rect 29854 5256 31024 5284
rect 31018 5244 31024 5256
rect 31076 5244 31082 5296
rect 33134 5284 33140 5296
rect 32784 5256 33140 5284
rect 20349 5219 20407 5225
rect 20349 5185 20361 5219
rect 20395 5216 20407 5219
rect 21085 5219 21143 5225
rect 21085 5216 21097 5219
rect 20395 5188 21097 5216
rect 20395 5185 20407 5188
rect 20349 5179 20407 5185
rect 21085 5185 21097 5188
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5185 21235 5219
rect 21177 5179 21235 5185
rect 21266 5176 21272 5228
rect 21324 5216 21330 5228
rect 22189 5219 22247 5225
rect 22189 5216 22201 5219
rect 21324 5188 22201 5216
rect 21324 5176 21330 5188
rect 22189 5185 22201 5188
rect 22235 5216 22247 5219
rect 22278 5216 22284 5228
rect 22235 5188 22284 5216
rect 22235 5185 22247 5188
rect 22189 5179 22247 5185
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 22738 5176 22744 5228
rect 22796 5216 22802 5228
rect 22833 5219 22891 5225
rect 22833 5216 22845 5219
rect 22796 5188 22845 5216
rect 22796 5176 22802 5188
rect 22833 5185 22845 5188
rect 22879 5185 22891 5219
rect 28350 5216 28356 5228
rect 24794 5188 27660 5216
rect 28311 5188 28356 5216
rect 22833 5179 22891 5185
rect 20530 5148 20536 5160
rect 20491 5120 20536 5148
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 23382 5148 23388 5160
rect 23343 5120 23388 5148
rect 23382 5108 23388 5120
rect 23440 5108 23446 5160
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 25133 5151 25191 5157
rect 23707 5120 25084 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 20165 5083 20223 5089
rect 20165 5049 20177 5083
rect 20211 5080 20223 5083
rect 20438 5080 20444 5092
rect 20211 5052 20444 5080
rect 20211 5049 20223 5052
rect 20165 5043 20223 5049
rect 20438 5040 20444 5052
rect 20496 5080 20502 5092
rect 20898 5080 20904 5092
rect 20496 5052 20904 5080
rect 20496 5040 20502 5052
rect 20898 5040 20904 5052
rect 20956 5040 20962 5092
rect 25056 5080 25084 5120
rect 25133 5117 25145 5151
rect 25179 5148 25191 5151
rect 25590 5148 25596 5160
rect 25179 5120 25596 5148
rect 25179 5117 25191 5120
rect 25133 5111 25191 5117
rect 25590 5108 25596 5120
rect 25648 5108 25654 5160
rect 27632 5148 27660 5188
rect 28350 5176 28356 5188
rect 28408 5176 28414 5228
rect 31113 5219 31171 5225
rect 31113 5185 31125 5219
rect 31159 5185 31171 5219
rect 31113 5179 31171 5185
rect 31757 5219 31815 5225
rect 31757 5185 31769 5219
rect 31803 5216 31815 5219
rect 32784 5216 32812 5256
rect 33134 5244 33140 5256
rect 33192 5244 33198 5296
rect 35345 5287 35403 5293
rect 35345 5284 35357 5287
rect 34256 5256 35357 5284
rect 31803 5188 32812 5216
rect 31803 5185 31815 5188
rect 31757 5179 31815 5185
rect 29086 5148 29092 5160
rect 27632 5120 29092 5148
rect 29086 5108 29092 5120
rect 29144 5108 29150 5160
rect 29270 5108 29276 5160
rect 29328 5148 29334 5160
rect 31021 5151 31079 5157
rect 31021 5148 31033 5151
rect 29328 5120 31033 5148
rect 29328 5108 29334 5120
rect 31021 5117 31033 5120
rect 31067 5117 31079 5151
rect 31128 5148 31156 5179
rect 32858 5176 32864 5228
rect 32916 5216 32922 5228
rect 34256 5225 34284 5256
rect 35345 5253 35357 5256
rect 35391 5284 35403 5287
rect 35526 5284 35532 5296
rect 35391 5256 35532 5284
rect 35391 5253 35403 5256
rect 35345 5247 35403 5253
rect 35526 5244 35532 5256
rect 35584 5284 35590 5296
rect 35897 5287 35955 5293
rect 35897 5284 35909 5287
rect 35584 5256 35909 5284
rect 35584 5244 35590 5256
rect 35897 5253 35909 5256
rect 35943 5284 35955 5287
rect 36446 5284 36452 5296
rect 35943 5256 36452 5284
rect 35943 5253 35955 5256
rect 35897 5247 35955 5253
rect 36446 5244 36452 5256
rect 36504 5244 36510 5296
rect 34241 5219 34299 5225
rect 34241 5216 34253 5219
rect 32916 5188 34253 5216
rect 32916 5176 32922 5188
rect 34241 5185 34253 5188
rect 34287 5185 34299 5219
rect 34241 5179 34299 5185
rect 34422 5176 34428 5228
rect 34480 5216 34486 5228
rect 34885 5219 34943 5225
rect 34885 5216 34897 5219
rect 34480 5188 34897 5216
rect 34480 5176 34486 5188
rect 34885 5185 34897 5188
rect 34931 5185 34943 5219
rect 34885 5179 34943 5185
rect 32876 5148 32904 5176
rect 31128 5120 32904 5148
rect 31021 5111 31079 5117
rect 33778 5108 33784 5160
rect 33836 5148 33842 5160
rect 33965 5151 34023 5157
rect 33965 5148 33977 5151
rect 33836 5120 33977 5148
rect 33836 5108 33842 5120
rect 33965 5117 33977 5120
rect 34011 5117 34023 5151
rect 33965 5111 34023 5117
rect 26970 5080 26976 5092
rect 25056 5052 26976 5080
rect 26970 5040 26976 5052
rect 27028 5040 27034 5092
rect 31386 5040 31392 5092
rect 31444 5080 31450 5092
rect 31444 5052 31984 5080
rect 31444 5040 31450 5052
rect 31956 5024 31984 5052
rect 22094 4972 22100 5024
rect 22152 5012 22158 5024
rect 22741 5015 22799 5021
rect 22741 5012 22753 5015
rect 22152 4984 22753 5012
rect 22152 4972 22158 4984
rect 22741 4981 22753 4984
rect 22787 4981 22799 5015
rect 22741 4975 22799 4981
rect 28994 4972 29000 5024
rect 29052 5012 29058 5024
rect 31665 5015 31723 5021
rect 31665 5012 31677 5015
rect 29052 4984 31677 5012
rect 29052 4972 29058 4984
rect 31665 4981 31677 4984
rect 31711 4981 31723 5015
rect 31665 4975 31723 4981
rect 31938 4972 31944 5024
rect 31996 5012 32002 5024
rect 32309 5015 32367 5021
rect 32309 5012 32321 5015
rect 31996 4984 32321 5012
rect 31996 4972 32002 4984
rect 32309 4981 32321 4984
rect 32355 4981 32367 5015
rect 32309 4975 32367 4981
rect 34514 4972 34520 5024
rect 34572 5012 34578 5024
rect 34793 5015 34851 5021
rect 34793 5012 34805 5015
rect 34572 4984 34805 5012
rect 34572 4972 34578 4984
rect 34793 4981 34805 4984
rect 34839 4981 34851 5015
rect 34793 4975 34851 4981
rect 36538 4972 36544 5024
rect 36596 5012 36602 5024
rect 37461 5015 37519 5021
rect 37461 5012 37473 5015
rect 36596 4984 37473 5012
rect 36596 4972 36602 4984
rect 37461 4981 37473 4984
rect 37507 4981 37519 5015
rect 38286 5012 38292 5024
rect 38247 4984 38292 5012
rect 37461 4975 37519 4981
rect 38286 4972 38292 4984
rect 38344 4972 38350 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 20898 4768 20904 4820
rect 20956 4808 20962 4820
rect 21637 4811 21695 4817
rect 21637 4808 21649 4811
rect 20956 4780 21649 4808
rect 20956 4768 20962 4780
rect 21637 4777 21649 4780
rect 21683 4777 21695 4811
rect 21637 4771 21695 4777
rect 24029 4811 24087 4817
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 24394 4808 24400 4820
rect 24075 4780 24400 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 24394 4768 24400 4780
rect 24452 4768 24458 4820
rect 26329 4811 26387 4817
rect 26329 4777 26341 4811
rect 26375 4808 26387 4811
rect 26786 4808 26792 4820
rect 26375 4780 26792 4808
rect 26375 4777 26387 4780
rect 26329 4771 26387 4777
rect 26786 4768 26792 4780
rect 26844 4768 26850 4820
rect 26896 4780 28120 4808
rect 24412 4740 24440 4768
rect 24412 4712 24716 4740
rect 22094 4632 22100 4684
rect 22152 4672 22158 4684
rect 24688 4672 24716 4712
rect 26050 4700 26056 4752
rect 26108 4740 26114 4752
rect 26896 4740 26924 4780
rect 26108 4712 26924 4740
rect 28092 4740 28120 4780
rect 28350 4768 28356 4820
rect 28408 4808 28414 4820
rect 28997 4811 29055 4817
rect 28997 4808 29009 4811
rect 28408 4780 29009 4808
rect 28408 4768 28414 4780
rect 28997 4777 29009 4780
rect 29043 4777 29055 4811
rect 28997 4771 29055 4777
rect 28534 4740 28540 4752
rect 28092 4712 28540 4740
rect 26108 4700 26114 4712
rect 28534 4700 28540 4712
rect 28592 4700 28598 4752
rect 24857 4675 24915 4681
rect 24857 4672 24869 4675
rect 22152 4644 22197 4672
rect 24688 4644 24869 4672
rect 22152 4632 22158 4644
rect 24857 4641 24869 4644
rect 24903 4672 24915 4675
rect 25406 4672 25412 4684
rect 24903 4644 25412 4672
rect 24903 4641 24915 4644
rect 24857 4635 24915 4641
rect 25406 4632 25412 4644
rect 25464 4632 25470 4684
rect 25866 4632 25872 4684
rect 25924 4672 25930 4684
rect 26142 4672 26148 4684
rect 25924 4644 26148 4672
rect 25924 4632 25930 4644
rect 26142 4632 26148 4644
rect 26200 4672 26206 4684
rect 27065 4675 27123 4681
rect 27065 4672 27077 4675
rect 26200 4644 27077 4672
rect 26200 4632 26206 4644
rect 27065 4641 27077 4644
rect 27111 4641 27123 4675
rect 29012 4672 29040 4771
rect 29086 4768 29092 4820
rect 29144 4808 29150 4820
rect 30742 4808 30748 4820
rect 29144 4780 30748 4808
rect 29144 4768 29150 4780
rect 30742 4768 30748 4780
rect 30800 4768 30806 4820
rect 31018 4768 31024 4820
rect 31076 4808 31082 4820
rect 31481 4811 31539 4817
rect 31481 4808 31493 4811
rect 31076 4780 31493 4808
rect 31076 4768 31082 4780
rect 31481 4777 31493 4780
rect 31527 4777 31539 4811
rect 32122 4808 32128 4820
rect 32083 4780 32128 4808
rect 31481 4771 31539 4777
rect 32122 4768 32128 4780
rect 32180 4768 32186 4820
rect 34054 4808 34060 4820
rect 34015 4780 34060 4808
rect 34054 4768 34060 4780
rect 34112 4768 34118 4820
rect 36446 4768 36452 4820
rect 36504 4808 36510 4820
rect 36541 4811 36599 4817
rect 36541 4808 36553 4811
rect 36504 4780 36553 4808
rect 36504 4768 36510 4780
rect 36541 4777 36553 4780
rect 36587 4777 36599 4811
rect 36541 4771 36599 4777
rect 31110 4700 31116 4752
rect 31168 4740 31174 4752
rect 32769 4743 32827 4749
rect 32769 4740 32781 4743
rect 31168 4712 32781 4740
rect 31168 4700 31174 4712
rect 32769 4709 32781 4712
rect 32815 4709 32827 4743
rect 32769 4703 32827 4709
rect 29733 4675 29791 4681
rect 29733 4672 29745 4675
rect 29012 4644 29745 4672
rect 27065 4635 27123 4641
rect 29733 4641 29745 4644
rect 29779 4672 29791 4675
rect 30098 4672 30104 4684
rect 29779 4644 30104 4672
rect 29779 4641 29791 4644
rect 29733 4635 29791 4641
rect 30098 4632 30104 4644
rect 30156 4632 30162 4684
rect 31294 4632 31300 4684
rect 31352 4672 31358 4684
rect 37093 4675 37151 4681
rect 37093 4672 37105 4675
rect 31352 4644 37105 4672
rect 31352 4632 31358 4644
rect 37093 4641 37105 4644
rect 37139 4641 37151 4675
rect 37093 4635 37151 4641
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 22244 4576 22293 4604
rect 22244 4564 22250 4576
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 24578 4604 24584 4616
rect 24539 4576 24584 4604
rect 22281 4567 22339 4573
rect 24578 4564 24584 4576
rect 24636 4564 24642 4616
rect 26694 4564 26700 4616
rect 26752 4604 26758 4616
rect 26789 4607 26847 4613
rect 26789 4604 26801 4607
rect 26752 4576 26801 4604
rect 26752 4564 26758 4576
rect 26789 4573 26801 4576
rect 26835 4573 26847 4607
rect 29270 4604 29276 4616
rect 28198 4576 29276 4604
rect 26789 4567 26847 4573
rect 29270 4564 29276 4576
rect 29328 4564 29334 4616
rect 32217 4607 32275 4613
rect 32217 4573 32229 4607
rect 32263 4573 32275 4607
rect 32858 4604 32864 4616
rect 32819 4576 32864 4604
rect 32217 4567 32275 4573
rect 26082 4508 27016 4536
rect 20622 4468 20628 4480
rect 20583 4440 20628 4468
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 22925 4471 22983 4477
rect 22925 4437 22937 4471
rect 22971 4468 22983 4471
rect 23382 4468 23388 4480
rect 22971 4440 23388 4468
rect 22971 4437 22983 4440
rect 22925 4431 22983 4437
rect 23382 4428 23388 4440
rect 23440 4428 23446 4480
rect 26988 4468 27016 4508
rect 28368 4508 28672 4536
rect 28368 4468 28396 4508
rect 26988 4440 28396 4468
rect 28644 4468 28672 4508
rect 29178 4496 29184 4548
rect 29236 4536 29242 4548
rect 30009 4539 30067 4545
rect 30009 4536 30021 4539
rect 29236 4508 30021 4536
rect 29236 4496 29242 4508
rect 30009 4505 30021 4508
rect 30055 4505 30067 4539
rect 32030 4536 32036 4548
rect 31234 4508 32036 4536
rect 30009 4499 30067 4505
rect 32030 4496 32036 4508
rect 32088 4496 32094 4548
rect 32232 4536 32260 4567
rect 32858 4564 32864 4576
rect 32916 4604 32922 4616
rect 33505 4607 33563 4613
rect 33505 4604 33517 4607
rect 32916 4576 33517 4604
rect 32916 4564 32922 4576
rect 33505 4573 33517 4576
rect 33551 4573 33563 4607
rect 33505 4567 33563 4573
rect 33778 4564 33784 4616
rect 33836 4604 33842 4616
rect 34149 4607 34207 4613
rect 34149 4604 34161 4607
rect 33836 4576 34161 4604
rect 33836 4564 33842 4576
rect 34149 4573 34161 4576
rect 34195 4573 34207 4607
rect 37826 4604 37832 4616
rect 37787 4576 37832 4604
rect 34149 4567 34207 4573
rect 37826 4564 37832 4576
rect 37884 4564 37890 4616
rect 33134 4536 33140 4548
rect 32232 4508 33140 4536
rect 33134 4496 33140 4508
rect 33192 4496 33198 4548
rect 34606 4536 34612 4548
rect 33244 4508 34612 4536
rect 33244 4468 33272 4508
rect 34606 4496 34612 4508
rect 34664 4496 34670 4548
rect 33410 4468 33416 4480
rect 28644 4440 33272 4468
rect 33371 4440 33416 4468
rect 33410 4428 33416 4440
rect 33468 4428 33474 4480
rect 34882 4468 34888 4480
rect 34843 4440 34888 4468
rect 34882 4428 34888 4440
rect 34940 4468 34946 4480
rect 35437 4471 35495 4477
rect 35437 4468 35449 4471
rect 34940 4440 35449 4468
rect 34940 4428 34946 4440
rect 35437 4437 35449 4440
rect 35483 4437 35495 4471
rect 35986 4468 35992 4480
rect 35947 4440 35992 4468
rect 35437 4431 35495 4437
rect 35986 4428 35992 4440
rect 36044 4428 36050 4480
rect 38010 4468 38016 4480
rect 37971 4440 38016 4468
rect 38010 4428 38016 4440
rect 38068 4428 38074 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 20349 4267 20407 4273
rect 20349 4233 20361 4267
rect 20395 4264 20407 4267
rect 20530 4264 20536 4276
rect 20395 4236 20536 4264
rect 20395 4233 20407 4236
rect 20349 4227 20407 4233
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 24578 4224 24584 4276
rect 24636 4264 24642 4276
rect 25869 4267 25927 4273
rect 25869 4264 25881 4267
rect 24636 4236 25881 4264
rect 24636 4224 24642 4236
rect 25869 4233 25881 4236
rect 25915 4233 25927 4267
rect 34422 4264 34428 4276
rect 25869 4227 25927 4233
rect 28276 4236 34428 4264
rect 28276 4196 28304 4236
rect 34422 4224 34428 4236
rect 34480 4224 34486 4276
rect 35526 4224 35532 4276
rect 35584 4264 35590 4276
rect 35989 4267 36047 4273
rect 35989 4264 36001 4267
rect 35584 4236 36001 4264
rect 35584 4224 35590 4236
rect 35989 4233 36001 4236
rect 36035 4233 36047 4267
rect 35989 4227 36047 4233
rect 31665 4199 31723 4205
rect 31665 4196 31677 4199
rect 24886 4168 28304 4196
rect 29486 4168 31677 4196
rect 31665 4165 31677 4168
rect 31711 4165 31723 4199
rect 31665 4159 31723 4165
rect 31864 4168 32352 4196
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 20530 4128 20536 4140
rect 20303 4100 20536 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 21085 4131 21143 4137
rect 21085 4097 21097 4131
rect 21131 4097 21143 4131
rect 21085 4091 21143 4097
rect 22373 4131 22431 4137
rect 22373 4097 22385 4131
rect 22419 4128 22431 4131
rect 22830 4128 22836 4140
rect 22419 4100 22836 4128
rect 22419 4097 22431 4100
rect 22373 4091 22431 4097
rect 21100 3992 21128 4091
rect 22830 4088 22836 4100
rect 22888 4088 22894 4140
rect 22925 4131 22983 4137
rect 22925 4097 22937 4131
rect 22971 4128 22983 4131
rect 23198 4128 23204 4140
rect 22971 4100 23204 4128
rect 22971 4097 22983 4100
rect 22925 4091 22983 4097
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 25406 4128 25412 4140
rect 25367 4100 25412 4128
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 25498 4088 25504 4140
rect 25556 4128 25562 4140
rect 26421 4131 26479 4137
rect 26421 4128 26433 4131
rect 25556 4100 26433 4128
rect 25556 4088 25562 4100
rect 26421 4097 26433 4100
rect 26467 4097 26479 4131
rect 26421 4091 26479 4097
rect 30190 4088 30196 4140
rect 30248 4128 30254 4140
rect 30742 4128 30748 4140
rect 30248 4100 30748 4128
rect 30248 4088 30254 4100
rect 30742 4088 30748 4100
rect 30800 4088 30806 4140
rect 31110 4128 31116 4140
rect 31071 4100 31116 4128
rect 31110 4088 31116 4100
rect 31168 4088 31174 4140
rect 31757 4131 31815 4137
rect 31757 4097 31769 4131
rect 31803 4126 31815 4131
rect 31864 4126 31892 4168
rect 32324 4137 32352 4168
rect 31803 4098 31892 4126
rect 32309 4131 32367 4137
rect 31803 4097 31815 4098
rect 31757 4091 31815 4097
rect 32309 4097 32321 4131
rect 32355 4128 32367 4131
rect 32858 4128 32864 4140
rect 32355 4100 32864 4128
rect 32355 4097 32367 4100
rect 32309 4091 32367 4097
rect 32858 4088 32864 4100
rect 32916 4128 32922 4140
rect 33137 4131 33195 4137
rect 33137 4128 33149 4131
rect 32916 4100 33149 4128
rect 32916 4088 32922 4100
rect 33137 4097 33149 4100
rect 33183 4097 33195 4131
rect 33778 4128 33784 4140
rect 33739 4100 33784 4128
rect 33137 4091 33195 4097
rect 33778 4088 33784 4100
rect 33836 4128 33842 4140
rect 34238 4128 34244 4140
rect 33836 4100 34244 4128
rect 33836 4088 33842 4100
rect 34238 4088 34244 4100
rect 34296 4128 34302 4140
rect 34425 4131 34483 4137
rect 34425 4128 34437 4131
rect 34296 4100 34437 4128
rect 34296 4088 34302 4100
rect 34425 4097 34437 4100
rect 34471 4097 34483 4131
rect 38010 4128 38016 4140
rect 37971 4100 38016 4128
rect 34425 4091 34483 4097
rect 38010 4088 38016 4100
rect 38068 4088 38074 4140
rect 23382 4060 23388 4072
rect 23343 4032 23388 4060
rect 23382 4020 23388 4032
rect 23440 4020 23446 4072
rect 23661 4063 23719 4069
rect 23661 4029 23673 4063
rect 23707 4060 23719 4063
rect 25516 4060 25544 4088
rect 23707 4032 25544 4060
rect 23707 4029 23719 4032
rect 23661 4023 23719 4029
rect 27338 4020 27344 4072
rect 27396 4060 27402 4072
rect 28445 4063 28503 4069
rect 28445 4060 28457 4063
rect 27396 4032 28457 4060
rect 27396 4020 27402 4032
rect 28445 4029 28457 4032
rect 28491 4029 28503 4063
rect 29914 4060 29920 4072
rect 29875 4032 29920 4060
rect 28445 4023 28503 4029
rect 29914 4020 29920 4032
rect 29972 4020 29978 4072
rect 30282 4020 30288 4072
rect 30340 4060 30346 4072
rect 34333 4063 34391 4069
rect 34333 4060 34345 4063
rect 30340 4032 34345 4060
rect 30340 4020 30346 4032
rect 34333 4029 34345 4032
rect 34379 4029 34391 4063
rect 36541 4063 36599 4069
rect 36541 4060 36553 4063
rect 34333 4023 34391 4029
rect 34440 4032 36553 4060
rect 21100 3964 23520 3992
rect 1486 3884 1492 3936
rect 1544 3924 1550 3936
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 1544 3896 1593 3924
rect 1544 3884 1550 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 1581 3887 1639 3893
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 20993 3927 21051 3933
rect 20993 3924 21005 3927
rect 20680 3896 21005 3924
rect 20680 3884 20686 3896
rect 20993 3893 21005 3896
rect 21039 3893 21051 3927
rect 23492 3924 23520 3964
rect 24762 3952 24768 4004
rect 24820 3992 24826 4004
rect 33045 3995 33103 4001
rect 33045 3992 33057 3995
rect 24820 3964 28580 3992
rect 24820 3952 24826 3964
rect 26234 3924 26240 3936
rect 23492 3896 26240 3924
rect 20993 3887 21051 3893
rect 26234 3884 26240 3896
rect 26292 3884 26298 3936
rect 27246 3924 27252 3936
rect 27207 3896 27252 3924
rect 27246 3884 27252 3896
rect 27304 3924 27310 3936
rect 27709 3927 27767 3933
rect 27709 3924 27721 3927
rect 27304 3896 27721 3924
rect 27304 3884 27310 3896
rect 27709 3893 27721 3896
rect 27755 3893 27767 3927
rect 28552 3924 28580 3964
rect 30116 3964 33057 3992
rect 30116 3924 30144 3964
rect 33045 3961 33057 3964
rect 33091 3961 33103 3995
rect 34440 3992 34468 4032
rect 36541 4029 36553 4032
rect 36587 4029 36599 4063
rect 36541 4023 36599 4029
rect 37461 3995 37519 4001
rect 37461 3992 37473 3995
rect 33045 3955 33103 3961
rect 33152 3964 34468 3992
rect 35544 3964 37473 3992
rect 28552 3896 30144 3924
rect 27709 3887 27767 3893
rect 30190 3884 30196 3936
rect 30248 3924 30254 3936
rect 31021 3927 31079 3933
rect 31021 3924 31033 3927
rect 30248 3896 31033 3924
rect 30248 3884 30254 3896
rect 31021 3893 31033 3896
rect 31067 3893 31079 3927
rect 31021 3887 31079 3893
rect 31202 3884 31208 3936
rect 31260 3924 31266 3936
rect 32214 3924 32220 3936
rect 31260 3896 32220 3924
rect 31260 3884 31266 3896
rect 32214 3884 32220 3896
rect 32272 3884 32278 3936
rect 32398 3924 32404 3936
rect 32359 3896 32404 3924
rect 32398 3884 32404 3896
rect 32456 3884 32462 3936
rect 32490 3884 32496 3936
rect 32548 3924 32554 3936
rect 33152 3924 33180 3964
rect 35544 3936 35572 3964
rect 37461 3961 37473 3964
rect 37507 3961 37519 3995
rect 37461 3955 37519 3961
rect 33686 3924 33692 3936
rect 32548 3896 33180 3924
rect 33647 3896 33692 3924
rect 32548 3884 32554 3896
rect 33686 3884 33692 3896
rect 33744 3884 33750 3936
rect 34146 3884 34152 3936
rect 34204 3924 34210 3936
rect 34882 3924 34888 3936
rect 34204 3896 34888 3924
rect 34204 3884 34210 3896
rect 34882 3884 34888 3896
rect 34940 3924 34946 3936
rect 35437 3927 35495 3933
rect 35437 3924 35449 3927
rect 34940 3896 35449 3924
rect 34940 3884 34946 3896
rect 35437 3893 35449 3896
rect 35483 3924 35495 3927
rect 35526 3924 35532 3936
rect 35483 3896 35532 3924
rect 35483 3893 35495 3896
rect 35437 3887 35495 3893
rect 35526 3884 35532 3896
rect 35584 3884 35590 3936
rect 37182 3884 37188 3936
rect 37240 3924 37246 3936
rect 38197 3927 38255 3933
rect 38197 3924 38209 3927
rect 37240 3896 38209 3924
rect 37240 3884 37246 3896
rect 38197 3893 38209 3896
rect 38243 3893 38255 3927
rect 38197 3887 38255 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 20438 3720 20444 3732
rect 20399 3692 20444 3720
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 20530 3680 20536 3732
rect 20588 3720 20594 3732
rect 21361 3723 21419 3729
rect 21361 3720 21373 3723
rect 20588 3692 21373 3720
rect 20588 3680 20594 3692
rect 21361 3689 21373 3692
rect 21407 3720 21419 3723
rect 28626 3720 28632 3732
rect 21407 3692 26740 3720
rect 28587 3692 28632 3720
rect 21407 3689 21419 3692
rect 21361 3683 21419 3689
rect 24118 3612 24124 3664
rect 24176 3652 24182 3664
rect 24176 3624 24716 3652
rect 24176 3612 24182 3624
rect 20622 3584 20628 3596
rect 20583 3556 20628 3584
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 24688 3584 24716 3624
rect 24857 3587 24915 3593
rect 24857 3584 24869 3587
rect 24688 3556 24869 3584
rect 24857 3553 24869 3556
rect 24903 3553 24915 3587
rect 24857 3547 24915 3553
rect 24946 3544 24952 3596
rect 25004 3584 25010 3596
rect 26418 3584 26424 3596
rect 25004 3556 26424 3584
rect 25004 3544 25010 3556
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 19705 3519 19763 3525
rect 1903 3488 6914 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 1578 3408 1584 3460
rect 1636 3448 1642 3460
rect 2317 3451 2375 3457
rect 2317 3448 2329 3451
rect 1636 3420 2329 3448
rect 1636 3408 1642 3420
rect 2317 3417 2329 3420
rect 2363 3417 2375 3451
rect 2317 3411 2375 3417
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 6886 3380 6914 3488
rect 19705 3485 19717 3519
rect 19751 3516 19763 3519
rect 20530 3516 20536 3528
rect 19751 3488 20536 3516
rect 19751 3485 19763 3488
rect 19705 3479 19763 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20809 3519 20867 3525
rect 20809 3485 20821 3519
rect 20855 3516 20867 3519
rect 21358 3516 21364 3528
rect 20855 3488 21364 3516
rect 20855 3485 20867 3488
rect 20809 3479 20867 3485
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 22186 3476 22192 3528
rect 22244 3516 22250 3528
rect 22281 3519 22339 3525
rect 22281 3516 22293 3519
rect 22244 3488 22293 3516
rect 22244 3476 22250 3488
rect 22281 3485 22293 3488
rect 22327 3485 22339 3519
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 22281 3479 22339 3485
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 22557 3451 22615 3457
rect 22557 3417 22569 3451
rect 22603 3448 22615 3451
rect 22646 3448 22652 3460
rect 22603 3420 22652 3448
rect 22603 3417 22615 3420
rect 22557 3411 22615 3417
rect 22646 3408 22652 3420
rect 22704 3408 22710 3460
rect 24762 3448 24768 3460
rect 23782 3420 24768 3448
rect 24762 3408 24768 3420
rect 24820 3408 24826 3460
rect 26602 3448 26608 3460
rect 26082 3420 26608 3448
rect 26602 3408 26608 3420
rect 26660 3408 26666 3460
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 6886 3352 19533 3380
rect 19521 3349 19533 3352
rect 19567 3349 19579 3383
rect 19521 3343 19579 3349
rect 24029 3383 24087 3389
rect 24029 3349 24041 3383
rect 24075 3380 24087 3383
rect 26142 3380 26148 3392
rect 24075 3352 26148 3380
rect 24075 3349 24087 3352
rect 24029 3343 24087 3349
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 26326 3380 26332 3392
rect 26287 3352 26332 3380
rect 26326 3340 26332 3352
rect 26384 3340 26390 3392
rect 26712 3380 26740 3692
rect 28626 3680 28632 3692
rect 28684 3720 28690 3732
rect 34241 3723 34299 3729
rect 34241 3720 34253 3723
rect 28684 3692 28994 3720
rect 28684 3680 28690 3692
rect 28966 3664 28994 3692
rect 29196 3692 34253 3720
rect 28966 3624 29000 3664
rect 28994 3612 29000 3624
rect 29052 3612 29058 3664
rect 26786 3544 26792 3596
rect 26844 3584 26850 3596
rect 26881 3587 26939 3593
rect 26881 3584 26893 3587
rect 26844 3556 26893 3584
rect 26844 3544 26850 3556
rect 26881 3553 26893 3556
rect 26927 3584 26939 3587
rect 27246 3584 27252 3596
rect 26927 3556 27252 3584
rect 26927 3553 26939 3556
rect 26881 3547 26939 3553
rect 27246 3544 27252 3556
rect 27304 3544 27310 3596
rect 29196 3584 29224 3692
rect 34241 3689 34253 3692
rect 34287 3689 34299 3723
rect 34241 3683 34299 3689
rect 34422 3680 34428 3732
rect 34480 3720 34486 3732
rect 34977 3723 35035 3729
rect 34977 3720 34989 3723
rect 34480 3692 34989 3720
rect 34480 3680 34486 3692
rect 34977 3689 34989 3692
rect 35023 3689 35035 3723
rect 35526 3720 35532 3732
rect 35487 3692 35532 3720
rect 34977 3683 35035 3689
rect 35526 3680 35532 3692
rect 35584 3720 35590 3732
rect 36081 3723 36139 3729
rect 36081 3720 36093 3723
rect 35584 3692 36093 3720
rect 35584 3680 35590 3692
rect 36081 3689 36093 3692
rect 36127 3689 36139 3723
rect 36081 3683 36139 3689
rect 31294 3612 31300 3664
rect 31352 3652 31358 3664
rect 31481 3655 31539 3661
rect 31481 3652 31493 3655
rect 31352 3624 31493 3652
rect 31352 3612 31358 3624
rect 31481 3621 31493 3624
rect 31527 3652 31539 3655
rect 33689 3655 33747 3661
rect 33689 3652 33701 3655
rect 31527 3624 32076 3652
rect 31527 3621 31539 3624
rect 31481 3615 31539 3621
rect 28276 3556 29224 3584
rect 28276 3502 28304 3556
rect 29270 3544 29276 3596
rect 29328 3584 29334 3596
rect 30009 3587 30067 3593
rect 30009 3584 30021 3587
rect 29328 3556 30021 3584
rect 29328 3544 29334 3556
rect 30009 3553 30021 3556
rect 30055 3553 30067 3587
rect 30009 3547 30067 3553
rect 30558 3544 30564 3596
rect 30616 3584 30622 3596
rect 31202 3584 31208 3596
rect 30616 3556 31208 3584
rect 30616 3544 30622 3556
rect 31202 3544 31208 3556
rect 31260 3544 31266 3596
rect 32048 3584 32076 3624
rect 33244 3624 33701 3652
rect 32217 3587 32275 3593
rect 32217 3584 32229 3587
rect 32048 3556 32229 3584
rect 32217 3553 32229 3556
rect 32263 3553 32275 3587
rect 32217 3547 32275 3553
rect 32582 3544 32588 3596
rect 32640 3584 32646 3596
rect 33244 3584 33272 3624
rect 33689 3621 33701 3624
rect 33735 3652 33747 3655
rect 35986 3652 35992 3664
rect 33735 3624 35992 3652
rect 33735 3621 33747 3624
rect 33689 3615 33747 3621
rect 35986 3612 35992 3624
rect 36044 3612 36050 3664
rect 34514 3584 34520 3596
rect 32640 3556 33272 3584
rect 33336 3556 34520 3584
rect 32640 3544 32646 3556
rect 28994 3476 29000 3528
rect 29052 3516 29058 3528
rect 29733 3519 29791 3525
rect 29733 3516 29745 3519
rect 29052 3488 29745 3516
rect 29052 3476 29058 3488
rect 29733 3485 29745 3488
rect 29779 3485 29791 3519
rect 31570 3516 31576 3528
rect 31142 3488 31576 3516
rect 29733 3479 29791 3485
rect 31570 3476 31576 3488
rect 31628 3476 31634 3528
rect 31938 3516 31944 3528
rect 31899 3488 31944 3516
rect 31938 3476 31944 3488
rect 31996 3476 32002 3528
rect 33336 3502 33364 3556
rect 34514 3544 34520 3556
rect 34572 3544 34578 3596
rect 34238 3476 34244 3528
rect 34296 3516 34302 3528
rect 34333 3519 34391 3525
rect 34333 3516 34345 3519
rect 34296 3488 34345 3516
rect 34296 3476 34302 3488
rect 34333 3485 34345 3488
rect 34379 3516 34391 3519
rect 34882 3516 34888 3528
rect 34379 3488 34888 3516
rect 34379 3485 34391 3488
rect 34333 3479 34391 3485
rect 34882 3476 34888 3488
rect 34940 3476 34946 3528
rect 38013 3519 38071 3525
rect 38013 3485 38025 3519
rect 38059 3485 38071 3519
rect 38286 3516 38292 3528
rect 38247 3488 38292 3516
rect 38013 3479 38071 3485
rect 27154 3408 27160 3460
rect 27212 3448 27218 3460
rect 38028 3448 38056 3479
rect 38286 3476 38292 3488
rect 38344 3476 38350 3528
rect 27212 3420 27257 3448
rect 28460 3420 29224 3448
rect 27212 3408 27218 3420
rect 28460 3380 28488 3420
rect 26712 3352 28488 3380
rect 28718 3340 28724 3392
rect 28776 3380 28782 3392
rect 29089 3383 29147 3389
rect 29089 3380 29101 3383
rect 28776 3352 29101 3380
rect 28776 3340 28782 3352
rect 29089 3349 29101 3352
rect 29135 3349 29147 3383
rect 29196 3380 29224 3420
rect 31312 3420 31754 3448
rect 31312 3380 31340 3420
rect 29196 3352 31340 3380
rect 31726 3380 31754 3420
rect 33612 3420 38056 3448
rect 33612 3380 33640 3420
rect 36630 3380 36636 3392
rect 31726 3352 33640 3380
rect 36591 3352 36636 3380
rect 29089 3343 29147 3349
rect 36630 3340 36636 3352
rect 36688 3340 36694 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 6886 3148 20637 3176
rect 3142 3068 3148 3120
rect 3200 3108 3206 3120
rect 3329 3111 3387 3117
rect 3329 3108 3341 3111
rect 3200 3080 3341 3108
rect 3200 3068 3206 3080
rect 3329 3077 3341 3080
rect 3375 3108 3387 3111
rect 6886 3108 6914 3148
rect 20625 3145 20637 3148
rect 20671 3145 20683 3179
rect 21358 3176 21364 3188
rect 21319 3148 21364 3176
rect 20625 3139 20683 3145
rect 21358 3136 21364 3148
rect 21416 3136 21422 3188
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 23382 3176 23388 3188
rect 22244 3148 23388 3176
rect 22244 3136 22250 3148
rect 3375 3080 6914 3108
rect 19521 3111 19579 3117
rect 3375 3077 3387 3080
rect 3329 3071 3387 3077
rect 19521 3077 19533 3111
rect 19567 3108 19579 3111
rect 21266 3108 21272 3120
rect 19567 3080 21272 3108
rect 19567 3077 19579 3080
rect 19521 3071 19579 3077
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 18322 3040 18328 3052
rect 17543 3012 18328 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 18322 3000 18328 3012
rect 18380 3040 18386 3052
rect 19242 3040 19248 3052
rect 18380 3012 19248 3040
rect 18380 3000 18386 3012
rect 19242 3000 19248 3012
rect 19300 3000 19306 3052
rect 14 2932 20 2984
rect 72 2972 78 2984
rect 1486 2972 1492 2984
rect 72 2944 1492 2972
rect 72 2932 78 2944
rect 1486 2932 1492 2944
rect 1544 2972 1550 2984
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 1544 2944 1593 2972
rect 1544 2932 1550 2944
rect 1581 2941 1593 2944
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 19536 2972 19564 3071
rect 19996 3049 20024 3080
rect 21266 3068 21272 3080
rect 21324 3068 21330 3120
rect 22557 3111 22615 3117
rect 22557 3077 22569 3111
rect 22603 3108 22615 3111
rect 23106 3108 23112 3120
rect 22603 3080 23112 3108
rect 22603 3077 22615 3080
rect 22557 3071 22615 3077
rect 23106 3068 23112 3080
rect 23164 3068 23170 3120
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21450 3040 21456 3052
rect 20855 3012 21456 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21450 3000 21456 3012
rect 21508 3000 21514 3052
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3040 22155 3043
rect 22741 3043 22799 3049
rect 22741 3040 22753 3043
rect 22143 3012 22753 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 22741 3009 22753 3012
rect 22787 3040 22799 3043
rect 23014 3040 23020 3052
rect 22787 3012 23020 3040
rect 22787 3009 22799 3012
rect 22741 3003 22799 3009
rect 23014 3000 23020 3012
rect 23072 3000 23078 3052
rect 23308 3049 23336 3148
rect 23382 3136 23388 3148
rect 23440 3136 23446 3188
rect 26326 3136 26332 3188
rect 26384 3176 26390 3188
rect 26513 3179 26571 3185
rect 26513 3176 26525 3179
rect 26384 3148 26525 3176
rect 26384 3136 26390 3148
rect 26513 3145 26525 3148
rect 26559 3145 26571 3179
rect 26513 3139 26571 3145
rect 26602 3136 26608 3188
rect 26660 3176 26666 3188
rect 27246 3176 27252 3188
rect 26660 3148 26924 3176
rect 27207 3148 27252 3176
rect 26660 3136 26666 3148
rect 23569 3111 23627 3117
rect 23569 3077 23581 3111
rect 23615 3108 23627 3111
rect 23658 3108 23664 3120
rect 23615 3080 23664 3108
rect 23615 3077 23627 3080
rect 23569 3071 23627 3077
rect 23658 3068 23664 3080
rect 23716 3068 23722 3120
rect 25222 3108 25228 3120
rect 24794 3080 25228 3108
rect 25222 3068 25228 3080
rect 25280 3068 25286 3120
rect 25317 3111 25375 3117
rect 25317 3077 25329 3111
rect 25363 3108 25375 3111
rect 25498 3108 25504 3120
rect 25363 3080 25504 3108
rect 25363 3077 25375 3080
rect 25317 3071 25375 3077
rect 25498 3068 25504 3080
rect 25556 3068 25562 3120
rect 23293 3043 23351 3049
rect 23293 3009 23305 3043
rect 23339 3009 23351 3043
rect 23293 3003 23351 3009
rect 24854 3000 24860 3052
rect 24912 3040 24918 3052
rect 25590 3040 25596 3052
rect 24912 3012 25596 3040
rect 24912 3000 24918 3012
rect 25590 3000 25596 3012
rect 25648 3000 25654 3052
rect 25777 3043 25835 3049
rect 25777 3009 25789 3043
rect 25823 3009 25835 3043
rect 25777 3003 25835 3009
rect 25792 2972 25820 3003
rect 25866 3000 25872 3052
rect 25924 3040 25930 3052
rect 26896 3040 26924 3148
rect 27246 3136 27252 3148
rect 27304 3136 27310 3188
rect 28074 3176 28080 3188
rect 28035 3148 28080 3176
rect 28074 3136 28080 3148
rect 28132 3136 28138 3188
rect 29086 3176 29092 3188
rect 28184 3148 29092 3176
rect 28184 3117 28212 3148
rect 29086 3136 29092 3148
rect 29144 3176 29150 3188
rect 31386 3176 31392 3188
rect 29144 3148 31392 3176
rect 29144 3136 29150 3148
rect 31386 3136 31392 3148
rect 31444 3136 31450 3188
rect 34146 3176 34152 3188
rect 31956 3148 34152 3176
rect 31956 3120 31984 3148
rect 34146 3136 34152 3148
rect 34204 3136 34210 3188
rect 35342 3176 35348 3188
rect 35303 3148 35348 3176
rect 35342 3136 35348 3148
rect 35400 3136 35406 3188
rect 35526 3136 35532 3188
rect 35584 3176 35590 3188
rect 36357 3179 36415 3185
rect 36357 3176 36369 3179
rect 35584 3148 36369 3176
rect 35584 3136 35590 3148
rect 36357 3145 36369 3148
rect 36403 3145 36415 3179
rect 36357 3139 36415 3145
rect 28169 3111 28227 3117
rect 28169 3077 28181 3111
rect 28215 3077 28227 3111
rect 30190 3108 30196 3120
rect 30038 3080 30196 3108
rect 28169 3071 28227 3077
rect 30190 3068 30196 3080
rect 30248 3068 30254 3120
rect 31938 3108 31944 3120
rect 30760 3080 31944 3108
rect 30760 3052 30788 3080
rect 31938 3068 31944 3080
rect 31996 3068 32002 3120
rect 32398 3068 32404 3120
rect 32456 3108 32462 3120
rect 32456 3080 32614 3108
rect 32456 3068 32462 3080
rect 25924 3012 26832 3040
rect 26896 3012 28856 3040
rect 25924 3000 25930 3012
rect 1903 2944 19564 2972
rect 20180 2944 25820 2972
rect 26804 2972 26832 3012
rect 28718 2972 28724 2984
rect 26804 2944 28724 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 5534 2864 5540 2916
rect 5592 2904 5598 2916
rect 5721 2907 5779 2913
rect 5721 2904 5733 2907
rect 5592 2876 5733 2904
rect 5592 2864 5598 2876
rect 5721 2873 5733 2876
rect 5767 2904 5779 2907
rect 20070 2904 20076 2916
rect 5767 2876 20076 2904
rect 5767 2873 5779 2876
rect 5721 2867 5779 2873
rect 20070 2864 20076 2876
rect 20128 2864 20134 2916
rect 20180 2913 20208 2944
rect 28718 2932 28724 2944
rect 28776 2932 28782 2984
rect 28828 2972 28856 3012
rect 30742 3000 30748 3052
rect 30800 3040 30806 3052
rect 31389 3043 31447 3049
rect 31389 3040 31401 3043
rect 30800 3012 30845 3040
rect 31128 3012 31401 3040
rect 30800 3000 30806 3012
rect 30374 2972 30380 2984
rect 28828 2944 30380 2972
rect 30374 2932 30380 2944
rect 30432 2932 30438 2984
rect 30466 2932 30472 2984
rect 30524 2972 30530 2984
rect 30524 2944 30569 2972
rect 30524 2932 30530 2944
rect 20165 2907 20223 2913
rect 20165 2873 20177 2907
rect 20211 2873 20223 2907
rect 20165 2867 20223 2873
rect 25222 2864 25228 2916
rect 25280 2904 25286 2916
rect 25280 2876 26832 2904
rect 25280 2864 25286 2876
rect 3786 2836 3792 2848
rect 3747 2808 3792 2836
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 17313 2839 17371 2845
rect 17313 2836 17325 2839
rect 14608 2808 17325 2836
rect 14608 2796 14614 2808
rect 17313 2805 17325 2808
rect 17359 2805 17371 2839
rect 17313 2799 17371 2805
rect 18049 2839 18107 2845
rect 18049 2805 18061 2839
rect 18095 2836 18107 2839
rect 18322 2836 18328 2848
rect 18095 2808 18328 2836
rect 18095 2805 18107 2808
rect 18049 2799 18107 2805
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 23658 2796 23664 2848
rect 23716 2836 23722 2848
rect 24762 2836 24768 2848
rect 23716 2808 24768 2836
rect 23716 2796 23722 2808
rect 24762 2796 24768 2808
rect 24820 2796 24826 2848
rect 25130 2796 25136 2848
rect 25188 2836 25194 2848
rect 25961 2839 26019 2845
rect 25961 2836 25973 2839
rect 25188 2808 25973 2836
rect 25188 2796 25194 2808
rect 25961 2805 25973 2808
rect 26007 2805 26019 2839
rect 26804 2836 26832 2876
rect 27062 2864 27068 2916
rect 27120 2904 27126 2916
rect 27246 2904 27252 2916
rect 27120 2876 27252 2904
rect 27120 2864 27126 2876
rect 27246 2864 27252 2876
rect 27304 2904 27310 2916
rect 28994 2904 29000 2916
rect 27304 2876 29000 2904
rect 27304 2864 27310 2876
rect 28994 2864 29000 2876
rect 29052 2864 29058 2916
rect 30098 2836 30104 2848
rect 26804 2808 30104 2836
rect 25961 2799 26019 2805
rect 30098 2796 30104 2808
rect 30156 2796 30162 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 31128 2836 31156 3012
rect 31389 3009 31401 3012
rect 31435 3040 31447 3043
rect 32490 3040 32496 3052
rect 31435 3012 32496 3040
rect 31435 3009 31447 3012
rect 31389 3003 31447 3009
rect 32490 3000 32496 3012
rect 32548 3000 32554 3052
rect 31205 2975 31263 2981
rect 31205 2941 31217 2975
rect 31251 2972 31263 2975
rect 31478 2972 31484 2984
rect 31251 2944 31484 2972
rect 31251 2941 31263 2944
rect 31205 2935 31263 2941
rect 31478 2932 31484 2944
rect 31536 2932 31542 2984
rect 31846 2932 31852 2984
rect 31904 2972 31910 2984
rect 33781 2975 33839 2981
rect 33781 2972 33793 2975
rect 31904 2944 33793 2972
rect 31904 2932 31910 2944
rect 33781 2941 33793 2944
rect 33827 2941 33839 2975
rect 33781 2935 33839 2941
rect 34057 2975 34115 2981
rect 34057 2941 34069 2975
rect 34103 2972 34115 2975
rect 34164 2972 34192 3136
rect 34606 3108 34612 3120
rect 34567 3080 34612 3108
rect 34606 3068 34612 3080
rect 34664 3068 34670 3120
rect 34701 3043 34759 3049
rect 34701 3009 34713 3043
rect 34747 3040 34759 3043
rect 34882 3040 34888 3052
rect 34747 3012 34888 3040
rect 34747 3009 34759 3012
rect 34701 3003 34759 3009
rect 34882 3000 34888 3012
rect 34940 3000 34946 3052
rect 35161 3043 35219 3049
rect 35161 3009 35173 3043
rect 35207 3040 35219 3043
rect 36538 3040 36544 3052
rect 35207 3012 36544 3040
rect 35207 3009 35219 3012
rect 35161 3003 35219 3009
rect 34103 2944 34192 2972
rect 34103 2941 34115 2944
rect 34057 2935 34115 2941
rect 34238 2932 34244 2984
rect 34296 2972 34302 2984
rect 35176 2972 35204 3003
rect 36538 3000 36544 3012
rect 36596 3000 36602 3052
rect 38010 3040 38016 3052
rect 37971 3012 38016 3040
rect 38010 3000 38016 3012
rect 38068 3000 38074 3052
rect 38194 3000 38200 3052
rect 38252 3040 38258 3052
rect 38289 3043 38347 3049
rect 38289 3040 38301 3043
rect 38252 3012 38301 3040
rect 38252 3000 38258 3012
rect 38289 3009 38301 3012
rect 38335 3040 38347 3043
rect 39298 3040 39304 3052
rect 38335 3012 39304 3040
rect 38335 3009 38347 3012
rect 38289 3003 38347 3009
rect 39298 3000 39304 3012
rect 39356 3000 39362 3052
rect 34296 2944 35204 2972
rect 34296 2932 34302 2944
rect 31386 2864 31392 2916
rect 31444 2904 31450 2916
rect 35805 2907 35863 2913
rect 35805 2904 35817 2907
rect 31444 2876 32444 2904
rect 31444 2864 31450 2876
rect 32306 2836 32312 2848
rect 30340 2808 31156 2836
rect 32267 2808 32312 2836
rect 30340 2796 30346 2808
rect 32306 2796 32312 2808
rect 32364 2796 32370 2848
rect 32416 2836 32444 2876
rect 33980 2876 35817 2904
rect 33980 2836 34008 2876
rect 35805 2873 35817 2876
rect 35851 2873 35863 2907
rect 35805 2867 35863 2873
rect 32416 2808 34008 2836
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 10778 2632 10784 2644
rect 4203 2604 10784 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 19150 2632 19156 2644
rect 14507 2604 19156 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 22922 2592 22928 2644
rect 22980 2632 22986 2644
rect 26326 2632 26332 2644
rect 22980 2604 26332 2632
rect 22980 2592 22986 2604
rect 26326 2592 26332 2604
rect 26384 2592 26390 2644
rect 26510 2592 26516 2644
rect 26568 2632 26574 2644
rect 27249 2635 27307 2641
rect 27249 2632 27261 2635
rect 26568 2604 27261 2632
rect 26568 2592 26574 2604
rect 27249 2601 27261 2604
rect 27295 2601 27307 2635
rect 27249 2595 27307 2601
rect 29362 2592 29368 2644
rect 29420 2632 29426 2644
rect 29733 2635 29791 2641
rect 29733 2632 29745 2635
rect 29420 2604 29745 2632
rect 29420 2592 29426 2604
rect 29733 2601 29745 2604
rect 29779 2601 29791 2635
rect 29733 2595 29791 2601
rect 30650 2592 30656 2644
rect 30708 2632 30714 2644
rect 33505 2635 33563 2641
rect 33505 2632 33517 2635
rect 30708 2604 33517 2632
rect 30708 2592 30714 2604
rect 33505 2601 33517 2604
rect 33551 2601 33563 2635
rect 33505 2595 33563 2601
rect 35526 2592 35532 2644
rect 35584 2632 35590 2644
rect 35621 2635 35679 2641
rect 35621 2632 35633 2635
rect 35584 2604 35633 2632
rect 35584 2592 35590 2604
rect 35621 2601 35633 2604
rect 35667 2601 35679 2635
rect 35621 2595 35679 2601
rect 9401 2567 9459 2573
rect 9401 2533 9413 2567
rect 9447 2564 9459 2567
rect 12066 2564 12072 2576
rect 9447 2536 12072 2564
rect 9447 2533 9459 2536
rect 9401 2527 9459 2533
rect 12066 2524 12072 2536
rect 12124 2524 12130 2576
rect 21542 2564 21548 2576
rect 12544 2536 21548 2564
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2496 1915 2499
rect 1946 2496 1952 2508
rect 1903 2468 1952 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 10318 2456 10324 2508
rect 10376 2496 10382 2508
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 10376 2468 11161 2496
rect 10376 2456 10382 2468
rect 11149 2465 11161 2468
rect 11195 2496 11207 2499
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11195 2468 11713 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11701 2459 11759 2465
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 3142 2428 3148 2440
rect 3103 2400 3148 2428
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 5534 2428 5540 2440
rect 5495 2400 5540 2428
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2428 7530 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7524 2400 7941 2428
rect 7524 2388 7530 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 12544 2428 12572 2536
rect 21542 2524 21548 2536
rect 21600 2524 21606 2576
rect 36449 2567 36507 2573
rect 36449 2533 36461 2567
rect 36495 2564 36507 2567
rect 37274 2564 37280 2576
rect 36495 2536 37280 2564
rect 36495 2533 36507 2536
rect 36449 2527 36507 2533
rect 37274 2524 37280 2536
rect 37332 2524 37338 2576
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 14660 2468 18337 2496
rect 10919 2400 12572 2428
rect 12621 2431 12679 2437
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 12621 2397 12633 2431
rect 12667 2428 12679 2431
rect 14550 2428 14556 2440
rect 12667 2400 14556 2428
rect 12667 2397 12679 2400
rect 12621 2391 12679 2397
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 3786 2360 3792 2372
rect 3292 2332 3792 2360
rect 3292 2320 3298 2332
rect 3786 2320 3792 2332
rect 3844 2360 3850 2372
rect 4065 2363 4123 2369
rect 4065 2360 4077 2363
rect 3844 2332 4077 2360
rect 3844 2320 3850 2332
rect 4065 2329 4077 2332
rect 4111 2329 4123 2363
rect 4065 2323 4123 2329
rect 8573 2363 8631 2369
rect 8573 2329 8585 2363
rect 8619 2360 8631 2363
rect 9030 2360 9036 2372
rect 8619 2332 9036 2360
rect 8619 2329 8631 2332
rect 8573 2323 8631 2329
rect 9030 2320 9036 2332
rect 9088 2360 9094 2372
rect 9217 2363 9275 2369
rect 9217 2360 9229 2363
rect 9088 2332 9229 2360
rect 9088 2320 9094 2332
rect 9217 2329 9229 2332
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 9858 2320 9864 2372
rect 9916 2360 9922 2372
rect 13725 2363 13783 2369
rect 9916 2332 12572 2360
rect 9916 2320 9922 2332
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 2961 2295 3019 2301
rect 2961 2292 2973 2295
rect 1360 2264 2973 2292
rect 1360 2252 1366 2264
rect 2961 2261 2973 2264
rect 3007 2261 3019 2295
rect 2961 2255 3019 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 5224 2264 5365 2292
rect 5224 2252 5230 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 7156 2264 7297 2292
rect 7156 2252 7162 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12308 2264 12449 2292
rect 12308 2252 12314 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12544 2292 12572 2332
rect 13725 2329 13737 2363
rect 13771 2360 13783 2363
rect 14182 2360 14188 2372
rect 13771 2332 14188 2360
rect 13771 2329 13783 2332
rect 13725 2323 13783 2329
rect 14182 2320 14188 2332
rect 14240 2360 14246 2372
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 14240 2332 14381 2360
rect 14240 2320 14246 2332
rect 14369 2329 14381 2332
rect 14415 2329 14427 2363
rect 14369 2323 14427 2329
rect 14660 2292 14688 2468
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 21818 2496 21824 2508
rect 18325 2459 18383 2465
rect 19720 2468 21824 2496
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 15988 2400 16865 2428
rect 15988 2388 15994 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 18046 2428 18052 2440
rect 17959 2400 18052 2428
rect 16853 2391 16911 2397
rect 18046 2388 18052 2400
rect 18104 2428 18110 2440
rect 19720 2437 19748 2468
rect 21818 2456 21824 2468
rect 21876 2456 21882 2508
rect 22186 2496 22192 2508
rect 22147 2468 22192 2496
rect 22186 2456 22192 2468
rect 22244 2456 22250 2508
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2496 22523 2499
rect 22922 2496 22928 2508
rect 22511 2468 22928 2496
rect 22511 2465 22523 2468
rect 22465 2459 22523 2465
rect 22922 2456 22928 2468
rect 22980 2456 22986 2508
rect 23474 2456 23480 2508
rect 23532 2496 23538 2508
rect 24578 2496 24584 2508
rect 23532 2468 24584 2496
rect 23532 2456 23538 2468
rect 24578 2456 24584 2468
rect 24636 2456 24642 2508
rect 26234 2496 26240 2508
rect 25976 2468 26240 2496
rect 19705 2431 19763 2437
rect 18104 2400 18276 2428
rect 18104 2388 18110 2400
rect 18248 2360 18276 2400
rect 19705 2397 19717 2431
rect 19751 2397 19763 2431
rect 21174 2428 21180 2440
rect 21135 2400 21180 2428
rect 19705 2391 19763 2397
rect 21174 2388 21180 2400
rect 21232 2388 21238 2440
rect 25976 2414 26004 2468
rect 26234 2456 26240 2468
rect 26292 2456 26298 2508
rect 26329 2499 26387 2505
rect 26329 2465 26341 2499
rect 26375 2496 26387 2499
rect 26418 2496 26424 2508
rect 26375 2468 26424 2496
rect 26375 2465 26387 2468
rect 26329 2459 26387 2465
rect 26418 2456 26424 2468
rect 26476 2496 26482 2508
rect 27154 2496 27160 2508
rect 26476 2468 27160 2496
rect 26476 2456 26482 2468
rect 27154 2456 27160 2468
rect 27212 2456 27218 2508
rect 27338 2456 27344 2508
rect 27396 2496 27402 2508
rect 28721 2499 28779 2505
rect 28721 2496 28733 2499
rect 27396 2468 28733 2496
rect 27396 2456 27402 2468
rect 28721 2465 28733 2468
rect 28767 2465 28779 2499
rect 28721 2459 28779 2465
rect 28994 2456 29000 2508
rect 29052 2496 29058 2508
rect 31481 2499 31539 2505
rect 29052 2468 29097 2496
rect 29052 2456 29058 2468
rect 31481 2465 31493 2499
rect 31527 2496 31539 2499
rect 31938 2496 31944 2508
rect 31527 2468 31944 2496
rect 31527 2465 31539 2468
rect 31481 2459 31539 2465
rect 31938 2456 31944 2468
rect 31996 2456 32002 2508
rect 37458 2496 37464 2508
rect 37419 2468 37464 2496
rect 37458 2456 37464 2468
rect 37516 2456 37522 2508
rect 37734 2496 37740 2508
rect 37695 2468 37740 2496
rect 37734 2456 37740 2468
rect 37792 2456 37798 2508
rect 32950 2428 32956 2440
rect 32911 2400 32956 2428
rect 32950 2388 32956 2400
rect 33008 2428 33014 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33008 2400 33609 2428
rect 33008 2388 33014 2400
rect 33597 2397 33609 2400
rect 33643 2428 33655 2431
rect 34241 2431 34299 2437
rect 34241 2428 34253 2431
rect 33643 2400 34253 2428
rect 33643 2397 33655 2400
rect 33597 2391 33655 2397
rect 34241 2397 34253 2400
rect 34287 2397 34299 2431
rect 34241 2391 34299 2397
rect 34422 2388 34428 2440
rect 34480 2428 34486 2440
rect 34698 2428 34704 2440
rect 34480 2400 34704 2428
rect 34480 2388 34486 2400
rect 34698 2388 34704 2400
rect 34756 2428 34762 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34756 2400 35081 2428
rect 34756 2388 34762 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35069 2391 35127 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36265 2431 36323 2437
rect 36265 2428 36277 2431
rect 36136 2400 36277 2428
rect 36136 2388 36142 2400
rect 36265 2397 36277 2400
rect 36311 2397 36323 2431
rect 37476 2428 37504 2456
rect 38010 2428 38016 2440
rect 37476 2400 38016 2428
rect 36265 2391 36323 2397
rect 38010 2388 38016 2400
rect 38068 2388 38074 2440
rect 20165 2363 20223 2369
rect 20165 2360 20177 2363
rect 18248 2332 20177 2360
rect 20165 2329 20177 2332
rect 20211 2329 20223 2363
rect 24578 2360 24584 2372
rect 23690 2332 24584 2360
rect 20165 2323 20223 2329
rect 24578 2320 24584 2332
rect 24636 2320 24642 2372
rect 24857 2363 24915 2369
rect 24857 2329 24869 2363
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 12544 2264 14688 2292
rect 12437 2255 12495 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16172 2264 17049 2292
rect 16172 2252 16178 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19521 2295 19579 2301
rect 19521 2292 19533 2295
rect 19392 2264 19533 2292
rect 19392 2252 19398 2264
rect 19521 2261 19533 2264
rect 19567 2261 19579 2295
rect 19521 2255 19579 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 21361 2295 21419 2301
rect 21361 2292 21373 2295
rect 21324 2264 21373 2292
rect 21324 2252 21330 2264
rect 21361 2261 21373 2264
rect 21407 2261 21419 2295
rect 21361 2255 21419 2261
rect 23290 2252 23296 2304
rect 23348 2292 23354 2304
rect 23937 2295 23995 2301
rect 23937 2292 23949 2295
rect 23348 2264 23949 2292
rect 23348 2252 23354 2264
rect 23937 2261 23949 2264
rect 23983 2292 23995 2295
rect 24872 2292 24900 2323
rect 28258 2320 28264 2372
rect 28316 2320 28322 2372
rect 30774 2332 31156 2360
rect 23983 2264 24900 2292
rect 31128 2292 31156 2332
rect 31202 2320 31208 2372
rect 31260 2360 31266 2372
rect 34149 2363 34207 2369
rect 34149 2360 34161 2363
rect 31260 2332 31305 2360
rect 31404 2332 34161 2360
rect 31260 2320 31266 2332
rect 31404 2292 31432 2332
rect 34149 2329 34161 2332
rect 34195 2329 34207 2363
rect 34149 2323 34207 2329
rect 32858 2292 32864 2304
rect 31128 2264 31432 2292
rect 32819 2264 32864 2292
rect 23983 2261 23995 2264
rect 23937 2255 23995 2261
rect 32858 2252 32864 2264
rect 32916 2252 32922 2304
rect 34974 2292 34980 2304
rect 34935 2264 34980 2292
rect 34974 2252 34980 2264
rect 35032 2252 35038 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 24578 2048 24584 2100
rect 24636 2088 24642 2100
rect 32858 2088 32864 2100
rect 24636 2060 32864 2088
rect 24636 2048 24642 2060
rect 32858 2048 32864 2060
rect 32916 2048 32922 2100
rect 18322 1980 18328 2032
rect 18380 2020 18386 2032
rect 34974 2020 34980 2032
rect 18380 1992 34980 2020
rect 18380 1980 18386 1992
rect 34974 1980 34980 1992
rect 35032 1980 35038 2032
rect 26234 1912 26240 1964
rect 26292 1952 26298 1964
rect 33686 1952 33692 1964
rect 26292 1924 33692 1952
rect 26292 1912 26298 1924
rect 33686 1912 33692 1924
rect 33744 1912 33750 1964
rect 28258 1844 28264 1896
rect 28316 1884 28322 1896
rect 33410 1884 33416 1896
rect 28316 1856 33416 1884
rect 28316 1844 28322 1856
rect 33410 1844 33416 1856
rect 33468 1844 33474 1896
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16120 37408 16172 37460
rect 2320 37247 2372 37256
rect 2320 37213 2329 37247
rect 2329 37213 2363 37247
rect 2363 37213 2372 37247
rect 2320 37204 2372 37213
rect 3424 37204 3476 37256
rect 5540 37247 5592 37256
rect 5540 37213 5549 37247
rect 5549 37213 5583 37247
rect 5583 37213 5592 37247
rect 5540 37204 5592 37213
rect 2412 37136 2464 37188
rect 9036 37204 9088 37256
rect 10324 37272 10376 37324
rect 11704 37272 11756 37324
rect 12256 37272 12308 37324
rect 27068 37408 27120 37460
rect 34152 37408 34204 37460
rect 19984 37272 20036 37324
rect 23204 37272 23256 37324
rect 26792 37272 26844 37324
rect 10876 37247 10928 37256
rect 10876 37213 10885 37247
rect 10885 37213 10919 37247
rect 10919 37213 10928 37247
rect 10876 37204 10928 37213
rect 14280 37247 14332 37256
rect 14280 37213 14289 37247
rect 14289 37213 14323 37247
rect 14323 37213 14332 37247
rect 14280 37204 14332 37213
rect 17132 37247 17184 37256
rect 17132 37213 17141 37247
rect 17141 37213 17175 37247
rect 17175 37213 17184 37247
rect 17132 37204 17184 37213
rect 17868 37204 17920 37256
rect 20720 37136 20772 37188
rect 21364 37204 21416 37256
rect 23388 37136 23440 37188
rect 24584 37136 24636 37188
rect 1308 37068 1360 37120
rect 2780 37068 2832 37120
rect 3240 37068 3292 37120
rect 5172 37068 5224 37120
rect 7104 37068 7156 37120
rect 8024 37111 8076 37120
rect 8024 37077 8033 37111
rect 8033 37077 8067 37111
rect 8067 37077 8076 37111
rect 8024 37068 8076 37077
rect 9312 37111 9364 37120
rect 9312 37077 9321 37111
rect 9321 37077 9355 37111
rect 9355 37077 9364 37111
rect 9312 37068 9364 37077
rect 14188 37068 14240 37120
rect 18052 37068 18104 37120
rect 21272 37068 21324 37120
rect 23848 37068 23900 37120
rect 27068 37204 27120 37256
rect 28724 37204 28776 37256
rect 30472 37247 30524 37256
rect 30472 37213 30481 37247
rect 30481 37213 30515 37247
rect 30515 37213 30524 37247
rect 30472 37204 30524 37213
rect 32312 37247 32364 37256
rect 32312 37213 32321 37247
rect 32321 37213 32355 37247
rect 32355 37213 32364 37247
rect 32312 37204 32364 37213
rect 34796 37272 34848 37324
rect 36268 37204 36320 37256
rect 36912 37204 36964 37256
rect 25136 37068 25188 37120
rect 29000 37068 29052 37120
rect 30380 37068 30432 37120
rect 32220 37068 32272 37120
rect 36084 37068 36136 37120
rect 38016 37068 38068 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 3424 36907 3476 36916
rect 3424 36873 3433 36907
rect 3433 36873 3467 36907
rect 3467 36873 3476 36907
rect 3424 36864 3476 36873
rect 11704 36907 11756 36916
rect 11704 36873 11713 36907
rect 11713 36873 11747 36907
rect 11747 36873 11756 36907
rect 11704 36864 11756 36873
rect 17868 36907 17920 36916
rect 17868 36873 17877 36907
rect 17877 36873 17911 36907
rect 17911 36873 17920 36907
rect 17868 36864 17920 36873
rect 20720 36907 20772 36916
rect 20720 36873 20729 36907
rect 20729 36873 20763 36907
rect 20763 36873 20772 36907
rect 20720 36864 20772 36873
rect 21364 36907 21416 36916
rect 21364 36873 21373 36907
rect 21373 36873 21407 36907
rect 21407 36873 21416 36907
rect 21364 36864 21416 36873
rect 32312 36864 32364 36916
rect 39304 36864 39356 36916
rect 20 36796 72 36848
rect 1676 36839 1728 36848
rect 1676 36805 1685 36839
rect 1685 36805 1719 36839
rect 1719 36805 1728 36839
rect 1676 36796 1728 36805
rect 2228 36592 2280 36644
rect 1492 36524 1544 36576
rect 2320 36567 2372 36576
rect 2320 36533 2329 36567
rect 2329 36533 2363 36567
rect 2363 36533 2372 36567
rect 2320 36524 2372 36533
rect 10876 36728 10928 36780
rect 17684 36771 17736 36780
rect 17684 36737 17693 36771
rect 17693 36737 17727 36771
rect 17727 36737 17736 36771
rect 17684 36728 17736 36737
rect 23388 36796 23440 36848
rect 22744 36728 22796 36780
rect 24032 36771 24084 36780
rect 24032 36737 24041 36771
rect 24041 36737 24075 36771
rect 24075 36737 24084 36771
rect 24032 36728 24084 36737
rect 26424 36796 26476 36848
rect 17132 36660 17184 36712
rect 26056 36660 26108 36712
rect 36912 36660 36964 36712
rect 4804 36524 4856 36576
rect 24216 36567 24268 36576
rect 24216 36533 24225 36567
rect 24225 36533 24259 36567
rect 24259 36533 24268 36567
rect 24216 36524 24268 36533
rect 36268 36524 36320 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1676 36320 1728 36372
rect 24216 36320 24268 36372
rect 30472 36320 30524 36372
rect 1860 36159 1912 36168
rect 1860 36125 1869 36159
rect 1869 36125 1903 36159
rect 1903 36125 1912 36159
rect 1860 36116 1912 36125
rect 37740 36116 37792 36168
rect 1676 36023 1728 36032
rect 1676 35989 1685 36023
rect 1685 35989 1719 36023
rect 1719 35989 1728 36023
rect 1676 35980 1728 35989
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1860 35776 1912 35828
rect 38292 35776 38344 35828
rect 2504 35640 2556 35692
rect 37924 35640 37976 35692
rect 2504 35479 2556 35488
rect 2504 35445 2513 35479
rect 2513 35445 2547 35479
rect 2547 35445 2556 35479
rect 2504 35436 2556 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2136 34484 2188 34536
rect 37464 34527 37516 34536
rect 37464 34493 37473 34527
rect 37473 34493 37507 34527
rect 37507 34493 37516 34527
rect 37464 34484 37516 34493
rect 1676 34391 1728 34400
rect 1676 34357 1685 34391
rect 1685 34357 1719 34391
rect 1719 34357 1728 34391
rect 1676 34348 1728 34357
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 1584 32376 1636 32428
rect 25504 32419 25556 32428
rect 25504 32385 25513 32419
rect 25513 32385 25547 32419
rect 25547 32385 25556 32419
rect 25504 32376 25556 32385
rect 38292 32351 38344 32360
rect 38292 32317 38301 32351
rect 38301 32317 38335 32351
rect 38335 32317 38344 32351
rect 38292 32308 38344 32317
rect 2688 32240 2740 32292
rect 8024 32172 8076 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1584 32011 1636 32020
rect 1584 31977 1593 32011
rect 1593 31977 1627 32011
rect 1627 31977 1636 32011
rect 1584 31968 1636 31977
rect 38292 32011 38344 32020
rect 38292 31977 38301 32011
rect 38301 31977 38335 32011
rect 38335 31977 38344 32011
rect 38292 31968 38344 31977
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 23848 31467 23900 31476
rect 23848 31433 23857 31467
rect 23857 31433 23891 31467
rect 23891 31433 23900 31467
rect 23848 31424 23900 31433
rect 24308 31288 24360 31340
rect 25504 31331 25556 31340
rect 25504 31297 25513 31331
rect 25513 31297 25547 31331
rect 25547 31297 25556 31331
rect 25504 31288 25556 31297
rect 24308 31127 24360 31136
rect 24308 31093 24317 31127
rect 24317 31093 24351 31127
rect 24351 31093 24360 31127
rect 24308 31084 24360 31093
rect 25136 31084 25188 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 9312 30676 9364 30728
rect 23388 30676 23440 30728
rect 33692 30608 33744 30660
rect 1676 30583 1728 30592
rect 1676 30549 1685 30583
rect 1685 30549 1719 30583
rect 1719 30549 1728 30583
rect 1676 30540 1728 30549
rect 2320 30583 2372 30592
rect 2320 30549 2329 30583
rect 2329 30549 2363 30583
rect 2363 30549 2372 30583
rect 2320 30540 2372 30549
rect 22928 30540 22980 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 17684 30200 17736 30252
rect 25780 30132 25832 30184
rect 38292 30175 38344 30184
rect 38292 30141 38301 30175
rect 38301 30141 38335 30175
rect 38335 30141 38344 30175
rect 38292 30132 38344 30141
rect 20076 29996 20128 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 38292 29835 38344 29844
rect 38292 29801 38301 29835
rect 38301 29801 38335 29835
rect 38335 29801 38344 29835
rect 38292 29792 38344 29801
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 14280 29248 14332 29300
rect 1860 29155 1912 29164
rect 1860 29121 1869 29155
rect 1869 29121 1903 29155
rect 1903 29121 1912 29155
rect 1860 29112 1912 29121
rect 22744 29155 22796 29164
rect 1676 29019 1728 29028
rect 1676 28985 1685 29019
rect 1685 28985 1719 29019
rect 1719 28985 1728 29019
rect 1676 28976 1728 28985
rect 22744 29121 22753 29155
rect 22753 29121 22787 29155
rect 22787 29121 22796 29155
rect 22744 29112 22796 29121
rect 38016 29155 38068 29164
rect 38016 29121 38025 29155
rect 38025 29121 38059 29155
rect 38059 29121 38068 29155
rect 38016 29112 38068 29121
rect 16580 28976 16632 29028
rect 23204 28976 23256 29028
rect 38200 29019 38252 29028
rect 38200 28985 38209 29019
rect 38209 28985 38243 29019
rect 38243 28985 38252 29019
rect 38200 28976 38252 28985
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2228 28500 2280 28552
rect 23112 28500 23164 28552
rect 38016 28364 38068 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 2688 27820 2740 27872
rect 24032 28160 24084 28212
rect 26056 28160 26108 28212
rect 22468 27863 22520 27872
rect 22468 27829 22477 27863
rect 22477 27829 22511 27863
rect 22511 27829 22520 27863
rect 22468 27820 22520 27829
rect 25688 27820 25740 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 1584 26911 1636 26920
rect 1584 26877 1593 26911
rect 1593 26877 1627 26911
rect 1627 26877 1636 26911
rect 1584 26868 1636 26877
rect 2228 26868 2280 26920
rect 38016 26911 38068 26920
rect 38016 26877 38025 26911
rect 38025 26877 38059 26911
rect 38059 26877 38068 26911
rect 38016 26868 38068 26877
rect 38292 26911 38344 26920
rect 38292 26877 38301 26911
rect 38301 26877 38335 26911
rect 38335 26877 38344 26911
rect 38292 26868 38344 26877
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 1584 26571 1636 26580
rect 1584 26537 1593 26571
rect 1593 26537 1627 26571
rect 1627 26537 1636 26571
rect 1584 26528 1636 26537
rect 23112 26571 23164 26580
rect 23112 26537 23121 26571
rect 23121 26537 23155 26571
rect 23155 26537 23164 26571
rect 23112 26528 23164 26537
rect 38292 26571 38344 26580
rect 38292 26537 38301 26571
rect 38301 26537 38335 26571
rect 38335 26537 38344 26571
rect 38292 26528 38344 26537
rect 1860 26392 1912 26444
rect 24124 26392 24176 26444
rect 23112 26324 23164 26376
rect 22652 26256 22704 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 2044 24760 2096 24812
rect 38200 24803 38252 24812
rect 38200 24769 38209 24803
rect 38209 24769 38243 24803
rect 38243 24769 38252 24803
rect 38200 24760 38252 24769
rect 1676 24599 1728 24608
rect 1676 24565 1685 24599
rect 1685 24565 1719 24599
rect 1719 24565 1728 24599
rect 1676 24556 1728 24565
rect 24124 24556 24176 24608
rect 24768 24556 24820 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 25780 24395 25832 24404
rect 25780 24361 25789 24395
rect 25789 24361 25823 24395
rect 25823 24361 25832 24395
rect 25780 24352 25832 24361
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4804 23808 4856 23860
rect 28724 23851 28776 23860
rect 28724 23817 28733 23851
rect 28733 23817 28767 23851
rect 28767 23817 28776 23851
rect 28724 23808 28776 23817
rect 24216 23740 24268 23792
rect 37464 23808 37516 23860
rect 22468 23672 22520 23724
rect 23296 23672 23348 23724
rect 22560 23647 22612 23656
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 25780 23672 25832 23724
rect 26332 23715 26384 23724
rect 26332 23681 26341 23715
rect 26341 23681 26375 23715
rect 26375 23681 26384 23715
rect 26332 23672 26384 23681
rect 28080 23672 28132 23724
rect 7472 23536 7524 23588
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 5540 23264 5592 23316
rect 23296 23307 23348 23316
rect 23296 23273 23305 23307
rect 23305 23273 23339 23307
rect 23339 23273 23348 23307
rect 23296 23264 23348 23273
rect 25780 23264 25832 23316
rect 22652 23171 22704 23180
rect 22652 23137 22661 23171
rect 22661 23137 22695 23171
rect 22695 23137 22704 23171
rect 22652 23128 22704 23137
rect 22836 23103 22888 23112
rect 1676 22967 1728 22976
rect 1676 22933 1685 22967
rect 1685 22933 1719 22967
rect 1719 22933 1728 22967
rect 1676 22924 1728 22933
rect 22836 23069 22845 23103
rect 22845 23069 22879 23103
rect 22879 23069 22888 23103
rect 22836 23060 22888 23069
rect 25780 23060 25832 23112
rect 12072 22924 12124 22976
rect 25504 22924 25556 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 25412 22695 25464 22704
rect 25412 22661 25421 22695
rect 25421 22661 25455 22695
rect 25455 22661 25464 22695
rect 25412 22652 25464 22661
rect 25504 22695 25556 22704
rect 25504 22661 25513 22695
rect 25513 22661 25547 22695
rect 25547 22661 25556 22695
rect 25504 22652 25556 22661
rect 1676 22627 1728 22636
rect 1676 22593 1685 22627
rect 1685 22593 1719 22627
rect 1719 22593 1728 22627
rect 1676 22584 1728 22593
rect 35716 22584 35768 22636
rect 23020 22559 23072 22568
rect 23020 22525 23029 22559
rect 23029 22525 23063 22559
rect 23063 22525 23072 22559
rect 23020 22516 23072 22525
rect 1860 22491 1912 22500
rect 1860 22457 1869 22491
rect 1869 22457 1903 22491
rect 1903 22457 1912 22491
rect 1860 22448 1912 22457
rect 24952 22491 25004 22500
rect 24952 22457 24961 22491
rect 24961 22457 24995 22491
rect 24995 22457 25004 22491
rect 24952 22448 25004 22457
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 22836 22176 22888 22228
rect 23296 22219 23348 22228
rect 23296 22185 23305 22219
rect 23305 22185 23339 22219
rect 23339 22185 23348 22219
rect 23296 22176 23348 22185
rect 25412 22176 25464 22228
rect 23020 22040 23072 22092
rect 2044 21879 2096 21888
rect 2044 21845 2053 21879
rect 2053 21845 2087 21879
rect 2087 21845 2096 21879
rect 2044 21836 2096 21845
rect 22284 22015 22336 22024
rect 22284 21981 22293 22015
rect 22293 21981 22327 22015
rect 22327 21981 22336 22015
rect 22284 21972 22336 21981
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 24032 21972 24084 22024
rect 10140 21836 10192 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 22560 21632 22612 21684
rect 23112 21675 23164 21684
rect 23112 21641 23121 21675
rect 23121 21641 23155 21675
rect 23155 21641 23164 21675
rect 23112 21632 23164 21641
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 22744 21496 22796 21548
rect 24032 21496 24084 21548
rect 24584 21292 24636 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 24492 20884 24544 20936
rect 1584 20816 1636 20868
rect 16580 20816 16632 20868
rect 19984 20816 20036 20868
rect 2320 20748 2372 20800
rect 22744 20791 22796 20800
rect 22744 20757 22753 20791
rect 22753 20757 22787 20791
rect 22787 20757 22796 20791
rect 22744 20748 22796 20757
rect 23388 20791 23440 20800
rect 23388 20757 23397 20791
rect 23397 20757 23431 20791
rect 23431 20757 23440 20791
rect 23388 20748 23440 20757
rect 24032 20791 24084 20800
rect 24032 20757 24041 20791
rect 24041 20757 24075 20791
rect 24075 20757 24084 20791
rect 24032 20748 24084 20757
rect 24400 20748 24452 20800
rect 38200 20791 38252 20800
rect 38200 20757 38209 20791
rect 38209 20757 38243 20791
rect 38243 20757 38252 20791
rect 38200 20748 38252 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1584 20519 1636 20528
rect 1584 20485 1593 20519
rect 1593 20485 1627 20519
rect 1627 20485 1636 20519
rect 1584 20476 1636 20485
rect 1860 20204 1912 20256
rect 24308 20544 24360 20596
rect 37924 20544 37976 20596
rect 23664 20476 23716 20528
rect 25320 20519 25372 20528
rect 25320 20485 25329 20519
rect 25329 20485 25363 20519
rect 25363 20485 25372 20519
rect 25320 20476 25372 20485
rect 37832 20451 37884 20460
rect 23388 20383 23440 20392
rect 23388 20349 23397 20383
rect 23397 20349 23431 20383
rect 23431 20349 23440 20383
rect 23388 20340 23440 20349
rect 24952 20383 25004 20392
rect 24952 20349 24961 20383
rect 24961 20349 24995 20383
rect 24995 20349 25004 20383
rect 24952 20340 25004 20349
rect 25228 20340 25280 20392
rect 23756 20204 23808 20256
rect 26424 20204 26476 20256
rect 37832 20417 37841 20451
rect 37841 20417 37875 20451
rect 37875 20417 37884 20451
rect 37832 20408 37884 20417
rect 28080 20204 28132 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 23664 20043 23716 20052
rect 23664 20009 23673 20043
rect 23673 20009 23707 20043
rect 23707 20009 23716 20043
rect 23664 20000 23716 20009
rect 25320 20000 25372 20052
rect 2136 19932 2188 19984
rect 22284 19864 22336 19916
rect 16580 19839 16632 19848
rect 16580 19805 16589 19839
rect 16589 19805 16623 19839
rect 16623 19805 16632 19839
rect 16580 19796 16632 19805
rect 22468 19839 22520 19848
rect 22468 19805 22477 19839
rect 22477 19805 22511 19839
rect 22511 19805 22520 19839
rect 22468 19796 22520 19805
rect 23296 19796 23348 19848
rect 23664 19796 23716 19848
rect 19248 19728 19300 19780
rect 22744 19728 22796 19780
rect 9864 19703 9916 19712
rect 9864 19669 9873 19703
rect 9873 19669 9907 19703
rect 9907 19669 9916 19703
rect 9864 19660 9916 19669
rect 23480 19660 23532 19712
rect 25504 19660 25556 19712
rect 37280 19660 37332 19712
rect 37832 19660 37884 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 23296 19499 23348 19508
rect 23296 19465 23305 19499
rect 23305 19465 23339 19499
rect 23339 19465 23348 19499
rect 23296 19456 23348 19465
rect 22192 19431 22244 19440
rect 22192 19397 22201 19431
rect 22201 19397 22235 19431
rect 22235 19397 22244 19431
rect 22192 19388 22244 19397
rect 24216 19431 24268 19440
rect 24216 19397 24225 19431
rect 24225 19397 24259 19431
rect 24259 19397 24268 19431
rect 24216 19388 24268 19397
rect 26884 19456 26936 19508
rect 25228 19431 25280 19440
rect 25228 19397 25237 19431
rect 25237 19397 25271 19431
rect 25271 19397 25280 19431
rect 26332 19431 26384 19440
rect 25228 19388 25280 19397
rect 26332 19397 26341 19431
rect 26341 19397 26375 19431
rect 26375 19397 26384 19431
rect 26332 19388 26384 19397
rect 26424 19431 26476 19440
rect 26424 19397 26433 19431
rect 26433 19397 26467 19431
rect 26467 19397 26476 19431
rect 26424 19388 26476 19397
rect 15752 19320 15804 19372
rect 20076 19320 20128 19372
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 23664 19320 23716 19372
rect 33140 19320 33192 19372
rect 22284 19184 22336 19236
rect 25412 19184 25464 19236
rect 38200 19159 38252 19168
rect 38200 19125 38209 19159
rect 38209 19125 38243 19159
rect 38243 19125 38252 19159
rect 38200 19116 38252 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 26332 18912 26384 18964
rect 37740 18912 37792 18964
rect 22468 18844 22520 18896
rect 22560 18844 22612 18896
rect 19248 18776 19300 18828
rect 22284 18819 22336 18828
rect 22284 18785 22293 18819
rect 22293 18785 22327 18819
rect 22327 18785 22336 18819
rect 22284 18776 22336 18785
rect 22928 18776 22980 18828
rect 23204 18776 23256 18828
rect 2228 18708 2280 18760
rect 25504 18708 25556 18760
rect 38108 18708 38160 18760
rect 21732 18683 21784 18692
rect 21732 18649 21741 18683
rect 21741 18649 21775 18683
rect 21775 18649 21784 18683
rect 21732 18640 21784 18649
rect 22652 18572 22704 18624
rect 24768 18572 24820 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 25412 18343 25464 18352
rect 25412 18309 25421 18343
rect 25421 18309 25455 18343
rect 25455 18309 25464 18343
rect 25412 18300 25464 18309
rect 26332 18300 26384 18352
rect 26516 18300 26568 18352
rect 22100 18232 22152 18284
rect 23756 18275 23808 18284
rect 23756 18241 23765 18275
rect 23765 18241 23799 18275
rect 23799 18241 23808 18275
rect 23756 18232 23808 18241
rect 24768 18232 24820 18284
rect 22652 18207 22704 18216
rect 22652 18173 22661 18207
rect 22661 18173 22695 18207
rect 22695 18173 22704 18207
rect 22652 18164 22704 18173
rect 23112 18207 23164 18216
rect 23112 18173 23121 18207
rect 23121 18173 23155 18207
rect 23155 18173 23164 18207
rect 23112 18164 23164 18173
rect 23480 18096 23532 18148
rect 22100 18071 22152 18080
rect 22100 18037 22109 18071
rect 22109 18037 22143 18071
rect 22143 18037 22152 18071
rect 27160 18071 27212 18080
rect 22100 18028 22152 18037
rect 27160 18037 27169 18071
rect 27169 18037 27203 18071
rect 27203 18037 27212 18071
rect 27160 18028 27212 18037
rect 38108 18071 38160 18080
rect 38108 18037 38117 18071
rect 38117 18037 38151 18071
rect 38151 18037 38160 18071
rect 38108 18028 38160 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 21732 17867 21784 17876
rect 21732 17833 21741 17867
rect 21741 17833 21775 17867
rect 21775 17833 21784 17867
rect 21732 17824 21784 17833
rect 22192 17824 22244 17876
rect 26332 17824 26384 17876
rect 33140 17824 33192 17876
rect 26884 17799 26936 17808
rect 26884 17765 26893 17799
rect 26893 17765 26927 17799
rect 26927 17765 26936 17799
rect 26884 17756 26936 17765
rect 22100 17688 22152 17740
rect 23480 17688 23532 17740
rect 24216 17688 24268 17740
rect 25688 17731 25740 17740
rect 25688 17697 25697 17731
rect 25697 17697 25731 17731
rect 25731 17697 25740 17731
rect 25688 17688 25740 17697
rect 26700 17688 26752 17740
rect 22744 17620 22796 17672
rect 24768 17663 24820 17672
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 22652 17484 22704 17536
rect 23296 17552 23348 17604
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 25872 17663 25924 17672
rect 25872 17629 25881 17663
rect 25881 17629 25915 17663
rect 25915 17629 25924 17663
rect 25872 17620 25924 17629
rect 26608 17620 26660 17672
rect 27160 17620 27212 17672
rect 26240 17484 26292 17536
rect 31208 17484 31260 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 23112 17280 23164 17332
rect 24768 17280 24820 17332
rect 25872 17280 25924 17332
rect 6828 17144 6880 17196
rect 22744 17144 22796 17196
rect 24400 17144 24452 17196
rect 26516 17212 26568 17264
rect 27436 17144 27488 17196
rect 27528 17144 27580 17196
rect 38292 17187 38344 17196
rect 38292 17153 38301 17187
rect 38301 17153 38335 17187
rect 38335 17153 38344 17187
rect 38292 17144 38344 17153
rect 23388 17076 23440 17128
rect 26332 17076 26384 17128
rect 1676 17051 1728 17060
rect 1676 17017 1685 17051
rect 1685 17017 1719 17051
rect 1719 17017 1728 17051
rect 1676 17008 1728 17017
rect 23204 17008 23256 17060
rect 21180 16940 21232 16992
rect 24400 17008 24452 17060
rect 25044 16940 25096 16992
rect 37924 16940 37976 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2228 16736 2280 16788
rect 10784 16643 10836 16652
rect 2228 16532 2280 16584
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 20076 16643 20128 16652
rect 20076 16609 20085 16643
rect 20085 16609 20119 16643
rect 20119 16609 20128 16643
rect 20076 16600 20128 16609
rect 23296 16736 23348 16788
rect 25320 16736 25372 16788
rect 34796 16736 34848 16788
rect 23112 16711 23164 16720
rect 23112 16677 23121 16711
rect 23121 16677 23155 16711
rect 23155 16677 23164 16711
rect 23112 16668 23164 16677
rect 10140 16532 10192 16541
rect 21180 16575 21232 16584
rect 21180 16541 21189 16575
rect 21189 16541 21223 16575
rect 21223 16541 21232 16575
rect 21180 16532 21232 16541
rect 23572 16532 23624 16584
rect 25044 16600 25096 16652
rect 26516 16600 26568 16652
rect 26976 16575 27028 16584
rect 20260 16507 20312 16516
rect 20260 16473 20269 16507
rect 20269 16473 20303 16507
rect 20303 16473 20312 16507
rect 20260 16464 20312 16473
rect 22560 16507 22612 16516
rect 1768 16439 1820 16448
rect 1768 16405 1777 16439
rect 1777 16405 1811 16439
rect 1811 16405 1820 16439
rect 1768 16396 1820 16405
rect 21824 16439 21876 16448
rect 21824 16405 21833 16439
rect 21833 16405 21867 16439
rect 21867 16405 21876 16439
rect 21824 16396 21876 16405
rect 22560 16473 22569 16507
rect 22569 16473 22603 16507
rect 22603 16473 22612 16507
rect 22560 16464 22612 16473
rect 23480 16464 23532 16516
rect 26976 16541 26985 16575
rect 26985 16541 27019 16575
rect 27019 16541 27028 16575
rect 26976 16532 27028 16541
rect 27160 16532 27212 16584
rect 27528 16532 27580 16584
rect 25320 16464 25372 16516
rect 27344 16464 27396 16516
rect 24768 16396 24820 16448
rect 24860 16396 24912 16448
rect 27528 16439 27580 16448
rect 27528 16405 27537 16439
rect 27537 16405 27571 16439
rect 27571 16405 27580 16439
rect 27528 16396 27580 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 22652 16192 22704 16244
rect 20260 16124 20312 16176
rect 37832 16192 37884 16244
rect 21456 16099 21508 16108
rect 21456 16065 21465 16099
rect 21465 16065 21499 16099
rect 21499 16065 21508 16099
rect 21456 16056 21508 16065
rect 23480 16124 23532 16176
rect 23940 16124 23992 16176
rect 27068 16124 27120 16176
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 24768 16099 24820 16108
rect 24768 16065 24777 16099
rect 24777 16065 24811 16099
rect 24811 16065 24820 16099
rect 24768 16056 24820 16065
rect 26700 16056 26752 16108
rect 27160 16099 27212 16108
rect 27160 16065 27169 16099
rect 27169 16065 27203 16099
rect 27203 16065 27212 16099
rect 27160 16056 27212 16065
rect 23756 15988 23808 16040
rect 23848 15920 23900 15972
rect 24032 15963 24084 15972
rect 24032 15929 24041 15963
rect 24041 15929 24075 15963
rect 24075 15929 24084 15963
rect 24032 15920 24084 15929
rect 26240 15988 26292 16040
rect 25688 15852 25740 15904
rect 27252 15895 27304 15904
rect 27252 15861 27261 15895
rect 27261 15861 27295 15895
rect 27295 15861 27304 15895
rect 27252 15852 27304 15861
rect 27896 15895 27948 15904
rect 27896 15861 27905 15895
rect 27905 15861 27939 15895
rect 27939 15861 27948 15895
rect 27896 15852 27948 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 6828 15648 6880 15700
rect 22560 15648 22612 15700
rect 21456 15580 21508 15632
rect 23020 15580 23072 15632
rect 26240 15580 26292 15632
rect 27436 15648 27488 15700
rect 29368 15580 29420 15632
rect 23112 15555 23164 15564
rect 23112 15521 23121 15555
rect 23121 15521 23155 15555
rect 23155 15521 23164 15555
rect 23112 15512 23164 15521
rect 24584 15555 24636 15564
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 24860 15512 24912 15564
rect 25688 15555 25740 15564
rect 25688 15521 25697 15555
rect 25697 15521 25731 15555
rect 25731 15521 25740 15555
rect 25688 15512 25740 15521
rect 27528 15512 27580 15564
rect 1676 15351 1728 15360
rect 1676 15317 1685 15351
rect 1685 15317 1719 15351
rect 1719 15317 1728 15351
rect 1676 15308 1728 15317
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 26332 15487 26384 15496
rect 22192 15444 22244 15453
rect 19156 15376 19208 15428
rect 12164 15308 12216 15360
rect 26332 15453 26341 15487
rect 26341 15453 26375 15487
rect 26375 15453 26384 15487
rect 26332 15444 26384 15453
rect 27896 15512 27948 15564
rect 30472 15512 30524 15564
rect 38016 15487 38068 15496
rect 22836 15419 22888 15428
rect 22836 15385 22845 15419
rect 22845 15385 22879 15419
rect 22879 15385 22888 15419
rect 22836 15376 22888 15385
rect 22928 15419 22980 15428
rect 22928 15385 22937 15419
rect 22937 15385 22971 15419
rect 22971 15385 22980 15419
rect 22928 15376 22980 15385
rect 25872 15376 25924 15428
rect 38016 15453 38025 15487
rect 38025 15453 38059 15487
rect 38059 15453 38068 15487
rect 38016 15444 38068 15453
rect 37280 15376 37332 15428
rect 23204 15308 23256 15360
rect 26332 15308 26384 15360
rect 28172 15351 28224 15360
rect 28172 15317 28181 15351
rect 28181 15317 28215 15351
rect 28215 15317 28224 15351
rect 28172 15308 28224 15317
rect 38200 15351 38252 15360
rect 38200 15317 38209 15351
rect 38209 15317 38243 15351
rect 38243 15317 38252 15351
rect 38200 15308 38252 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 12164 15147 12216 15156
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 22928 15104 22980 15156
rect 23572 15104 23624 15156
rect 23848 15104 23900 15156
rect 27344 15104 27396 15156
rect 23480 15079 23532 15088
rect 23480 15045 23489 15079
rect 23489 15045 23523 15079
rect 23523 15045 23532 15079
rect 23480 15036 23532 15045
rect 24032 15079 24084 15088
rect 24032 15045 24041 15079
rect 24041 15045 24075 15079
rect 24075 15045 24084 15079
rect 24032 15036 24084 15045
rect 24584 15079 24636 15088
rect 24584 15045 24593 15079
rect 24593 15045 24627 15079
rect 24627 15045 24636 15079
rect 24584 15036 24636 15045
rect 22560 14968 22612 15020
rect 25596 14968 25648 15020
rect 25872 15011 25924 15020
rect 25872 14977 25881 15011
rect 25881 14977 25915 15011
rect 25915 14977 25924 15011
rect 25872 14968 25924 14977
rect 26240 14968 26292 15020
rect 27252 14968 27304 15020
rect 28540 14968 28592 15020
rect 23388 14943 23440 14952
rect 23388 14909 23397 14943
rect 23397 14909 23431 14943
rect 23431 14909 23440 14943
rect 23388 14900 23440 14909
rect 26424 14900 26476 14952
rect 27620 14900 27672 14952
rect 28172 14900 28224 14952
rect 22192 14832 22244 14884
rect 27712 14807 27764 14816
rect 27712 14773 27721 14807
rect 27721 14773 27755 14807
rect 27755 14773 27764 14807
rect 27712 14764 27764 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1860 14560 1912 14612
rect 35716 14603 35768 14612
rect 35716 14569 35725 14603
rect 35725 14569 35759 14603
rect 35759 14569 35768 14603
rect 35716 14560 35768 14569
rect 22100 14467 22152 14476
rect 22100 14433 22109 14467
rect 22109 14433 22143 14467
rect 22143 14433 22152 14467
rect 22100 14424 22152 14433
rect 23112 14424 23164 14476
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 23388 14399 23440 14408
rect 23388 14365 23397 14399
rect 23397 14365 23431 14399
rect 23431 14365 23440 14399
rect 23388 14356 23440 14365
rect 23572 14399 23624 14408
rect 23572 14365 23581 14399
rect 23581 14365 23615 14399
rect 23615 14365 23624 14399
rect 23572 14356 23624 14365
rect 27712 14492 27764 14544
rect 26332 14424 26384 14476
rect 26424 14467 26476 14476
rect 26424 14433 26433 14467
rect 26433 14433 26467 14467
rect 26467 14433 26476 14467
rect 26424 14424 26476 14433
rect 27620 14424 27672 14476
rect 25136 14356 25188 14408
rect 35348 14356 35400 14408
rect 1952 14288 2004 14340
rect 22192 14331 22244 14340
rect 22192 14297 22201 14331
rect 22201 14297 22235 14331
rect 22235 14297 22244 14331
rect 26700 14331 26752 14340
rect 22192 14288 22244 14297
rect 26700 14297 26709 14331
rect 26709 14297 26743 14331
rect 26743 14297 26752 14331
rect 26700 14288 26752 14297
rect 26792 14288 26844 14340
rect 27896 14331 27948 14340
rect 27896 14297 27905 14331
rect 27905 14297 27939 14331
rect 27939 14297 27948 14331
rect 27896 14288 27948 14297
rect 22652 14220 22704 14272
rect 22836 14220 22888 14272
rect 23664 14220 23716 14272
rect 26976 14220 27028 14272
rect 37740 14220 37792 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 22192 14059 22244 14068
rect 22192 14025 22201 14059
rect 22201 14025 22235 14059
rect 22235 14025 22244 14059
rect 22192 14016 22244 14025
rect 23572 14016 23624 14068
rect 23940 14059 23992 14068
rect 23940 14025 23949 14059
rect 23949 14025 23983 14059
rect 23983 14025 23992 14059
rect 23940 14016 23992 14025
rect 26332 14016 26384 14068
rect 27068 14016 27120 14068
rect 38016 14059 38068 14068
rect 38016 14025 38025 14059
rect 38025 14025 38059 14059
rect 38059 14025 38068 14059
rect 38016 14016 38068 14025
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 25688 13948 25740 14000
rect 28448 13948 28500 14000
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 21180 13880 21232 13932
rect 23204 13880 23256 13932
rect 23664 13880 23716 13932
rect 22376 13812 22428 13864
rect 26792 13880 26844 13932
rect 27528 13880 27580 13932
rect 37740 13880 37792 13932
rect 24492 13855 24544 13864
rect 24492 13821 24501 13855
rect 24501 13821 24535 13855
rect 24535 13821 24544 13855
rect 24492 13812 24544 13821
rect 26240 13812 26292 13864
rect 22836 13676 22888 13728
rect 26884 13676 26936 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 23480 13472 23532 13524
rect 25688 13472 25740 13524
rect 26700 13472 26752 13524
rect 24308 13404 24360 13456
rect 24492 13404 24544 13456
rect 22376 13379 22428 13388
rect 22376 13345 22385 13379
rect 22385 13345 22419 13379
rect 22419 13345 22428 13379
rect 22376 13336 22428 13345
rect 23388 13336 23440 13388
rect 4620 13268 4672 13320
rect 1952 13200 2004 13252
rect 1676 13175 1728 13184
rect 1676 13141 1685 13175
rect 1685 13141 1719 13175
rect 1719 13141 1728 13175
rect 1676 13132 1728 13141
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 20904 13132 20956 13184
rect 25780 13311 25832 13320
rect 25780 13277 25789 13311
rect 25789 13277 25823 13311
rect 25823 13277 25832 13311
rect 25780 13268 25832 13277
rect 25964 13311 26016 13320
rect 25964 13277 25973 13311
rect 25973 13277 26007 13311
rect 26007 13277 26016 13311
rect 25964 13268 26016 13277
rect 27252 13268 27304 13320
rect 38016 13311 38068 13320
rect 38016 13277 38025 13311
rect 38025 13277 38059 13311
rect 38059 13277 38068 13311
rect 38016 13268 38068 13277
rect 24584 13243 24636 13252
rect 24584 13209 24593 13243
rect 24593 13209 24627 13243
rect 24627 13209 24636 13243
rect 24584 13200 24636 13209
rect 24768 13200 24820 13252
rect 25228 13243 25280 13252
rect 25228 13209 25237 13243
rect 25237 13209 25271 13243
rect 25271 13209 25280 13243
rect 25228 13200 25280 13209
rect 25872 13132 25924 13184
rect 38200 13175 38252 13184
rect 38200 13141 38209 13175
rect 38209 13141 38243 13175
rect 38243 13141 38252 13175
rect 38200 13132 38252 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 10600 12928 10652 12980
rect 22100 12928 22152 12980
rect 25964 12928 26016 12980
rect 26332 12971 26384 12980
rect 26332 12937 26341 12971
rect 26341 12937 26375 12971
rect 26375 12937 26384 12971
rect 26332 12928 26384 12937
rect 27896 12971 27948 12980
rect 20812 12903 20864 12912
rect 20812 12869 20821 12903
rect 20821 12869 20855 12903
rect 20855 12869 20864 12903
rect 20812 12860 20864 12869
rect 23756 12903 23808 12912
rect 23756 12869 23765 12903
rect 23765 12869 23799 12903
rect 23799 12869 23808 12903
rect 23756 12860 23808 12869
rect 24032 12860 24084 12912
rect 27896 12937 27905 12971
rect 27905 12937 27939 12971
rect 27939 12937 27948 12971
rect 27896 12928 27948 12937
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 22284 12724 22336 12776
rect 22836 12792 22888 12844
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 22100 12588 22152 12640
rect 22928 12724 22980 12776
rect 27252 12792 27304 12844
rect 29184 12860 29236 12912
rect 27896 12724 27948 12776
rect 25228 12656 25280 12708
rect 26516 12656 26568 12708
rect 27620 12588 27672 12640
rect 37740 12588 37792 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 4620 12384 4672 12436
rect 20812 12384 20864 12436
rect 22284 12384 22336 12436
rect 28448 12427 28500 12436
rect 2504 12248 2556 12300
rect 20720 12248 20772 12300
rect 22284 12291 22336 12300
rect 22284 12257 22293 12291
rect 22293 12257 22327 12291
rect 22327 12257 22336 12291
rect 22284 12248 22336 12257
rect 23112 12316 23164 12368
rect 23296 12316 23348 12368
rect 24952 12291 25004 12300
rect 24952 12257 24961 12291
rect 24961 12257 24995 12291
rect 24995 12257 25004 12291
rect 24952 12248 25004 12257
rect 28448 12393 28457 12427
rect 28457 12393 28491 12427
rect 28491 12393 28500 12427
rect 28448 12384 28500 12393
rect 27620 12248 27672 12300
rect 15752 12180 15804 12232
rect 16396 12180 16448 12232
rect 20812 12180 20864 12232
rect 27896 12223 27948 12232
rect 27896 12189 27905 12223
rect 27905 12189 27939 12223
rect 27939 12189 27948 12223
rect 27896 12180 27948 12189
rect 29460 12180 29512 12232
rect 22376 12112 22428 12164
rect 4988 12087 5040 12096
rect 4988 12053 4997 12087
rect 4997 12053 5031 12087
rect 5031 12053 5040 12087
rect 4988 12044 5040 12053
rect 22652 12044 22704 12096
rect 23296 12155 23348 12164
rect 23296 12121 23305 12155
rect 23305 12121 23339 12155
rect 23339 12121 23348 12155
rect 23296 12112 23348 12121
rect 24124 12112 24176 12164
rect 24584 12112 24636 12164
rect 25688 12112 25740 12164
rect 29092 12112 29144 12164
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 22100 11840 22152 11892
rect 25780 11840 25832 11892
rect 26516 11840 26568 11892
rect 22192 11815 22244 11824
rect 22192 11781 22201 11815
rect 22201 11781 22235 11815
rect 22235 11781 22244 11815
rect 22192 11772 22244 11781
rect 23020 11772 23072 11824
rect 24032 11772 24084 11824
rect 24584 11815 24636 11824
rect 24584 11781 24593 11815
rect 24593 11781 24627 11815
rect 24627 11781 24636 11815
rect 24584 11772 24636 11781
rect 25872 11772 25924 11824
rect 24860 11679 24912 11688
rect 19984 11568 20036 11620
rect 21180 11500 21232 11552
rect 21548 11568 21600 11620
rect 24860 11645 24869 11679
rect 24869 11645 24903 11679
rect 24903 11645 24912 11679
rect 24860 11636 24912 11645
rect 25136 11636 25188 11688
rect 27068 11704 27120 11756
rect 27436 11704 27488 11756
rect 22652 11568 22704 11620
rect 22928 11568 22980 11620
rect 26700 11568 26752 11620
rect 38016 11568 38068 11620
rect 26792 11500 26844 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 4988 11296 5040 11348
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 22376 11339 22428 11348
rect 22376 11305 22385 11339
rect 22385 11305 22419 11339
rect 22419 11305 22428 11339
rect 22376 11296 22428 11305
rect 23020 11339 23072 11348
rect 23020 11305 23029 11339
rect 23029 11305 23063 11339
rect 23063 11305 23072 11339
rect 23020 11296 23072 11305
rect 23756 11296 23808 11348
rect 24860 11228 24912 11280
rect 24952 11203 25004 11212
rect 24952 11169 24961 11203
rect 24961 11169 24995 11203
rect 24995 11169 25004 11203
rect 24952 11160 25004 11169
rect 26424 11203 26476 11212
rect 26424 11169 26433 11203
rect 26433 11169 26467 11203
rect 26467 11169 26476 11203
rect 26424 11160 26476 11169
rect 26792 11160 26844 11212
rect 1768 11092 1820 11144
rect 16396 11092 16448 11144
rect 21548 11135 21600 11144
rect 21548 11101 21557 11135
rect 21557 11101 21591 11135
rect 21591 11101 21600 11135
rect 21548 11092 21600 11101
rect 22100 11092 22152 11144
rect 23480 11092 23532 11144
rect 24216 11092 24268 11144
rect 27068 11092 27120 11144
rect 31484 11092 31536 11144
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 21916 11024 21968 11076
rect 24308 11024 24360 11076
rect 24676 11067 24728 11076
rect 24676 11033 24685 11067
rect 24685 11033 24719 11067
rect 24719 11033 24728 11067
rect 24676 11024 24728 11033
rect 26700 11067 26752 11076
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 24492 10956 24544 11008
rect 26700 11033 26709 11067
rect 26709 11033 26743 11067
rect 26743 11033 26752 11067
rect 26700 11024 26752 11033
rect 26792 11067 26844 11076
rect 26792 11033 26801 11067
rect 26801 11033 26835 11067
rect 26835 11033 26844 11067
rect 26792 11024 26844 11033
rect 27436 11024 27488 11076
rect 38108 11024 38160 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 23296 10795 23348 10804
rect 23296 10761 23305 10795
rect 23305 10761 23339 10795
rect 23339 10761 23348 10795
rect 23296 10752 23348 10761
rect 24768 10752 24820 10804
rect 24860 10752 24912 10804
rect 25320 10752 25372 10804
rect 36268 10795 36320 10804
rect 2412 10684 2464 10736
rect 17224 10684 17276 10736
rect 21916 10684 21968 10736
rect 22192 10727 22244 10736
rect 22192 10693 22201 10727
rect 22201 10693 22235 10727
rect 22235 10693 22244 10727
rect 25412 10727 25464 10736
rect 22192 10684 22244 10693
rect 25412 10693 25421 10727
rect 25421 10693 25455 10727
rect 25455 10693 25464 10727
rect 25412 10684 25464 10693
rect 36268 10761 36277 10795
rect 36277 10761 36311 10795
rect 36311 10761 36320 10795
rect 36268 10752 36320 10761
rect 38292 10795 38344 10804
rect 38292 10761 38301 10795
rect 38301 10761 38335 10795
rect 38335 10761 38344 10795
rect 38292 10752 38344 10761
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 14280 10616 14332 10668
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 14372 10548 14424 10600
rect 22744 10616 22796 10668
rect 24216 10616 24268 10668
rect 22100 10548 22152 10600
rect 26424 10616 26476 10668
rect 29092 10659 29144 10668
rect 29092 10625 29101 10659
rect 29101 10625 29135 10659
rect 29135 10625 29144 10659
rect 29092 10616 29144 10625
rect 29552 10616 29604 10668
rect 36176 10659 36228 10668
rect 36176 10625 36185 10659
rect 36185 10625 36219 10659
rect 36219 10625 36228 10659
rect 36176 10616 36228 10625
rect 33600 10548 33652 10600
rect 26608 10480 26660 10532
rect 20812 10412 20864 10464
rect 27804 10412 27856 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 17224 10251 17276 10260
rect 17224 10217 17233 10251
rect 17233 10217 17267 10251
rect 17267 10217 17276 10251
rect 17224 10208 17276 10217
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 20812 10208 20864 10260
rect 33600 10251 33652 10260
rect 33600 10217 33609 10251
rect 33609 10217 33643 10251
rect 33643 10217 33652 10251
rect 33600 10208 33652 10217
rect 21548 10140 21600 10192
rect 24676 10072 24728 10124
rect 23480 10004 23532 10056
rect 27068 10140 27120 10192
rect 24952 10072 25004 10124
rect 26608 10115 26660 10124
rect 26608 10081 26617 10115
rect 26617 10081 26651 10115
rect 26651 10081 26660 10115
rect 26608 10072 26660 10081
rect 29092 10004 29144 10056
rect 36176 10004 36228 10056
rect 22284 9979 22336 9988
rect 22284 9945 22293 9979
rect 22293 9945 22327 9979
rect 22327 9945 22336 9979
rect 22284 9936 22336 9945
rect 22376 9979 22428 9988
rect 22376 9945 22385 9979
rect 22385 9945 22419 9979
rect 22419 9945 22428 9979
rect 26516 9979 26568 9988
rect 22376 9936 22428 9945
rect 26516 9945 26525 9979
rect 26525 9945 26559 9979
rect 26559 9945 26568 9979
rect 26516 9936 26568 9945
rect 24676 9911 24728 9920
rect 24676 9877 24685 9911
rect 24685 9877 24719 9911
rect 24719 9877 24728 9911
rect 24676 9868 24728 9877
rect 26240 9868 26292 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 22376 9664 22428 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 24676 9639 24728 9648
rect 24676 9605 24685 9639
rect 24685 9605 24719 9639
rect 24719 9605 24728 9639
rect 24676 9596 24728 9605
rect 25320 9639 25372 9648
rect 25320 9605 25329 9639
rect 25329 9605 25363 9639
rect 25363 9605 25372 9639
rect 25320 9596 25372 9605
rect 26240 9639 26292 9648
rect 26240 9605 26249 9639
rect 26249 9605 26283 9639
rect 26283 9605 26292 9639
rect 26240 9596 26292 9605
rect 22100 9528 22152 9580
rect 23296 9528 23348 9580
rect 24124 9503 24176 9512
rect 24124 9469 24133 9503
rect 24133 9469 24167 9503
rect 24167 9469 24176 9503
rect 24124 9460 24176 9469
rect 26332 9503 26384 9512
rect 26332 9469 26341 9503
rect 26341 9469 26375 9503
rect 26375 9469 26384 9503
rect 26332 9460 26384 9469
rect 25044 9392 25096 9444
rect 26792 9392 26844 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 22284 9120 22336 9172
rect 24492 9120 24544 9172
rect 25044 9163 25096 9172
rect 25044 9129 25053 9163
rect 25053 9129 25087 9163
rect 25087 9129 25096 9163
rect 25044 9120 25096 9129
rect 24124 8984 24176 9036
rect 20812 8959 20864 8968
rect 20812 8925 20821 8959
rect 20821 8925 20855 8959
rect 20855 8925 20864 8959
rect 20812 8916 20864 8925
rect 24860 8916 24912 8968
rect 37832 9120 37884 9172
rect 38108 9163 38160 9172
rect 38108 9129 38117 9163
rect 38117 9129 38151 9163
rect 38151 9129 38160 9163
rect 38108 9120 38160 9129
rect 25688 9095 25740 9104
rect 25688 9061 25697 9095
rect 25697 9061 25731 9095
rect 25731 9061 25740 9095
rect 25688 9052 25740 9061
rect 26332 8984 26384 9036
rect 28816 8916 28868 8968
rect 29368 8916 29420 8968
rect 21456 8891 21508 8900
rect 21456 8857 21465 8891
rect 21465 8857 21499 8891
rect 21499 8857 21508 8891
rect 21456 8848 21508 8857
rect 28540 8848 28592 8900
rect 30472 8848 30524 8900
rect 38200 8891 38252 8900
rect 38200 8857 38209 8891
rect 38209 8857 38243 8891
rect 38243 8857 38252 8891
rect 38200 8848 38252 8857
rect 22468 8780 22520 8832
rect 27252 8823 27304 8832
rect 27252 8789 27261 8823
rect 27261 8789 27295 8823
rect 27295 8789 27304 8823
rect 27252 8780 27304 8789
rect 29276 8780 29328 8832
rect 30932 8780 30984 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 25412 8619 25464 8628
rect 25412 8585 25421 8619
rect 25421 8585 25455 8619
rect 25455 8585 25464 8619
rect 25412 8576 25464 8585
rect 26516 8576 26568 8628
rect 27068 8576 27120 8628
rect 22192 8508 22244 8560
rect 23296 8508 23348 8560
rect 22744 8440 22796 8492
rect 22284 8372 22336 8424
rect 19248 8304 19300 8356
rect 20812 8304 20864 8356
rect 26056 8440 26108 8492
rect 28540 8508 28592 8560
rect 29092 8508 29144 8560
rect 29276 8483 29328 8492
rect 29276 8449 29285 8483
rect 29285 8449 29319 8483
rect 29319 8449 29328 8483
rect 29276 8440 29328 8449
rect 24860 8415 24912 8424
rect 24860 8381 24869 8415
rect 24869 8381 24903 8415
rect 24903 8381 24912 8415
rect 24860 8372 24912 8381
rect 28908 8372 28960 8424
rect 30932 8508 30984 8560
rect 30104 8440 30156 8492
rect 31208 8415 31260 8424
rect 31208 8381 31217 8415
rect 31217 8381 31251 8415
rect 31251 8381 31260 8415
rect 31208 8372 31260 8381
rect 27436 8304 27488 8356
rect 28816 8236 28868 8288
rect 30012 8236 30064 8288
rect 32128 8236 32180 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 23296 8032 23348 8084
rect 24584 8032 24636 8084
rect 26516 8032 26568 8084
rect 27528 7964 27580 8016
rect 29552 7964 29604 8016
rect 31208 8032 31260 8084
rect 31576 7964 31628 8016
rect 31668 7964 31720 8016
rect 21456 7939 21508 7948
rect 21456 7905 21465 7939
rect 21465 7905 21499 7939
rect 21499 7905 21508 7939
rect 21456 7896 21508 7905
rect 22652 7896 22704 7948
rect 14096 7828 14148 7880
rect 22284 7871 22336 7880
rect 22284 7837 22293 7871
rect 22293 7837 22327 7871
rect 22327 7837 22336 7871
rect 22284 7828 22336 7837
rect 30012 7896 30064 7948
rect 30748 7896 30800 7948
rect 37832 7896 37884 7948
rect 25688 7828 25740 7880
rect 27252 7871 27304 7880
rect 27252 7837 27261 7871
rect 27261 7837 27295 7871
rect 27295 7837 27304 7871
rect 27252 7828 27304 7837
rect 21364 7760 21416 7812
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 22376 7692 22428 7744
rect 24124 7692 24176 7744
rect 26516 7760 26568 7812
rect 27528 7760 27580 7812
rect 26608 7692 26660 7744
rect 27712 7735 27764 7744
rect 27712 7701 27721 7735
rect 27721 7701 27755 7735
rect 27755 7701 27764 7735
rect 27712 7692 27764 7701
rect 29276 7828 29328 7880
rect 33140 7828 33192 7880
rect 38292 7871 38344 7880
rect 38292 7837 38301 7871
rect 38301 7837 38335 7871
rect 38335 7837 38344 7871
rect 38292 7828 38344 7837
rect 29000 7760 29052 7812
rect 32036 7760 32088 7812
rect 29552 7692 29604 7744
rect 30196 7692 30248 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 14096 7531 14148 7540
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 21364 7531 21416 7540
rect 21364 7497 21373 7531
rect 21373 7497 21407 7531
rect 21407 7497 21416 7531
rect 21364 7488 21416 7497
rect 22468 7531 22520 7540
rect 22468 7497 22477 7531
rect 22477 7497 22511 7531
rect 22511 7497 22520 7531
rect 22468 7488 22520 7497
rect 22744 7488 22796 7540
rect 26148 7488 26200 7540
rect 33692 7531 33744 7540
rect 33692 7497 33701 7531
rect 33701 7497 33735 7531
rect 33735 7497 33744 7531
rect 33692 7488 33744 7497
rect 38292 7531 38344 7540
rect 38292 7497 38301 7531
rect 38301 7497 38335 7531
rect 38335 7497 38344 7531
rect 38292 7488 38344 7497
rect 22376 7420 22428 7472
rect 27252 7420 27304 7472
rect 27436 7420 27488 7472
rect 29000 7420 29052 7472
rect 30656 7463 30708 7472
rect 30656 7429 30665 7463
rect 30665 7429 30699 7463
rect 30699 7429 30708 7463
rect 30656 7420 30708 7429
rect 23940 7284 23992 7336
rect 24216 7284 24268 7336
rect 24492 7284 24544 7336
rect 25688 7284 25740 7336
rect 27988 7284 28040 7336
rect 25136 7148 25188 7200
rect 25780 7191 25832 7200
rect 25780 7157 25789 7191
rect 25789 7157 25823 7191
rect 25823 7157 25832 7191
rect 27712 7216 27764 7268
rect 28448 7284 28500 7336
rect 29000 7284 29052 7336
rect 30656 7284 30708 7336
rect 32220 7352 32272 7404
rect 33140 7395 33192 7404
rect 33140 7361 33149 7395
rect 33149 7361 33183 7395
rect 33183 7361 33192 7395
rect 33140 7352 33192 7361
rect 34060 7284 34112 7336
rect 25780 7148 25832 7157
rect 27804 7148 27856 7200
rect 29368 7148 29420 7200
rect 29644 7148 29696 7200
rect 30656 7148 30708 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 22744 6944 22796 6996
rect 25596 6944 25648 6996
rect 28816 6944 28868 6996
rect 28908 6944 28960 6996
rect 31668 6944 31720 6996
rect 20720 6808 20772 6860
rect 21456 6808 21508 6860
rect 22284 6851 22336 6860
rect 22284 6817 22293 6851
rect 22293 6817 22327 6851
rect 22327 6817 22336 6851
rect 22284 6808 22336 6817
rect 23296 6808 23348 6860
rect 26148 6808 26200 6860
rect 27160 6808 27212 6860
rect 28448 6808 28500 6860
rect 20812 6715 20864 6724
rect 20812 6681 20821 6715
rect 20821 6681 20855 6715
rect 20855 6681 20864 6715
rect 20812 6672 20864 6681
rect 20904 6715 20956 6724
rect 20904 6681 20913 6715
rect 20913 6681 20947 6715
rect 20947 6681 20956 6715
rect 20904 6672 20956 6681
rect 23388 6604 23440 6656
rect 30104 6808 30156 6860
rect 29736 6783 29788 6792
rect 29736 6749 29745 6783
rect 29745 6749 29779 6783
rect 29779 6749 29788 6783
rect 29736 6740 29788 6749
rect 32036 6740 32088 6792
rect 32220 6783 32272 6792
rect 32220 6749 32229 6783
rect 32229 6749 32263 6783
rect 32263 6749 32272 6783
rect 32220 6740 32272 6749
rect 27160 6672 27212 6724
rect 24032 6647 24084 6656
rect 24032 6613 24041 6647
rect 24041 6613 24075 6647
rect 24075 6613 24084 6647
rect 26976 6647 27028 6656
rect 24032 6604 24084 6613
rect 26976 6613 26985 6647
rect 26985 6613 27019 6647
rect 27019 6613 27028 6647
rect 26976 6604 27028 6613
rect 28448 6672 28500 6724
rect 31944 6672 31996 6724
rect 29920 6604 29972 6656
rect 30196 6604 30248 6656
rect 31576 6604 31628 6656
rect 32404 6604 32456 6656
rect 37924 6808 37976 6860
rect 34704 6604 34756 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 20812 6400 20864 6452
rect 24124 6400 24176 6452
rect 27160 6400 27212 6452
rect 31944 6400 31996 6452
rect 22192 6375 22244 6384
rect 22192 6341 22201 6375
rect 22201 6341 22235 6375
rect 22235 6341 22244 6375
rect 22192 6332 22244 6341
rect 24584 6332 24636 6384
rect 26240 6332 26292 6384
rect 27068 6332 27120 6384
rect 27804 6332 27856 6384
rect 28356 6332 28408 6384
rect 29644 6332 29696 6384
rect 29736 6332 29788 6384
rect 30472 6332 30524 6384
rect 32220 6264 32272 6316
rect 33140 6307 33192 6316
rect 22100 6239 22152 6248
rect 22100 6205 22109 6239
rect 22109 6205 22143 6239
rect 22143 6205 22152 6239
rect 22100 6196 22152 6205
rect 22652 6171 22704 6180
rect 22652 6137 22661 6171
rect 22661 6137 22695 6171
rect 22695 6137 22704 6171
rect 22652 6128 22704 6137
rect 32404 6196 32456 6248
rect 33140 6273 33149 6307
rect 33149 6273 33183 6307
rect 33183 6273 33192 6307
rect 33140 6264 33192 6273
rect 29920 6128 29972 6180
rect 23572 6103 23624 6112
rect 23572 6069 23581 6103
rect 23581 6069 23615 6103
rect 23615 6069 23624 6103
rect 23572 6060 23624 6069
rect 24492 6060 24544 6112
rect 25780 6103 25832 6112
rect 25780 6069 25789 6103
rect 25789 6069 25823 6103
rect 25823 6069 25832 6103
rect 25780 6060 25832 6069
rect 27988 6060 28040 6112
rect 30840 6060 30892 6112
rect 31024 6103 31076 6112
rect 31024 6069 31033 6103
rect 31033 6069 31067 6103
rect 31067 6069 31076 6103
rect 31024 6060 31076 6069
rect 31116 6060 31168 6112
rect 31668 6060 31720 6112
rect 32036 6060 32088 6112
rect 34796 6060 34848 6112
rect 35532 6103 35584 6112
rect 35532 6069 35541 6103
rect 35541 6069 35575 6103
rect 35575 6069 35584 6103
rect 35532 6060 35584 6069
rect 36084 6103 36136 6112
rect 36084 6069 36093 6103
rect 36093 6069 36127 6103
rect 36127 6069 36136 6103
rect 36084 6060 36136 6069
rect 37464 6060 37516 6112
rect 38200 6103 38252 6112
rect 38200 6069 38209 6103
rect 38209 6069 38243 6103
rect 38243 6069 38252 6103
rect 38200 6060 38252 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 24584 5856 24636 5908
rect 36176 5856 36228 5908
rect 26608 5788 26660 5840
rect 29184 5831 29236 5840
rect 29184 5797 29193 5831
rect 29193 5797 29227 5831
rect 29227 5797 29236 5831
rect 29184 5788 29236 5797
rect 24032 5720 24084 5772
rect 27252 5720 27304 5772
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 27436 5695 27488 5704
rect 27436 5661 27445 5695
rect 27445 5661 27479 5695
rect 27479 5661 27488 5695
rect 27436 5652 27488 5661
rect 20720 5516 20772 5568
rect 22192 5516 22244 5568
rect 22284 5559 22336 5568
rect 22284 5525 22293 5559
rect 22293 5525 22327 5559
rect 22327 5525 22336 5559
rect 24584 5559 24636 5568
rect 22284 5516 22336 5525
rect 24584 5525 24593 5559
rect 24593 5525 24627 5559
rect 24627 5525 24636 5559
rect 24584 5516 24636 5525
rect 31116 5584 31168 5636
rect 31208 5627 31260 5636
rect 31208 5593 31217 5627
rect 31217 5593 31251 5627
rect 31251 5593 31260 5627
rect 31208 5584 31260 5593
rect 28724 5516 28776 5568
rect 29092 5516 29144 5568
rect 31392 5516 31444 5568
rect 31668 5720 31720 5772
rect 32312 5720 32364 5772
rect 33692 5788 33744 5840
rect 32220 5652 32272 5704
rect 32864 5695 32916 5704
rect 32864 5661 32873 5695
rect 32873 5661 32907 5695
rect 32907 5661 32916 5695
rect 32864 5652 32916 5661
rect 31668 5584 31720 5636
rect 33232 5652 33284 5704
rect 34428 5652 34480 5704
rect 38292 5695 38344 5704
rect 38292 5661 38301 5695
rect 38301 5661 38335 5695
rect 38335 5661 38344 5695
rect 38292 5652 38344 5661
rect 32220 5516 32272 5568
rect 34796 5584 34848 5636
rect 35532 5559 35584 5568
rect 35532 5525 35541 5559
rect 35541 5525 35575 5559
rect 35575 5525 35584 5559
rect 35532 5516 35584 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 22100 5355 22152 5364
rect 22100 5321 22109 5355
rect 22109 5321 22143 5355
rect 22143 5321 22152 5355
rect 22100 5312 22152 5321
rect 24584 5312 24636 5364
rect 25780 5312 25832 5364
rect 26700 5312 26752 5364
rect 27436 5312 27488 5364
rect 28356 5312 28408 5364
rect 29460 5312 29512 5364
rect 29920 5312 29972 5364
rect 23572 5244 23624 5296
rect 27528 5244 27580 5296
rect 28908 5244 28960 5296
rect 31024 5244 31076 5296
rect 33140 5287 33192 5296
rect 21272 5176 21324 5228
rect 22284 5176 22336 5228
rect 22744 5176 22796 5228
rect 28356 5219 28408 5228
rect 20536 5151 20588 5160
rect 20536 5117 20545 5151
rect 20545 5117 20579 5151
rect 20579 5117 20588 5151
rect 20536 5108 20588 5117
rect 23388 5151 23440 5160
rect 23388 5117 23397 5151
rect 23397 5117 23431 5151
rect 23431 5117 23440 5151
rect 23388 5108 23440 5117
rect 20444 5040 20496 5092
rect 20904 5040 20956 5092
rect 25596 5108 25648 5160
rect 28356 5185 28365 5219
rect 28365 5185 28399 5219
rect 28399 5185 28408 5219
rect 28356 5176 28408 5185
rect 33140 5253 33149 5287
rect 33149 5253 33183 5287
rect 33183 5253 33192 5287
rect 33140 5244 33192 5253
rect 29092 5108 29144 5160
rect 29276 5108 29328 5160
rect 32864 5219 32916 5228
rect 32864 5185 32873 5219
rect 32873 5185 32907 5219
rect 32907 5185 32916 5219
rect 35532 5244 35584 5296
rect 36452 5287 36504 5296
rect 36452 5253 36461 5287
rect 36461 5253 36495 5287
rect 36495 5253 36504 5287
rect 36452 5244 36504 5253
rect 32864 5176 32916 5185
rect 34428 5176 34480 5228
rect 33784 5108 33836 5160
rect 26976 5040 27028 5092
rect 31392 5040 31444 5092
rect 22100 4972 22152 5024
rect 29000 4972 29052 5024
rect 31944 4972 31996 5024
rect 34520 4972 34572 5024
rect 36544 4972 36596 5024
rect 38292 5015 38344 5024
rect 38292 4981 38301 5015
rect 38301 4981 38335 5015
rect 38335 4981 38344 5015
rect 38292 4972 38344 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 20904 4768 20956 4820
rect 24400 4768 24452 4820
rect 26792 4768 26844 4820
rect 22100 4675 22152 4684
rect 22100 4641 22109 4675
rect 22109 4641 22143 4675
rect 22143 4641 22152 4675
rect 26056 4700 26108 4752
rect 28356 4768 28408 4820
rect 28540 4743 28592 4752
rect 28540 4709 28549 4743
rect 28549 4709 28583 4743
rect 28583 4709 28592 4743
rect 28540 4700 28592 4709
rect 22100 4632 22152 4641
rect 25412 4632 25464 4684
rect 25872 4632 25924 4684
rect 26148 4632 26200 4684
rect 29092 4768 29144 4820
rect 30748 4768 30800 4820
rect 31024 4768 31076 4820
rect 32128 4811 32180 4820
rect 32128 4777 32137 4811
rect 32137 4777 32171 4811
rect 32171 4777 32180 4811
rect 32128 4768 32180 4777
rect 34060 4811 34112 4820
rect 34060 4777 34069 4811
rect 34069 4777 34103 4811
rect 34103 4777 34112 4811
rect 34060 4768 34112 4777
rect 36452 4768 36504 4820
rect 31116 4700 31168 4752
rect 30104 4632 30156 4684
rect 31300 4632 31352 4684
rect 22192 4564 22244 4616
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 26700 4564 26752 4616
rect 29276 4564 29328 4616
rect 32864 4607 32916 4616
rect 20628 4471 20680 4480
rect 20628 4437 20637 4471
rect 20637 4437 20671 4471
rect 20671 4437 20680 4471
rect 20628 4428 20680 4437
rect 23388 4471 23440 4480
rect 23388 4437 23397 4471
rect 23397 4437 23431 4471
rect 23431 4437 23440 4471
rect 23388 4428 23440 4437
rect 29184 4496 29236 4548
rect 32036 4496 32088 4548
rect 32864 4573 32873 4607
rect 32873 4573 32907 4607
rect 32907 4573 32916 4607
rect 32864 4564 32916 4573
rect 33784 4564 33836 4616
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 37832 4564 37884 4573
rect 33140 4496 33192 4548
rect 34612 4496 34664 4548
rect 33416 4471 33468 4480
rect 33416 4437 33425 4471
rect 33425 4437 33459 4471
rect 33459 4437 33468 4471
rect 33416 4428 33468 4437
rect 34888 4471 34940 4480
rect 34888 4437 34897 4471
rect 34897 4437 34931 4471
rect 34931 4437 34940 4471
rect 34888 4428 34940 4437
rect 35992 4471 36044 4480
rect 35992 4437 36001 4471
rect 36001 4437 36035 4471
rect 36035 4437 36044 4471
rect 35992 4428 36044 4437
rect 38016 4471 38068 4480
rect 38016 4437 38025 4471
rect 38025 4437 38059 4471
rect 38059 4437 38068 4471
rect 38016 4428 38068 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 20536 4224 20588 4276
rect 24584 4224 24636 4276
rect 34428 4224 34480 4276
rect 35532 4224 35584 4276
rect 20536 4088 20588 4140
rect 22836 4088 22888 4140
rect 23204 4088 23256 4140
rect 25412 4131 25464 4140
rect 25412 4097 25421 4131
rect 25421 4097 25455 4131
rect 25455 4097 25464 4131
rect 25412 4088 25464 4097
rect 25504 4088 25556 4140
rect 30196 4131 30248 4140
rect 30196 4097 30205 4131
rect 30205 4097 30239 4131
rect 30239 4097 30248 4131
rect 30196 4088 30248 4097
rect 30748 4088 30800 4140
rect 31116 4131 31168 4140
rect 31116 4097 31125 4131
rect 31125 4097 31159 4131
rect 31159 4097 31168 4131
rect 31116 4088 31168 4097
rect 32864 4088 32916 4140
rect 33784 4131 33836 4140
rect 33784 4097 33793 4131
rect 33793 4097 33827 4131
rect 33827 4097 33836 4131
rect 33784 4088 33836 4097
rect 34244 4088 34296 4140
rect 38016 4131 38068 4140
rect 38016 4097 38025 4131
rect 38025 4097 38059 4131
rect 38059 4097 38068 4131
rect 38016 4088 38068 4097
rect 23388 4063 23440 4072
rect 23388 4029 23397 4063
rect 23397 4029 23431 4063
rect 23431 4029 23440 4063
rect 23388 4020 23440 4029
rect 27344 4020 27396 4072
rect 29920 4063 29972 4072
rect 29920 4029 29929 4063
rect 29929 4029 29963 4063
rect 29963 4029 29972 4063
rect 29920 4020 29972 4029
rect 30288 4020 30340 4072
rect 1492 3884 1544 3936
rect 20628 3884 20680 3936
rect 24768 3952 24820 4004
rect 26240 3884 26292 3936
rect 27252 3927 27304 3936
rect 27252 3893 27261 3927
rect 27261 3893 27295 3927
rect 27295 3893 27304 3927
rect 27252 3884 27304 3893
rect 30196 3884 30248 3936
rect 31208 3884 31260 3936
rect 32220 3884 32272 3936
rect 32404 3927 32456 3936
rect 32404 3893 32413 3927
rect 32413 3893 32447 3927
rect 32447 3893 32456 3927
rect 32404 3884 32456 3893
rect 32496 3884 32548 3936
rect 33692 3927 33744 3936
rect 33692 3893 33701 3927
rect 33701 3893 33735 3927
rect 33735 3893 33744 3927
rect 33692 3884 33744 3893
rect 34152 3884 34204 3936
rect 34888 3927 34940 3936
rect 34888 3893 34897 3927
rect 34897 3893 34931 3927
rect 34931 3893 34940 3927
rect 34888 3884 34940 3893
rect 35532 3884 35584 3936
rect 37188 3884 37240 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 20444 3723 20496 3732
rect 20444 3689 20453 3723
rect 20453 3689 20487 3723
rect 20487 3689 20496 3723
rect 20444 3680 20496 3689
rect 20536 3680 20588 3732
rect 28632 3723 28684 3732
rect 24124 3612 24176 3664
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 24952 3544 25004 3596
rect 26424 3544 26476 3596
rect 1584 3408 1636 3460
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 20536 3476 20588 3528
rect 21364 3476 21416 3528
rect 22192 3476 22244 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 22652 3408 22704 3460
rect 24768 3408 24820 3460
rect 26608 3408 26660 3460
rect 26148 3340 26200 3392
rect 26332 3383 26384 3392
rect 26332 3349 26341 3383
rect 26341 3349 26375 3383
rect 26375 3349 26384 3383
rect 26332 3340 26384 3349
rect 28632 3689 28641 3723
rect 28641 3689 28675 3723
rect 28675 3689 28684 3723
rect 28632 3680 28684 3689
rect 29000 3612 29052 3664
rect 26792 3544 26844 3596
rect 27252 3544 27304 3596
rect 34428 3680 34480 3732
rect 35532 3723 35584 3732
rect 35532 3689 35541 3723
rect 35541 3689 35575 3723
rect 35575 3689 35584 3723
rect 35532 3680 35584 3689
rect 31300 3612 31352 3664
rect 29276 3544 29328 3596
rect 30564 3544 30616 3596
rect 31208 3544 31260 3596
rect 32588 3544 32640 3596
rect 35992 3612 36044 3664
rect 29000 3476 29052 3528
rect 31576 3476 31628 3528
rect 31944 3519 31996 3528
rect 31944 3485 31953 3519
rect 31953 3485 31987 3519
rect 31987 3485 31996 3519
rect 31944 3476 31996 3485
rect 34520 3544 34572 3596
rect 34244 3476 34296 3528
rect 34888 3519 34940 3528
rect 34888 3485 34897 3519
rect 34897 3485 34931 3519
rect 34931 3485 34940 3519
rect 34888 3476 34940 3485
rect 38292 3519 38344 3528
rect 27160 3451 27212 3460
rect 27160 3417 27169 3451
rect 27169 3417 27203 3451
rect 27203 3417 27212 3451
rect 38292 3485 38301 3519
rect 38301 3485 38335 3519
rect 38335 3485 38344 3519
rect 38292 3476 38344 3485
rect 27160 3408 27212 3417
rect 28724 3340 28776 3392
rect 36636 3383 36688 3392
rect 36636 3349 36645 3383
rect 36645 3349 36679 3383
rect 36679 3349 36688 3383
rect 36636 3340 36688 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3148 3068 3200 3120
rect 21364 3179 21416 3188
rect 21364 3145 21373 3179
rect 21373 3145 21407 3179
rect 21407 3145 21416 3179
rect 21364 3136 21416 3145
rect 22192 3136 22244 3188
rect 18328 3000 18380 3052
rect 19248 3000 19300 3052
rect 20 2932 72 2984
rect 1492 2932 1544 2984
rect 21272 3068 21324 3120
rect 23112 3068 23164 3120
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 23020 3000 23072 3052
rect 23388 3136 23440 3188
rect 26332 3136 26384 3188
rect 26608 3136 26660 3188
rect 27252 3179 27304 3188
rect 23664 3068 23716 3120
rect 25228 3068 25280 3120
rect 25504 3068 25556 3120
rect 24860 3000 24912 3052
rect 25596 3000 25648 3052
rect 25872 3000 25924 3052
rect 27252 3145 27261 3179
rect 27261 3145 27295 3179
rect 27295 3145 27304 3179
rect 27252 3136 27304 3145
rect 28080 3179 28132 3188
rect 28080 3145 28089 3179
rect 28089 3145 28123 3179
rect 28123 3145 28132 3179
rect 28080 3136 28132 3145
rect 29092 3136 29144 3188
rect 31392 3136 31444 3188
rect 34152 3136 34204 3188
rect 35348 3179 35400 3188
rect 35348 3145 35357 3179
rect 35357 3145 35391 3179
rect 35391 3145 35400 3179
rect 35348 3136 35400 3145
rect 35532 3136 35584 3188
rect 30196 3068 30248 3120
rect 31944 3068 31996 3120
rect 32404 3068 32456 3120
rect 28724 2975 28776 2984
rect 5540 2864 5592 2916
rect 20076 2864 20128 2916
rect 28724 2941 28733 2975
rect 28733 2941 28767 2975
rect 28767 2941 28776 2975
rect 28724 2932 28776 2941
rect 30748 3043 30800 3052
rect 30748 3009 30757 3043
rect 30757 3009 30791 3043
rect 30791 3009 30800 3043
rect 30748 3000 30800 3009
rect 30380 2932 30432 2984
rect 30472 2975 30524 2984
rect 30472 2941 30481 2975
rect 30481 2941 30515 2975
rect 30515 2941 30524 2975
rect 30472 2932 30524 2941
rect 25228 2864 25280 2916
rect 3792 2839 3844 2848
rect 3792 2805 3801 2839
rect 3801 2805 3835 2839
rect 3835 2805 3844 2839
rect 3792 2796 3844 2805
rect 14556 2796 14608 2848
rect 18328 2796 18380 2848
rect 23664 2796 23716 2848
rect 24768 2796 24820 2848
rect 25136 2796 25188 2848
rect 27068 2864 27120 2916
rect 27252 2864 27304 2916
rect 29000 2864 29052 2916
rect 30104 2796 30156 2848
rect 30288 2796 30340 2848
rect 32496 3000 32548 3052
rect 31484 2932 31536 2984
rect 31852 2932 31904 2984
rect 34612 3111 34664 3120
rect 34612 3077 34621 3111
rect 34621 3077 34655 3111
rect 34655 3077 34664 3111
rect 34612 3068 34664 3077
rect 34888 3000 34940 3052
rect 34244 2932 34296 2984
rect 36544 3000 36596 3052
rect 38016 3043 38068 3052
rect 38016 3009 38025 3043
rect 38025 3009 38059 3043
rect 38059 3009 38068 3043
rect 38016 3000 38068 3009
rect 38200 3000 38252 3052
rect 39304 3000 39356 3052
rect 31392 2864 31444 2916
rect 32312 2839 32364 2848
rect 32312 2805 32321 2839
rect 32321 2805 32355 2839
rect 32355 2805 32364 2839
rect 32312 2796 32364 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 10784 2592 10836 2644
rect 19156 2592 19208 2644
rect 22928 2592 22980 2644
rect 26332 2592 26384 2644
rect 26516 2592 26568 2644
rect 29368 2592 29420 2644
rect 30656 2592 30708 2644
rect 35532 2592 35584 2644
rect 12072 2524 12124 2576
rect 1952 2456 2004 2508
rect 10324 2456 10376 2508
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 21548 2524 21600 2576
rect 37280 2524 37332 2576
rect 14556 2388 14608 2440
rect 3240 2320 3292 2372
rect 3792 2320 3844 2372
rect 9036 2320 9088 2372
rect 9864 2320 9916 2372
rect 1308 2252 1360 2304
rect 5172 2252 5224 2304
rect 7104 2252 7156 2304
rect 12256 2252 12308 2304
rect 14188 2320 14240 2372
rect 15936 2388 15988 2440
rect 18052 2431 18104 2440
rect 18052 2397 18061 2431
rect 18061 2397 18095 2431
rect 18095 2397 18104 2431
rect 21824 2456 21876 2508
rect 22192 2499 22244 2508
rect 22192 2465 22201 2499
rect 22201 2465 22235 2499
rect 22235 2465 22244 2499
rect 22192 2456 22244 2465
rect 22928 2456 22980 2508
rect 23480 2456 23532 2508
rect 24584 2499 24636 2508
rect 24584 2465 24593 2499
rect 24593 2465 24627 2499
rect 24627 2465 24636 2499
rect 24584 2456 24636 2465
rect 18052 2388 18104 2397
rect 21180 2431 21232 2440
rect 21180 2397 21189 2431
rect 21189 2397 21223 2431
rect 21223 2397 21232 2431
rect 21180 2388 21232 2397
rect 26240 2456 26292 2508
rect 26424 2456 26476 2508
rect 27160 2456 27212 2508
rect 27344 2456 27396 2508
rect 29000 2499 29052 2508
rect 29000 2465 29009 2499
rect 29009 2465 29043 2499
rect 29043 2465 29052 2499
rect 29000 2456 29052 2465
rect 31944 2456 31996 2508
rect 37464 2499 37516 2508
rect 37464 2465 37473 2499
rect 37473 2465 37507 2499
rect 37507 2465 37516 2499
rect 37464 2456 37516 2465
rect 37740 2499 37792 2508
rect 37740 2465 37749 2499
rect 37749 2465 37783 2499
rect 37783 2465 37792 2499
rect 37740 2456 37792 2465
rect 32956 2431 33008 2440
rect 32956 2397 32965 2431
rect 32965 2397 32999 2431
rect 32999 2397 33008 2431
rect 32956 2388 33008 2397
rect 34428 2388 34480 2440
rect 34704 2388 34756 2440
rect 36084 2388 36136 2440
rect 38016 2388 38068 2440
rect 24584 2320 24636 2372
rect 16120 2252 16172 2304
rect 19340 2252 19392 2304
rect 21272 2252 21324 2304
rect 23296 2252 23348 2304
rect 28264 2320 28316 2372
rect 31208 2363 31260 2372
rect 31208 2329 31217 2363
rect 31217 2329 31251 2363
rect 31251 2329 31260 2363
rect 31208 2320 31260 2329
rect 32864 2295 32916 2304
rect 32864 2261 32873 2295
rect 32873 2261 32907 2295
rect 32907 2261 32916 2295
rect 32864 2252 32916 2261
rect 34980 2295 35032 2304
rect 34980 2261 34989 2295
rect 34989 2261 35023 2295
rect 35023 2261 35032 2295
rect 34980 2252 35032 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 24584 2048 24636 2100
rect 32864 2048 32916 2100
rect 18328 1980 18380 2032
rect 34980 1980 35032 2032
rect 26240 1912 26292 1964
rect 33692 1912 33744 1964
rect 28264 1844 28316 1896
rect 33416 1844 33468 1896
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 3238 39200 3294 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 14186 39200 14242 39800
rect 16118 39200 16174 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 23202 39200 23258 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 34150 39200 34206 39800
rect 36082 39200 36138 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 32 36854 60 39200
rect 1320 37126 1348 39200
rect 2778 38176 2834 38185
rect 2778 38111 2834 38120
rect 2320 37256 2372 37262
rect 2320 37198 2372 37204
rect 1308 37120 1360 37126
rect 1308 37062 1360 37068
rect 20 36848 72 36854
rect 20 36790 72 36796
rect 1676 36848 1728 36854
rect 1676 36790 1728 36796
rect 1492 36576 1544 36582
rect 1492 36518 1544 36524
rect 1504 35894 1532 36518
rect 1688 36378 1716 36790
rect 2228 36644 2280 36650
rect 2228 36586 2280 36592
rect 1676 36372 1728 36378
rect 1676 36314 1728 36320
rect 1860 36168 1912 36174
rect 1674 36136 1730 36145
rect 1860 36110 1912 36116
rect 1674 36071 1730 36080
rect 1688 36038 1716 36071
rect 1676 36032 1728 36038
rect 1676 35974 1728 35980
rect 1504 35866 1808 35894
rect 1676 34400 1728 34406
rect 1676 34342 1728 34348
rect 1688 34105 1716 34342
rect 1674 34096 1730 34105
rect 1674 34031 1730 34040
rect 1584 32428 1636 32434
rect 1584 32370 1636 32376
rect 1596 32065 1624 32370
rect 1582 32056 1638 32065
rect 1582 31991 1584 32000
rect 1636 31991 1638 32000
rect 1584 31962 1636 31968
rect 1674 30696 1730 30705
rect 1674 30631 1730 30640
rect 1688 30598 1716 30631
rect 1676 30592 1728 30598
rect 1676 30534 1728 30540
rect 1676 29028 1728 29034
rect 1676 28970 1728 28976
rect 1688 28665 1716 28970
rect 1674 28656 1730 28665
rect 1674 28591 1730 28600
rect 1584 26920 1636 26926
rect 1584 26862 1636 26868
rect 1596 26625 1624 26862
rect 1582 26616 1638 26625
rect 1582 26551 1584 26560
rect 1636 26551 1638 26560
rect 1584 26522 1636 26528
rect 1676 24608 1728 24614
rect 1674 24576 1676 24585
rect 1728 24576 1730 24585
rect 1674 24511 1730 24520
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1688 22642 1716 22918
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 1688 22545 1716 22578
rect 1674 22536 1730 22545
rect 1674 22471 1730 22480
rect 1584 20868 1636 20874
rect 1584 20810 1636 20816
rect 1596 20534 1624 20810
rect 1584 20528 1636 20534
rect 1582 20496 1584 20505
rect 1636 20496 1638 20505
rect 1582 20431 1638 20440
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 19145 1624 19246
rect 1582 19136 1638 19145
rect 1582 19071 1638 19080
rect 1596 18970 1624 19071
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1674 17096 1730 17105
rect 1674 17031 1676 17040
rect 1728 17031 1730 17040
rect 1676 17002 1728 17008
rect 1780 16574 1808 35866
rect 1872 35834 1900 36110
rect 1860 35828 1912 35834
rect 1860 35770 1912 35776
rect 2136 34536 2188 34542
rect 2136 34478 2188 34484
rect 1860 29164 1912 29170
rect 1860 29106 1912 29112
rect 1872 26450 1900 29106
rect 1860 26444 1912 26450
rect 1860 26386 1912 26392
rect 2044 24812 2096 24818
rect 2044 24754 2096 24760
rect 1860 22500 1912 22506
rect 1860 22442 1912 22448
rect 1872 20262 1900 22442
rect 2056 21894 2084 24754
rect 2044 21888 2096 21894
rect 2044 21830 2096 21836
rect 1860 20256 1912 20262
rect 1860 20198 1912 20204
rect 2148 19990 2176 34478
rect 2240 28558 2268 36586
rect 2332 36582 2360 37198
rect 2412 37188 2464 37194
rect 2412 37130 2464 37136
rect 2320 36576 2372 36582
rect 2320 36518 2372 36524
rect 2320 30592 2372 30598
rect 2320 30534 2372 30540
rect 2228 28552 2280 28558
rect 2228 28494 2280 28500
rect 2228 26920 2280 26926
rect 2228 26862 2280 26868
rect 2136 19984 2188 19990
rect 2136 19926 2188 19932
rect 2240 18766 2268 26862
rect 2332 20806 2360 30534
rect 2320 20800 2372 20806
rect 2320 20742 2372 20748
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2240 16794 2268 18702
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2240 16590 2268 16730
rect 2228 16584 2280 16590
rect 1780 16546 1900 16574
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1688 15065 1716 15302
rect 1674 15056 1730 15065
rect 1674 14991 1730 15000
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1688 13025 1716 13126
rect 1674 13016 1730 13025
rect 1674 12951 1730 12960
rect 1780 11150 1808 16390
rect 1872 14618 1900 16546
rect 2228 16526 2280 16532
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1964 13258 1992 14282
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1676 11008 1728 11014
rect 1674 10976 1676 10985
rect 1728 10976 1730 10985
rect 1674 10911 1730 10920
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1872 10130 1900 10610
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9654 1624 9998
rect 1584 9648 1636 9654
rect 1582 9616 1584 9625
rect 1636 9616 1638 9625
rect 1582 9551 1638 9560
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7585 1716 7686
rect 1674 7576 1730 7585
rect 1674 7511 1730 7520
rect 1676 5568 1728 5574
rect 1674 5536 1676 5545
rect 1728 5536 1730 5545
rect 1674 5471 1730 5480
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1504 2990 1532 3878
rect 1674 3496 1730 3505
rect 1584 3460 1636 3466
rect 1674 3431 1730 3440
rect 1584 3402 1636 3408
rect 20 2984 72 2990
rect 20 2926 72 2932
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 32 800 60 2926
rect 1596 2446 1624 3402
rect 1688 3398 1716 3431
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1964 2514 1992 13194
rect 2424 10742 2452 37130
rect 2792 37126 2820 38111
rect 3252 37126 3280 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3424 37256 3476 37262
rect 3424 37198 3476 37204
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 3240 37120 3292 37126
rect 3240 37062 3292 37068
rect 3436 36922 3464 37198
rect 5184 37126 5212 39200
rect 5540 37256 5592 37262
rect 5540 37198 5592 37204
rect 5172 37120 5224 37126
rect 5172 37062 5224 37068
rect 3424 36916 3476 36922
rect 3424 36858 3476 36864
rect 4804 36576 4856 36582
rect 4804 36518 4856 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 2504 35692 2556 35698
rect 2504 35634 2556 35640
rect 2516 35494 2544 35634
rect 2504 35488 2556 35494
rect 2504 35430 2556 35436
rect 2516 12306 2544 35430
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 2688 32292 2740 32298
rect 2688 32234 2740 32240
rect 2700 27878 2728 32234
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4816 23866 4844 36518
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5552 23322 5580 37198
rect 7116 37126 7144 39200
rect 9048 37262 9076 39200
rect 10336 37330 10364 39200
rect 12268 37330 12296 39200
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 11704 37324 11756 37330
rect 11704 37266 11756 37272
rect 12256 37324 12308 37330
rect 12256 37266 12308 37272
rect 9036 37256 9088 37262
rect 9036 37198 9088 37204
rect 10876 37256 10928 37262
rect 10876 37198 10928 37204
rect 7104 37120 7156 37126
rect 7104 37062 7156 37068
rect 8024 37120 8076 37126
rect 8024 37062 8076 37068
rect 9312 37120 9364 37126
rect 9312 37062 9364 37068
rect 8036 32230 8064 37062
rect 8024 32224 8076 32230
rect 8024 32166 8076 32172
rect 9324 30734 9352 37062
rect 10888 36786 10916 37198
rect 11716 36922 11744 37266
rect 14200 37126 14228 39200
rect 16132 37466 16160 39200
rect 16120 37460 16172 37466
rect 16120 37402 16172 37408
rect 14280 37256 14332 37262
rect 14280 37198 14332 37204
rect 17132 37256 17184 37262
rect 17132 37198 17184 37204
rect 17868 37256 17920 37262
rect 17868 37198 17920 37204
rect 14188 37120 14240 37126
rect 14188 37062 14240 37068
rect 11704 36916 11756 36922
rect 11704 36858 11756 36864
rect 10876 36780 10928 36786
rect 10876 36722 10928 36728
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 14292 29306 14320 37198
rect 17144 36718 17172 37198
rect 17880 36922 17908 37198
rect 18064 37126 18092 39200
rect 19996 37330 20024 39200
rect 19984 37324 20036 37330
rect 19984 37266 20036 37272
rect 20720 37188 20772 37194
rect 20720 37130 20772 37136
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20732 36922 20760 37130
rect 21284 37126 21312 39200
rect 23216 37330 23244 39200
rect 23204 37324 23256 37330
rect 23204 37266 23256 37272
rect 21364 37256 21416 37262
rect 21364 37198 21416 37204
rect 21272 37120 21324 37126
rect 21272 37062 21324 37068
rect 21376 36922 21404 37198
rect 23388 37188 23440 37194
rect 23388 37130 23440 37136
rect 24584 37188 24636 37194
rect 24584 37130 24636 37136
rect 17868 36916 17920 36922
rect 17868 36858 17920 36864
rect 20720 36916 20772 36922
rect 20720 36858 20772 36864
rect 21364 36916 21416 36922
rect 21364 36858 21416 36864
rect 23400 36854 23428 37130
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 23388 36848 23440 36854
rect 23388 36790 23440 36796
rect 17684 36780 17736 36786
rect 17684 36722 17736 36728
rect 22744 36780 22796 36786
rect 22744 36722 22796 36728
rect 17132 36712 17184 36718
rect 17132 36654 17184 36660
rect 17696 30258 17724 36722
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 17684 30252 17736 30258
rect 17684 30194 17736 30200
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 16580 29028 16632 29034
rect 16580 28970 16632 28976
rect 7472 23588 7524 23594
rect 7472 23530 7524 23536
rect 5540 23316 5592 23322
rect 5540 23258 5592 23264
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 6840 15706 6868 17138
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12442 4660 13262
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5000 11354 5028 12038
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 3160 2446 3188 3062
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 1596 1465 1624 2382
rect 3804 2378 3832 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5552 2446 5580 2858
rect 7484 2446 7512 23530
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 9876 2378 9904 19654
rect 10152 16590 10180 21830
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10612 12986 10640 13126
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10796 2650 10824 16594
rect 12084 14414 12112 22918
rect 16592 20874 16620 28970
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 16592 19854 16620 20810
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12176 15162 12204 15302
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 12084 2582 12112 14350
rect 15764 12238 15792 19314
rect 19260 18834 19288 19722
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19156 15428 19208 15434
rect 19156 15370 19208 15376
rect 19168 13938 19196 15370
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16408 11354 16436 12174
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16408 11150 16436 11290
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 10062 14320 10610
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14384 10266 14412 10542
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14108 7546 14136 7822
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 12072 2576 12124 2582
rect 12072 2518 12124 2524
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 3252 800 3280 2314
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 5184 800 5212 2246
rect 7116 800 7144 2246
rect 9048 800 9076 2314
rect 10336 800 10364 2450
rect 14568 2446 14596 2790
rect 15948 2446 15976 10950
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17236 10266 17264 10678
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18340 2854 18368 2994
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 800 12296 2246
rect 14200 800 14228 2314
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16132 800 16160 2246
rect 18064 800 18092 2382
rect 18340 2038 18368 2790
rect 19168 2650 19196 13874
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11626 20024 20810
rect 20088 19378 20116 29990
rect 22756 29170 22784 36722
rect 23400 30734 23428 36790
rect 23860 31482 23888 37062
rect 24032 36780 24084 36786
rect 24032 36722 24084 36728
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 22928 30592 22980 30598
rect 22928 30534 22980 30540
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22468 27872 22520 27878
rect 22468 27814 22520 27820
rect 22480 23730 22508 27814
rect 22652 26308 22704 26314
rect 22652 26250 22704 26256
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22296 19922 22324 21966
rect 22572 21690 22600 23598
rect 22664 23186 22692 26250
rect 22652 23180 22704 23186
rect 22652 23122 22704 23128
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22848 22234 22876 23054
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22756 20806 22784 21490
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 21732 18692 21784 18698
rect 21732 18634 21784 18640
rect 21744 17882 21772 18634
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22112 18086 22140 18226
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 22112 17746 22140 18022
rect 22204 17882 22232 19382
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22296 18834 22324 19178
rect 22480 18902 22508 19790
rect 22756 19786 22784 20742
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22468 18896 22520 18902
rect 22468 18838 22520 18844
rect 22560 18896 22612 18902
rect 22560 18838 22612 18844
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22572 18714 22600 18838
rect 22940 18834 22968 30534
rect 23204 29028 23256 29034
rect 23204 28970 23256 28976
rect 23112 28552 23164 28558
rect 23112 28494 23164 28500
rect 23124 26586 23152 28494
rect 23112 26580 23164 26586
rect 23112 26522 23164 26528
rect 23124 26382 23152 26522
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 23020 22568 23072 22574
rect 23020 22510 23072 22516
rect 23032 22098 23060 22510
rect 23020 22092 23072 22098
rect 23020 22034 23072 22040
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23124 21690 23152 21966
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 23216 18986 23244 28970
rect 24044 28218 24072 36722
rect 24216 36576 24268 36582
rect 24216 36518 24268 36524
rect 24228 36378 24256 36518
rect 24216 36372 24268 36378
rect 24216 36314 24268 36320
rect 24308 31340 24360 31346
rect 24308 31282 24360 31288
rect 24320 31142 24348 31282
rect 24308 31136 24360 31142
rect 24308 31078 24360 31084
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 24124 26444 24176 26450
rect 24124 26386 24176 26392
rect 24136 24614 24164 26386
rect 24124 24608 24176 24614
rect 24124 24550 24176 24556
rect 24216 23792 24268 23798
rect 24216 23734 24268 23740
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 23308 23322 23336 23666
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23308 22234 23336 23258
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 24044 21554 24072 21966
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 24044 20806 24072 21490
rect 23388 20800 23440 20806
rect 23388 20742 23440 20748
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 23400 20398 23428 20742
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23308 19514 23336 19790
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23032 18958 23244 18986
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 22480 18686 22600 18714
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21192 16998 21220 17478
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19260 3058 19288 8298
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 20088 2922 20116 16594
rect 21192 16590 21220 16934
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 20260 16516 20312 16522
rect 20260 16458 20312 16464
rect 20272 16182 20300 16458
rect 20260 16176 20312 16182
rect 20260 16118 20312 16124
rect 21192 13938 21220 16526
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21468 15638 21496 16050
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20732 12306 20760 12718
rect 20824 12442 20852 12854
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20916 12322 20944 13126
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20824 12294 20944 12322
rect 20824 12238 20852 12294
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20824 10470 20852 12174
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20824 10266 20852 10406
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20824 8362 20852 8910
rect 20812 8356 20864 8362
rect 20812 8298 20864 8304
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20732 5574 20760 6802
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20824 6458 20852 6666
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 20456 3738 20484 5034
rect 20548 4282 20576 5102
rect 20916 5098 20944 6666
rect 20904 5092 20956 5098
rect 20904 5034 20956 5040
rect 20916 4826 20944 5034
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20640 4162 20668 4422
rect 20548 4146 20668 4162
rect 20536 4140 20668 4146
rect 20588 4134 20668 4140
rect 20536 4082 20588 4088
rect 20548 3738 20576 4082
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 20548 3534 20576 3674
rect 20640 3602 20668 3878
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20076 2916 20128 2922
rect 20076 2858 20128 2864
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 21192 2446 21220 11494
rect 21560 11150 21588 11562
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21362 10704 21418 10713
rect 21362 10639 21364 10648
rect 21416 10639 21418 10648
rect 21364 10610 21416 10616
rect 21560 10198 21588 11086
rect 21548 10192 21600 10198
rect 21548 10134 21600 10140
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 21468 7954 21496 8842
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21364 7812 21416 7818
rect 21364 7754 21416 7760
rect 21376 7546 21404 7754
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21468 6866 21496 7890
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21284 3126 21312 5170
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21376 3194 21404 3470
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21272 3120 21324 3126
rect 21272 3062 21324 3068
rect 21454 3088 21510 3097
rect 21454 3023 21456 3032
rect 21508 3023 21510 3032
rect 21456 2994 21508 3000
rect 21560 2582 21588 10134
rect 21548 2576 21600 2582
rect 21548 2518 21600 2524
rect 21836 2514 21864 16390
rect 22480 15586 22508 18686
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22664 18222 22692 18566
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22572 15706 22600 16458
rect 22664 16250 22692 17478
rect 22756 17202 22784 17614
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22480 15558 22600 15586
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22204 14890 22232 15438
rect 22572 15026 22600 15558
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22192 14884 22244 14890
rect 22192 14826 22244 14832
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22112 12986 22140 14418
rect 22192 14340 22244 14346
rect 22192 14282 22244 14288
rect 22204 14074 22232 14282
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 22388 13394 22416 13806
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22112 12866 22140 12922
rect 22112 12838 22232 12866
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 11898 22140 12582
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22204 11830 22232 12838
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22296 12442 22324 12718
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22296 12306 22324 12378
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 22388 11354 22416 12106
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21928 10742 21956 11018
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 22112 10606 22140 11086
rect 22192 10736 22244 10742
rect 22190 10704 22192 10713
rect 22244 10704 22246 10713
rect 22190 10639 22246 10648
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 22112 9586 22140 10542
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 22376 9988 22428 9994
rect 22376 9930 22428 9936
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22296 9178 22324 9930
rect 22388 9722 22416 9930
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22192 8560 22244 8566
rect 22192 8502 22244 8508
rect 22204 6390 22232 8502
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22296 7886 22324 8366
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22296 6866 22324 7822
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22388 7478 22416 7686
rect 22480 7546 22508 8774
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22192 6384 22244 6390
rect 22192 6326 22244 6332
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22112 5370 22140 6190
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22112 4690 22140 4966
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 22204 4622 22232 5510
rect 22296 5234 22324 5510
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 22204 3194 22232 3470
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22204 2514 22232 3130
rect 22572 2774 22600 14962
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22664 12102 22692 14214
rect 22756 12434 22784 17138
rect 23032 15638 23060 18958
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23216 18714 23244 18770
rect 23124 18686 23244 18714
rect 23124 18222 23152 18686
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 23124 17338 23152 18158
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23124 16726 23152 17274
rect 23204 17060 23256 17066
rect 23204 17002 23256 17008
rect 23112 16720 23164 16726
rect 23112 16662 23164 16668
rect 23216 16538 23244 17002
rect 23308 16794 23336 17546
rect 23400 17134 23428 20334
rect 23676 20058 23704 20470
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23492 18154 23520 19654
rect 23676 19378 23704 19790
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23492 17746 23520 18090
rect 23480 17740 23532 17746
rect 23480 17682 23532 17688
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 23124 16510 23244 16538
rect 23020 15632 23072 15638
rect 23020 15574 23072 15580
rect 23124 15570 23152 16510
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 22836 15428 22888 15434
rect 22836 15370 22888 15376
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 22848 14278 22876 15370
rect 22940 15162 22968 15370
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 23124 14482 23152 15506
rect 23204 15360 23256 15366
rect 23204 15302 23256 15308
rect 23216 14906 23244 15302
rect 23308 15042 23336 16730
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23480 16516 23532 16522
rect 23480 16458 23532 16464
rect 23492 16182 23520 16458
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 23584 15162 23612 16526
rect 23676 15858 23704 19314
rect 23768 18290 23796 20198
rect 24228 19446 24256 23734
rect 24320 20602 24348 31078
rect 24596 22094 24624 37130
rect 25148 37126 25176 39200
rect 27080 37466 27108 39200
rect 27068 37460 27120 37466
rect 27068 37402 27120 37408
rect 26792 37324 26844 37330
rect 26792 37266 26844 37272
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 26424 36848 26476 36854
rect 26424 36790 26476 36796
rect 26056 36712 26108 36718
rect 26056 36654 26108 36660
rect 25504 32428 25556 32434
rect 25504 32370 25556 32376
rect 25516 31346 25544 32370
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25136 31136 25188 31142
rect 25136 31078 25188 31084
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24504 22066 24624 22094
rect 24504 20942 24532 22066
rect 24780 21690 24808 24550
rect 24952 22500 25004 22506
rect 24952 22442 25004 22448
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24400 20800 24452 20806
rect 24400 20742 24452 20748
rect 24308 20596 24360 20602
rect 24308 20538 24360 20544
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23768 16046 23796 18226
rect 24228 17746 24256 19382
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24412 17202 24440 20742
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24412 17066 24440 17138
rect 24400 17060 24452 17066
rect 24400 17002 24452 17008
rect 23940 16176 23992 16182
rect 23940 16118 23992 16124
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23848 15972 23900 15978
rect 23848 15914 23900 15920
rect 23676 15830 23796 15858
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23480 15088 23532 15094
rect 23308 15014 23428 15042
rect 23480 15030 23532 15036
rect 23400 14958 23428 15014
rect 23388 14952 23440 14958
rect 23216 14878 23336 14906
rect 23388 14894 23440 14900
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22848 12850 22876 13670
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 22756 12406 22876 12434
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22652 11620 22704 11626
rect 22652 11562 22704 11568
rect 22664 7954 22692 11562
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22756 8498 22784 10610
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22664 6186 22692 7890
rect 22756 7546 22784 8434
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22756 7002 22784 7482
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22652 6180 22704 6186
rect 22652 6122 22704 6128
rect 22756 5234 22784 6938
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22848 4146 22876 12406
rect 22940 11626 22968 12718
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 22928 11620 22980 11626
rect 22928 11562 22980 11568
rect 23032 11354 23060 11766
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22848 3641 22876 4082
rect 22834 3632 22890 3641
rect 22834 3567 22890 3576
rect 22650 3496 22706 3505
rect 22650 3431 22652 3440
rect 22704 3431 22706 3440
rect 22652 3402 22704 3408
rect 23124 3126 23152 12310
rect 23216 4146 23244 13874
rect 23308 12374 23336 14878
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23400 13394 23428 14350
rect 23492 13530 23520 15030
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23584 14074 23612 14350
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 23676 13938 23704 14214
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23768 13818 23796 15830
rect 23860 15162 23888 15914
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23952 14074 23980 16118
rect 24032 15972 24084 15978
rect 24032 15914 24084 15920
rect 24044 15094 24072 15914
rect 24032 15088 24084 15094
rect 24032 15030 24084 15036
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 23676 13790 23796 13818
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 23296 12164 23348 12170
rect 23296 12106 23348 12112
rect 23308 10810 23336 12106
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 23492 10062 23520 11086
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23308 8566 23336 9522
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23308 8090 23336 8502
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23296 6860 23348 6866
rect 23348 6820 23428 6848
rect 23296 6802 23348 6808
rect 23400 6662 23428 6820
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23400 5166 23428 6598
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23584 5302 23612 6054
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23400 4486 23428 5102
rect 23388 4480 23440 4486
rect 23388 4422 23440 4428
rect 23204 4140 23256 4146
rect 23256 4100 23336 4128
rect 23204 4082 23256 4088
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 23032 2904 23060 2994
rect 23032 2876 23244 2904
rect 22572 2746 22968 2774
rect 22940 2650 22968 2746
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 22940 2514 22968 2586
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22928 2508 22980 2514
rect 22928 2450 22980 2456
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 18328 2032 18380 2038
rect 18328 1974 18380 1980
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21284 800 21312 2246
rect 23216 800 23244 2876
rect 23308 2310 23336 4100
rect 23400 4078 23428 4422
rect 23388 4072 23440 4078
rect 23388 4014 23440 4020
rect 23400 3194 23428 4014
rect 23388 3188 23440 3194
rect 23440 3148 23520 3176
rect 23388 3130 23440 3136
rect 23492 2514 23520 3148
rect 23676 3126 23704 13790
rect 24044 12918 24072 15030
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 23768 11354 23796 12854
rect 24044 11830 24072 12854
rect 24124 12164 24176 12170
rect 24124 12106 24176 12112
rect 24032 11824 24084 11830
rect 24032 11766 24084 11772
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 24136 9518 24164 12106
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24228 10674 24256 11086
rect 24320 11082 24348 13398
rect 24308 11076 24360 11082
rect 24308 11018 24360 11024
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 24136 9042 24164 9454
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 23940 7336 23992 7342
rect 23992 7284 24072 7290
rect 23940 7278 24072 7284
rect 23952 7262 24072 7278
rect 24044 6662 24072 7262
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 24044 5778 24072 6598
rect 24136 6458 24164 7686
rect 24228 7342 24256 10610
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 24124 6452 24176 6458
rect 24124 6394 24176 6400
rect 24032 5772 24084 5778
rect 24032 5714 24084 5720
rect 24136 3670 24164 6394
rect 24412 4826 24440 17002
rect 24596 16114 24624 21286
rect 24964 20398 24992 22442
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24780 18290 24808 18566
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24780 17338 24808 17614
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25056 16658 25084 16934
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24780 16114 24808 16390
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24872 15570 24900 16390
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24596 15094 24624 15506
rect 24584 15088 24636 15094
rect 24584 15030 24636 15036
rect 25148 14414 25176 31078
rect 25780 30184 25832 30190
rect 25780 30126 25832 30132
rect 25688 27872 25740 27878
rect 25688 27814 25740 27820
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25516 22710 25544 22918
rect 25412 22704 25464 22710
rect 25412 22646 25464 22652
rect 25504 22704 25556 22710
rect 25504 22646 25556 22652
rect 25424 22234 25452 22646
rect 25412 22228 25464 22234
rect 25412 22170 25464 22176
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25240 19446 25268 20334
rect 25332 20058 25360 20470
rect 25320 20052 25372 20058
rect 25320 19994 25372 20000
rect 25504 19712 25556 19718
rect 25504 19654 25556 19660
rect 25228 19440 25280 19446
rect 25228 19382 25280 19388
rect 25412 19236 25464 19242
rect 25412 19178 25464 19184
rect 25424 18358 25452 19178
rect 25516 18766 25544 19654
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 25412 18352 25464 18358
rect 25412 18294 25464 18300
rect 25320 16788 25372 16794
rect 25320 16730 25372 16736
rect 25332 16522 25360 16730
rect 25320 16516 25372 16522
rect 25320 16458 25372 16464
rect 25136 14408 25188 14414
rect 25136 14350 25188 14356
rect 25148 14006 25176 14350
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24504 13462 24532 13806
rect 24492 13456 24544 13462
rect 24492 13398 24544 13404
rect 24584 13252 24636 13258
rect 24584 13194 24636 13200
rect 24768 13252 24820 13258
rect 24768 13194 24820 13200
rect 25228 13252 25280 13258
rect 25228 13194 25280 13200
rect 24596 12170 24624 13194
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24492 11008 24544 11014
rect 24492 10950 24544 10956
rect 24504 9178 24532 10950
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24596 8090 24624 11766
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24688 10130 24716 11018
rect 24780 10810 24808 13194
rect 25240 12714 25268 13194
rect 25228 12708 25280 12714
rect 25228 12650 25280 12656
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24872 11286 24900 11630
rect 24860 11280 24912 11286
rect 24860 11222 24912 11228
rect 24872 10810 24900 11222
rect 24964 11218 24992 12242
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24964 10130 24992 11154
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24688 9654 24716 9862
rect 24676 9648 24728 9654
rect 24676 9590 24728 9596
rect 25044 9444 25096 9450
rect 25044 9386 25096 9392
rect 25056 9178 25084 9386
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24872 8430 24900 8910
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24584 8084 24636 8090
rect 24584 8026 24636 8032
rect 24492 7336 24544 7342
rect 24492 7278 24544 7284
rect 24504 6118 24532 7278
rect 25148 7206 25176 11630
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25332 9654 25360 10746
rect 25412 10736 25464 10742
rect 25412 10678 25464 10684
rect 25320 9648 25372 9654
rect 25320 9590 25372 9596
rect 25424 8634 25452 10678
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 24584 6384 24636 6390
rect 24584 6326 24636 6332
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24596 5914 24624 6326
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24596 5370 24624 5510
rect 24584 5364 24636 5370
rect 24584 5306 24636 5312
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 24596 4622 24624 5306
rect 25412 4684 25464 4690
rect 25412 4626 25464 4632
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24596 4282 24624 4558
rect 24584 4276 24636 4282
rect 24584 4218 24636 4224
rect 24124 3664 24176 3670
rect 24124 3606 24176 3612
rect 24596 3534 24624 4218
rect 25424 4146 25452 4626
rect 25516 4146 25544 18702
rect 25700 17746 25728 27814
rect 25792 24410 25820 30126
rect 26068 28218 26096 36654
rect 26436 35894 26464 36790
rect 26436 35866 26556 35894
rect 26056 28212 26108 28218
rect 26056 28154 26108 28160
rect 25780 24404 25832 24410
rect 25780 24346 25832 24352
rect 25792 23730 25820 24346
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 26332 23724 26384 23730
rect 26332 23666 26384 23672
rect 25792 23322 25820 23666
rect 26344 23633 26372 23666
rect 26330 23624 26386 23633
rect 26330 23559 26386 23568
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 25792 23118 25820 23258
rect 25780 23112 25832 23118
rect 25780 23054 25832 23060
rect 26424 20256 26476 20262
rect 26424 20198 26476 20204
rect 26436 19446 26464 20198
rect 26332 19440 26384 19446
rect 26332 19382 26384 19388
rect 26424 19440 26476 19446
rect 26424 19382 26476 19388
rect 26344 18970 26372 19382
rect 26332 18964 26384 18970
rect 26332 18906 26384 18912
rect 26528 18358 26556 35866
rect 26332 18352 26384 18358
rect 26332 18294 26384 18300
rect 26516 18352 26568 18358
rect 26516 18294 26568 18300
rect 26344 17882 26372 18294
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 25688 17740 25740 17746
rect 25688 17682 25740 17688
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25884 17338 25912 17614
rect 26240 17536 26292 17542
rect 26240 17478 26292 17484
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 26252 16046 26280 17478
rect 26528 17270 26556 18294
rect 26700 17740 26752 17746
rect 26700 17682 26752 17688
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26516 17264 26568 17270
rect 26516 17206 26568 17212
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26240 16040 26292 16046
rect 26240 15982 26292 15988
rect 25688 15904 25740 15910
rect 25688 15846 25740 15852
rect 25700 15570 25728 15846
rect 26252 15638 26280 15982
rect 26240 15632 26292 15638
rect 26240 15574 26292 15580
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25608 12850 25636 14962
rect 25700 14006 25728 15506
rect 26344 15502 26372 17070
rect 26528 16658 26556 17206
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 25872 15428 25924 15434
rect 25872 15370 25924 15376
rect 25884 15026 25912 15370
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 25872 15020 25924 15026
rect 25872 14962 25924 14968
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25700 13530 25728 13942
rect 26252 13870 26280 14962
rect 26344 14482 26372 15302
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26436 14482 26464 14894
rect 26332 14476 26384 14482
rect 26332 14418 26384 14424
rect 26424 14476 26476 14482
rect 26424 14418 26476 14424
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26240 13864 26292 13870
rect 26240 13806 26292 13812
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25608 7002 25636 12786
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25700 9110 25728 12106
rect 25792 11898 25820 13262
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25884 11830 25912 13126
rect 25976 12986 26004 13262
rect 25964 12980 26016 12986
rect 25964 12922 26016 12928
rect 26252 12434 26280 13806
rect 26344 12986 26372 14010
rect 26332 12980 26384 12986
rect 26332 12922 26384 12928
rect 26252 12406 26372 12434
rect 25872 11824 25924 11830
rect 25872 11766 25924 11772
rect 25688 9104 25740 9110
rect 25688 9046 25740 9052
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25700 7342 25728 7822
rect 25688 7336 25740 7342
rect 25688 7278 25740 7284
rect 25780 7200 25832 7206
rect 25780 7142 25832 7148
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 25608 5166 25636 6938
rect 25792 6118 25820 7142
rect 25780 6112 25832 6118
rect 25780 6054 25832 6060
rect 25792 5370 25820 6054
rect 25780 5364 25832 5370
rect 25780 5306 25832 5312
rect 25596 5160 25648 5166
rect 25596 5102 25648 5108
rect 25884 4690 25912 11766
rect 26240 9920 26292 9926
rect 26240 9862 26292 9868
rect 26252 9654 26280 9862
rect 26344 9674 26372 12406
rect 26436 11218 26464 14418
rect 26516 12708 26568 12714
rect 26516 12650 26568 12656
rect 26528 11898 26556 12650
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 26436 10674 26464 11154
rect 26620 10690 26648 17614
rect 26712 16114 26740 17682
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26712 14498 26740 16050
rect 26804 14634 26832 37266
rect 27080 37262 27108 37402
rect 27068 37256 27120 37262
rect 27068 37198 27120 37204
rect 28724 37256 28776 37262
rect 28724 37198 28776 37204
rect 28736 23866 28764 37198
rect 29012 37126 29040 39200
rect 29000 37120 29052 37126
rect 30300 37108 30328 39200
rect 30472 37256 30524 37262
rect 30472 37198 30524 37204
rect 30380 37120 30432 37126
rect 30300 37080 30380 37108
rect 29000 37062 29052 37068
rect 30380 37062 30432 37068
rect 30484 36378 30512 37198
rect 32232 37126 32260 39200
rect 34164 37466 34192 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34152 37460 34204 37466
rect 34152 37402 34204 37408
rect 34796 37324 34848 37330
rect 34796 37266 34848 37272
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 32324 36922 32352 37198
rect 32312 36916 32364 36922
rect 32312 36858 32364 36864
rect 30472 36372 30524 36378
rect 30472 36314 30524 36320
rect 33692 30660 33744 30666
rect 33692 30602 33744 30608
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 28080 23724 28132 23730
rect 28080 23666 28132 23672
rect 28092 20262 28120 23666
rect 28080 20256 28132 20262
rect 28080 20198 28132 20204
rect 26884 19508 26936 19514
rect 26884 19450 26936 19456
rect 26896 17814 26924 19450
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 26884 17808 26936 17814
rect 26884 17750 26936 17756
rect 27172 17678 27200 18022
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 26976 16584 27028 16590
rect 26976 16526 27028 16532
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 26804 14606 26924 14634
rect 26712 14470 26832 14498
rect 26804 14346 26832 14470
rect 26700 14340 26752 14346
rect 26700 14282 26752 14288
rect 26792 14340 26844 14346
rect 26792 14282 26844 14288
rect 26712 13530 26740 14282
rect 26804 13938 26832 14282
rect 26792 13932 26844 13938
rect 26792 13874 26844 13880
rect 26896 13734 26924 14606
rect 26988 14278 27016 16526
rect 27068 16176 27120 16182
rect 27068 16118 27120 16124
rect 26976 14272 27028 14278
rect 26976 14214 27028 14220
rect 26884 13728 26936 13734
rect 26884 13670 26936 13676
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 26700 11620 26752 11626
rect 26700 11562 26752 11568
rect 26712 11082 26740 11562
rect 26792 11552 26844 11558
rect 26792 11494 26844 11500
rect 26804 11218 26832 11494
rect 26792 11212 26844 11218
rect 26792 11154 26844 11160
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26792 11076 26844 11082
rect 26792 11018 26844 11024
rect 26424 10668 26476 10674
rect 26620 10662 26740 10690
rect 26424 10610 26476 10616
rect 26608 10532 26660 10538
rect 26608 10474 26660 10480
rect 26620 10130 26648 10474
rect 26608 10124 26660 10130
rect 26608 10066 26660 10072
rect 26516 9988 26568 9994
rect 26516 9930 26568 9936
rect 26240 9648 26292 9654
rect 26344 9646 26464 9674
rect 26240 9590 26292 9596
rect 26332 9512 26384 9518
rect 26332 9454 26384 9460
rect 26344 9042 26372 9454
rect 26332 9036 26384 9042
rect 26332 8978 26384 8984
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 26068 4758 26096 8434
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 26160 6866 26188 7482
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 26240 6384 26292 6390
rect 26240 6326 26292 6332
rect 26056 4752 26108 4758
rect 26056 4694 26108 4700
rect 25872 4684 25924 4690
rect 25872 4626 25924 4632
rect 26148 4684 26200 4690
rect 26148 4626 26200 4632
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 24768 4004 24820 4010
rect 24768 3946 24820 3952
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 23664 3120 23716 3126
rect 23664 3062 23716 3068
rect 23676 2854 23704 3062
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 24596 2514 24624 3470
rect 24780 3466 24808 3946
rect 24950 3632 25006 3641
rect 24950 3567 24952 3576
rect 25004 3567 25006 3576
rect 24952 3538 25004 3544
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 25516 3126 25544 4082
rect 26160 3398 26188 4626
rect 26252 3942 26280 6326
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 26436 3754 26464 9646
rect 26528 8634 26556 9930
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26528 7818 26556 8026
rect 26516 7812 26568 7818
rect 26516 7754 26568 7760
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26620 5846 26648 7686
rect 26608 5840 26660 5846
rect 26608 5782 26660 5788
rect 26712 5794 26740 10662
rect 26804 9450 26832 11018
rect 26792 9444 26844 9450
rect 26792 9386 26844 9392
rect 26988 6662 27016 14214
rect 27080 14074 27108 16118
rect 27172 16114 27200 16526
rect 27344 16516 27396 16522
rect 27344 16458 27396 16464
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27068 14068 27120 14074
rect 27068 14010 27120 14016
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 27080 11150 27108 11698
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 27068 10192 27120 10198
rect 27068 10134 27120 10140
rect 27080 8634 27108 10134
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 26976 6656 27028 6662
rect 26976 6598 27028 6604
rect 26712 5766 26832 5794
rect 26700 5364 26752 5370
rect 26700 5306 26752 5312
rect 26712 4622 26740 5306
rect 26804 4826 26832 5766
rect 26988 5098 27016 6598
rect 27080 6390 27108 8570
rect 27172 6882 27200 16050
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 27264 15026 27292 15846
rect 27356 15162 27384 16458
rect 27448 15706 27476 17138
rect 27540 16590 27568 17138
rect 27528 16584 27580 16590
rect 27528 16526 27580 16532
rect 27528 16448 27580 16454
rect 27528 16390 27580 16396
rect 27436 15700 27488 15706
rect 27436 15642 27488 15648
rect 27540 15570 27568 16390
rect 27896 15904 27948 15910
rect 27896 15846 27948 15852
rect 27908 15570 27936 15846
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 27896 15564 27948 15570
rect 27896 15506 27948 15512
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27620 14952 27672 14958
rect 27620 14894 27672 14900
rect 27632 14482 27660 14894
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 27724 14550 27752 14758
rect 27712 14544 27764 14550
rect 27712 14486 27764 14492
rect 27620 14476 27672 14482
rect 27620 14418 27672 14424
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27252 13320 27304 13326
rect 27252 13262 27304 13268
rect 27264 12850 27292 13262
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27264 12434 27292 12786
rect 27264 12406 27384 12434
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27264 7886 27292 8774
rect 27252 7880 27304 7886
rect 27252 7822 27304 7828
rect 27252 7472 27304 7478
rect 27252 7414 27304 7420
rect 27264 7177 27292 7414
rect 27250 7168 27306 7177
rect 27250 7103 27306 7112
rect 27172 6866 27292 6882
rect 27160 6860 27292 6866
rect 27212 6854 27292 6860
rect 27160 6802 27212 6808
rect 27160 6724 27212 6730
rect 27160 6666 27212 6672
rect 27172 6458 27200 6666
rect 27160 6452 27212 6458
rect 27160 6394 27212 6400
rect 27068 6384 27120 6390
rect 27068 6326 27120 6332
rect 27264 5778 27292 6854
rect 27252 5772 27304 5778
rect 27252 5714 27304 5720
rect 26976 5092 27028 5098
rect 26976 5034 27028 5040
rect 26792 4820 26844 4826
rect 26844 4780 26924 4808
rect 26792 4762 26844 4768
rect 26700 4616 26752 4622
rect 26700 4558 26752 4564
rect 26436 3726 26556 3754
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26344 3194 26372 3334
rect 26332 3188 26384 3194
rect 26332 3130 26384 3136
rect 25228 3120 25280 3126
rect 24780 3058 24900 3074
rect 25228 3062 25280 3068
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 24780 3052 24912 3058
rect 24780 3046 24860 3052
rect 24780 2854 24808 3046
rect 24860 2994 24912 3000
rect 25240 2922 25268 3062
rect 25608 3058 25912 3074
rect 25596 3052 25924 3058
rect 25648 3046 25872 3052
rect 25596 2994 25648 3000
rect 25872 2994 25924 3000
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 25136 2848 25188 2854
rect 25136 2790 25188 2796
rect 23480 2508 23532 2514
rect 23480 2450 23532 2456
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24584 2372 24636 2378
rect 24584 2314 24636 2320
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 24596 2106 24624 2314
rect 24584 2100 24636 2106
rect 24584 2042 24636 2048
rect 25148 800 25176 2790
rect 26344 2650 26372 3130
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 26436 2514 26464 3538
rect 26528 3505 26556 3726
rect 26712 3584 26740 4558
rect 26792 3596 26844 3602
rect 26712 3556 26792 3584
rect 26792 3538 26844 3544
rect 26896 3505 26924 4780
rect 27356 4078 27384 12406
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27448 11082 27476 11698
rect 27436 11076 27488 11082
rect 27436 11018 27488 11024
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27448 7478 27476 8298
rect 27540 8106 27568 13874
rect 27908 12986 27936 14282
rect 27896 12980 27948 12986
rect 27896 12922 27948 12928
rect 27896 12776 27948 12782
rect 27896 12718 27948 12724
rect 27620 12640 27672 12646
rect 27620 12582 27672 12588
rect 27632 12306 27660 12582
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27908 12238 27936 12718
rect 27896 12232 27948 12238
rect 27896 12174 27948 12180
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 27540 8078 27660 8106
rect 27528 8016 27580 8022
rect 27528 7958 27580 7964
rect 27540 7818 27568 7958
rect 27528 7812 27580 7818
rect 27528 7754 27580 7760
rect 27632 7698 27660 8078
rect 27540 7670 27660 7698
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 27436 7472 27488 7478
rect 27436 7414 27488 7420
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27448 5370 27476 5646
rect 27436 5364 27488 5370
rect 27436 5306 27488 5312
rect 27540 5302 27568 7670
rect 27724 7274 27752 7686
rect 27712 7268 27764 7274
rect 27712 7210 27764 7216
rect 27816 7206 27844 10406
rect 27988 7336 28040 7342
rect 27988 7278 28040 7284
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 27816 6390 27844 7142
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 28000 6118 28028 7278
rect 27988 6112 28040 6118
rect 27988 6054 28040 6060
rect 27528 5296 27580 5302
rect 27528 5238 27580 5244
rect 27344 4072 27396 4078
rect 27344 4014 27396 4020
rect 27252 3936 27304 3942
rect 27252 3878 27304 3884
rect 27264 3602 27292 3878
rect 27252 3596 27304 3602
rect 27252 3538 27304 3544
rect 26514 3496 26570 3505
rect 26882 3496 26938 3505
rect 26514 3431 26570 3440
rect 26608 3460 26660 3466
rect 26528 2650 26556 3431
rect 26882 3431 26938 3440
rect 27160 3460 27212 3466
rect 26608 3402 26660 3408
rect 27160 3402 27212 3408
rect 26620 3194 26648 3402
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 27068 2916 27120 2922
rect 27068 2858 27120 2864
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 26424 2508 26476 2514
rect 26424 2450 26476 2456
rect 26252 1970 26280 2450
rect 26240 1964 26292 1970
rect 26240 1906 26292 1912
rect 27080 800 27108 2858
rect 27172 2514 27200 3402
rect 27264 3194 27292 3538
rect 27252 3188 27304 3194
rect 27252 3130 27304 3136
rect 27264 2922 27292 3130
rect 27252 2916 27304 2922
rect 27252 2858 27304 2864
rect 27356 2514 27384 4014
rect 28092 3194 28120 20198
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 33152 17882 33180 19314
rect 33140 17876 33192 17882
rect 33140 17818 33192 17824
rect 31208 17536 31260 17542
rect 31208 17478 31260 17484
rect 29368 15632 29420 15638
rect 29368 15574 29420 15580
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 28184 14958 28212 15302
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28172 14952 28224 14958
rect 28172 14894 28224 14900
rect 28448 14000 28500 14006
rect 28448 13942 28500 13948
rect 28460 12442 28488 13942
rect 28448 12436 28500 12442
rect 28552 12434 28580 14962
rect 29184 12912 29236 12918
rect 29184 12854 29236 12860
rect 28552 12406 28672 12434
rect 28448 12378 28500 12384
rect 28540 8900 28592 8906
rect 28540 8842 28592 8848
rect 28552 8566 28580 8842
rect 28540 8560 28592 8566
rect 28540 8502 28592 8508
rect 28448 7336 28500 7342
rect 28448 7278 28500 7284
rect 28460 6866 28488 7278
rect 28448 6860 28500 6866
rect 28448 6802 28500 6808
rect 28448 6724 28500 6730
rect 28368 6684 28448 6712
rect 28368 6390 28396 6684
rect 28448 6666 28500 6672
rect 28356 6384 28408 6390
rect 28356 6326 28408 6332
rect 28356 5364 28408 5370
rect 28356 5306 28408 5312
rect 28368 5234 28396 5306
rect 28356 5228 28408 5234
rect 28356 5170 28408 5176
rect 28368 4826 28396 5170
rect 28356 4820 28408 4826
rect 28356 4762 28408 4768
rect 28540 4752 28592 4758
rect 28540 4694 28592 4700
rect 28552 3233 28580 4694
rect 28644 3738 28672 12406
rect 29092 12164 29144 12170
rect 29092 12106 29144 12112
rect 29104 10674 29132 12106
rect 29092 10668 29144 10674
rect 29092 10610 29144 10616
rect 29092 10056 29144 10062
rect 29092 9998 29144 10004
rect 28816 8968 28868 8974
rect 28816 8910 28868 8916
rect 28828 8294 28856 8910
rect 29104 8566 29132 9998
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 28908 8424 28960 8430
rect 28960 8372 29040 8378
rect 28908 8366 29040 8372
rect 28920 8350 29040 8366
rect 28816 8288 28868 8294
rect 28816 8230 28868 8236
rect 28828 7002 28856 8230
rect 29012 7818 29040 8350
rect 29000 7812 29052 7818
rect 29000 7754 29052 7760
rect 29000 7472 29052 7478
rect 29000 7414 29052 7420
rect 29012 7342 29040 7414
rect 29000 7336 29052 7342
rect 29000 7278 29052 7284
rect 28906 7168 28962 7177
rect 28962 7126 29040 7154
rect 28906 7103 28962 7112
rect 28816 6996 28868 7002
rect 28816 6938 28868 6944
rect 28908 6996 28960 7002
rect 28908 6938 28960 6944
rect 28920 5658 28948 6938
rect 28736 5630 28948 5658
rect 28736 5574 28764 5630
rect 28724 5568 28776 5574
rect 28724 5510 28776 5516
rect 28908 5296 28960 5302
rect 28908 5238 28960 5244
rect 28920 5137 28948 5238
rect 28906 5128 28962 5137
rect 28906 5063 28962 5072
rect 29012 5030 29040 7126
rect 29104 5574 29132 8502
rect 29196 5846 29224 12854
rect 29380 8974 29408 15574
rect 30472 15564 30524 15570
rect 30472 15506 30524 15512
rect 30484 12434 30512 15506
rect 31220 12434 31248 17478
rect 30484 12406 30604 12434
rect 31220 12406 31340 12434
rect 29460 12232 29512 12238
rect 29460 12174 29512 12180
rect 29368 8968 29420 8974
rect 29368 8910 29420 8916
rect 29276 8832 29328 8838
rect 29276 8774 29328 8780
rect 29288 8498 29316 8774
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29288 7886 29316 8434
rect 29276 7880 29328 7886
rect 29276 7822 29328 7828
rect 29380 7206 29408 8910
rect 29368 7200 29420 7206
rect 29368 7142 29420 7148
rect 29184 5840 29236 5846
rect 29184 5782 29236 5788
rect 29092 5568 29144 5574
rect 29092 5510 29144 5516
rect 29092 5160 29144 5166
rect 29092 5102 29144 5108
rect 29000 5024 29052 5030
rect 29000 4966 29052 4972
rect 29104 4826 29132 5102
rect 29092 4820 29144 4826
rect 29092 4762 29144 4768
rect 29196 4554 29224 5782
rect 29276 5160 29328 5166
rect 29276 5102 29328 5108
rect 29288 4622 29316 5102
rect 29276 4616 29328 4622
rect 29276 4558 29328 4564
rect 29184 4548 29236 4554
rect 29184 4490 29236 4496
rect 28632 3732 28684 3738
rect 28632 3674 28684 3680
rect 29000 3664 29052 3670
rect 29052 3612 29132 3618
rect 29000 3606 29132 3612
rect 29012 3590 29132 3606
rect 29104 3584 29132 3590
rect 29276 3596 29328 3602
rect 29104 3556 29276 3584
rect 29276 3538 29328 3544
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 28724 3392 28776 3398
rect 28724 3334 28776 3340
rect 28538 3224 28594 3233
rect 28080 3188 28132 3194
rect 28538 3159 28594 3168
rect 28080 3130 28132 3136
rect 28736 2990 28764 3334
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 29012 2922 29040 3470
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 29000 2916 29052 2922
rect 29000 2858 29052 2864
rect 29012 2514 29040 2858
rect 27160 2508 27212 2514
rect 27160 2450 27212 2456
rect 27344 2508 27396 2514
rect 27344 2450 27396 2456
rect 29000 2508 29052 2514
rect 29000 2450 29052 2456
rect 28264 2372 28316 2378
rect 28264 2314 28316 2320
rect 28276 1902 28304 2314
rect 29104 2122 29132 3130
rect 29380 2650 29408 7142
rect 29472 5370 29500 12174
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 29564 8022 29592 10610
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 30012 8288 30064 8294
rect 30012 8230 30064 8236
rect 29552 8016 29604 8022
rect 29552 7958 29604 7964
rect 29564 7750 29592 7958
rect 30024 7954 30052 8230
rect 30012 7948 30064 7954
rect 30012 7890 30064 7896
rect 29552 7744 29604 7750
rect 29552 7686 29604 7692
rect 29644 7200 29696 7206
rect 29644 7142 29696 7148
rect 29656 6390 29684 7142
rect 30116 6866 30144 8434
rect 30196 7744 30248 7750
rect 30196 7686 30248 7692
rect 30104 6860 30156 6866
rect 30104 6802 30156 6808
rect 29736 6792 29788 6798
rect 29736 6734 29788 6740
rect 29748 6390 29776 6734
rect 30208 6662 30236 7686
rect 29920 6656 29972 6662
rect 29920 6598 29972 6604
rect 30196 6656 30248 6662
rect 30196 6598 30248 6604
rect 29644 6384 29696 6390
rect 29644 6326 29696 6332
rect 29736 6384 29788 6390
rect 29736 6326 29788 6332
rect 29932 6186 29960 6598
rect 30484 6390 30512 8842
rect 30472 6384 30524 6390
rect 30472 6326 30524 6332
rect 29920 6180 29972 6186
rect 29920 6122 29972 6128
rect 29460 5364 29512 5370
rect 29460 5306 29512 5312
rect 29920 5364 29972 5370
rect 29920 5306 29972 5312
rect 29932 4078 29960 5306
rect 30104 4684 30156 4690
rect 30104 4626 30156 4632
rect 30116 4128 30144 4626
rect 30196 4140 30248 4146
rect 30116 4100 30196 4128
rect 30196 4082 30248 4088
rect 29920 4072 29972 4078
rect 30288 4072 30340 4078
rect 29920 4014 29972 4020
rect 30116 4020 30288 4026
rect 30116 4014 30340 4020
rect 30116 3998 30328 4014
rect 30116 2854 30144 3998
rect 30196 3936 30248 3942
rect 30196 3878 30248 3884
rect 30208 3126 30236 3878
rect 30576 3602 30604 12406
rect 30932 8832 30984 8838
rect 30932 8774 30984 8780
rect 30944 8566 30972 8774
rect 30932 8560 30984 8566
rect 30932 8502 30984 8508
rect 31208 8424 31260 8430
rect 31208 8366 31260 8372
rect 31220 8090 31248 8366
rect 31208 8084 31260 8090
rect 31208 8026 31260 8032
rect 30748 7948 30800 7954
rect 30748 7890 30800 7896
rect 30654 7576 30710 7585
rect 30654 7511 30710 7520
rect 30668 7478 30696 7511
rect 30656 7472 30708 7478
rect 30656 7414 30708 7420
rect 30656 7336 30708 7342
rect 30656 7278 30708 7284
rect 30668 7206 30696 7278
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 30760 4826 30788 7890
rect 30944 6174 31156 6202
rect 30840 6112 30892 6118
rect 30944 6100 30972 6174
rect 31128 6118 31156 6174
rect 30892 6072 30972 6100
rect 31024 6112 31076 6118
rect 30840 6054 30892 6060
rect 31024 6054 31076 6060
rect 31116 6112 31168 6118
rect 31116 6054 31168 6060
rect 31036 5302 31064 6054
rect 31128 5794 31156 6054
rect 31128 5766 31248 5794
rect 31220 5642 31248 5766
rect 31116 5636 31168 5642
rect 31116 5578 31168 5584
rect 31208 5636 31260 5642
rect 31208 5578 31260 5584
rect 31024 5296 31076 5302
rect 31024 5238 31076 5244
rect 31022 5128 31078 5137
rect 31022 5063 31078 5072
rect 31036 4826 31064 5063
rect 30748 4820 30800 4826
rect 30748 4762 30800 4768
rect 31024 4820 31076 4826
rect 31024 4762 31076 4768
rect 31128 4758 31156 5578
rect 31116 4752 31168 4758
rect 31116 4694 31168 4700
rect 31312 4690 31340 12406
rect 31484 11144 31536 11150
rect 31484 11086 31536 11092
rect 31392 5568 31444 5574
rect 31392 5510 31444 5516
rect 31404 5098 31432 5510
rect 31392 5092 31444 5098
rect 31392 5034 31444 5040
rect 31300 4684 31352 4690
rect 31300 4626 31352 4632
rect 31114 4176 31170 4185
rect 30748 4140 30800 4146
rect 31114 4111 31116 4120
rect 30748 4082 30800 4088
rect 31168 4111 31170 4120
rect 31116 4082 31168 4088
rect 30564 3596 30616 3602
rect 30564 3538 30616 3544
rect 30196 3120 30248 3126
rect 30196 3062 30248 3068
rect 30380 2984 30432 2990
rect 30380 2926 30432 2932
rect 30472 2984 30524 2990
rect 30576 2972 30604 3538
rect 30760 3058 30788 4082
rect 31208 3936 31260 3942
rect 31208 3878 31260 3884
rect 31220 3602 31248 3878
rect 31312 3670 31340 4626
rect 31300 3664 31352 3670
rect 31300 3606 31352 3612
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 31206 3496 31262 3505
rect 31206 3431 31262 3440
rect 30748 3052 30800 3058
rect 30748 2994 30800 3000
rect 30524 2944 30604 2972
rect 31220 2961 31248 3431
rect 31392 3188 31444 3194
rect 31392 3130 31444 3136
rect 31206 2952 31262 2961
rect 30472 2926 30524 2932
rect 30104 2848 30156 2854
rect 30104 2790 30156 2796
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29012 2094 29132 2122
rect 28264 1896 28316 1902
rect 28264 1838 28316 1844
rect 29012 800 29040 2094
rect 30300 800 30328 2790
rect 30392 2774 30420 2926
rect 31404 2922 31432 3130
rect 31496 2990 31524 11086
rect 33600 10600 33652 10606
rect 33600 10542 33652 10548
rect 33612 10266 33640 10542
rect 33600 10260 33652 10266
rect 33600 10202 33652 10208
rect 32128 8288 32180 8294
rect 32128 8230 32180 8236
rect 31576 8016 31628 8022
rect 31576 7958 31628 7964
rect 31668 8016 31720 8022
rect 31668 7958 31720 7964
rect 31588 6662 31616 7958
rect 31680 7002 31708 7958
rect 32036 7812 32088 7818
rect 32036 7754 32088 7760
rect 31668 6996 31720 7002
rect 31668 6938 31720 6944
rect 32048 6798 32076 7754
rect 32036 6792 32088 6798
rect 32036 6734 32088 6740
rect 31944 6724 31996 6730
rect 31944 6666 31996 6672
rect 31576 6656 31628 6662
rect 31576 6598 31628 6604
rect 31956 6458 31984 6666
rect 31944 6452 31996 6458
rect 31944 6394 31996 6400
rect 31668 6112 31720 6118
rect 31668 6054 31720 6060
rect 32036 6112 32088 6118
rect 32036 6054 32088 6060
rect 31680 5778 31708 6054
rect 31668 5772 31720 5778
rect 31668 5714 31720 5720
rect 31668 5636 31720 5642
rect 31668 5578 31720 5584
rect 31680 3754 31708 5578
rect 31944 5024 31996 5030
rect 31944 4966 31996 4972
rect 31588 3726 31708 3754
rect 31588 3534 31616 3726
rect 31956 3534 31984 4966
rect 32048 4554 32076 6054
rect 32140 4826 32168 8230
rect 33140 7880 33192 7886
rect 33140 7822 33192 7828
rect 33152 7410 33180 7822
rect 33704 7546 33732 30602
rect 34808 16794 34836 37266
rect 36096 37126 36124 39200
rect 36268 37256 36320 37262
rect 36268 37198 36320 37204
rect 36912 37256 36964 37262
rect 36912 37198 36964 37204
rect 36084 37120 36136 37126
rect 36084 37062 36136 37068
rect 36280 36582 36308 37198
rect 36924 36718 36952 37198
rect 38028 37126 38056 39200
rect 38290 38176 38346 38185
rect 38290 38111 38346 38120
rect 38016 37120 38068 37126
rect 38016 37062 38068 37068
rect 36912 36712 36964 36718
rect 36912 36654 36964 36660
rect 36268 36576 36320 36582
rect 36268 36518 36320 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35716 22636 35768 22642
rect 35716 22578 35768 22584
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35728 14618 35756 22578
rect 35716 14612 35768 14618
rect 35716 14554 35768 14560
rect 35348 14408 35400 14414
rect 35348 14350 35400 14356
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 33692 7540 33744 7546
rect 33692 7482 33744 7488
rect 32220 7404 32272 7410
rect 32220 7346 32272 7352
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 32232 6798 32260 7346
rect 32220 6792 32272 6798
rect 32220 6734 32272 6740
rect 32232 6322 32260 6734
rect 32404 6656 32456 6662
rect 32404 6598 32456 6604
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 32232 5710 32260 6258
rect 32416 6254 32444 6598
rect 33152 6322 33180 7346
rect 33140 6316 33192 6322
rect 33140 6258 33192 6264
rect 32404 6248 32456 6254
rect 32404 6190 32456 6196
rect 32312 5772 32364 5778
rect 32312 5714 32364 5720
rect 32220 5704 32272 5710
rect 32220 5646 32272 5652
rect 32232 5574 32260 5646
rect 32220 5568 32272 5574
rect 32220 5510 32272 5516
rect 32128 4820 32180 4826
rect 32128 4762 32180 4768
rect 32036 4548 32088 4554
rect 32036 4490 32088 4496
rect 32220 3936 32272 3942
rect 32218 3904 32220 3913
rect 32272 3904 32274 3913
rect 32218 3839 32274 3848
rect 31576 3528 31628 3534
rect 31576 3470 31628 3476
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 31850 3224 31906 3233
rect 31850 3159 31906 3168
rect 31864 2990 31892 3159
rect 31956 3126 31984 3470
rect 31944 3120 31996 3126
rect 31944 3062 31996 3068
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 31852 2984 31904 2990
rect 31852 2926 31904 2932
rect 31206 2887 31262 2896
rect 31392 2916 31444 2922
rect 30392 2746 30696 2774
rect 30668 2650 30696 2746
rect 30656 2644 30708 2650
rect 30656 2586 30708 2592
rect 31220 2378 31248 2887
rect 31392 2858 31444 2864
rect 31956 2514 31984 3062
rect 32324 2854 32352 5714
rect 32864 5704 32916 5710
rect 32864 5646 32916 5652
rect 33152 5692 33180 6258
rect 33704 5846 33732 7482
rect 34060 7336 34112 7342
rect 34060 7278 34112 7284
rect 33692 5840 33744 5846
rect 33692 5782 33744 5788
rect 33232 5704 33284 5710
rect 33152 5664 33232 5692
rect 32876 5234 32904 5646
rect 33152 5302 33180 5664
rect 33232 5646 33284 5652
rect 33140 5296 33192 5302
rect 33140 5238 33192 5244
rect 32864 5228 32916 5234
rect 32864 5170 32916 5176
rect 32876 4622 32904 5170
rect 32864 4616 32916 4622
rect 32864 4558 32916 4564
rect 32876 4146 32904 4558
rect 33152 4554 33180 5238
rect 33784 5160 33836 5166
rect 33784 5102 33836 5108
rect 33796 4622 33824 5102
rect 34072 4826 34100 7278
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 34428 5704 34480 5710
rect 34428 5646 34480 5652
rect 34440 5234 34468 5646
rect 34428 5228 34480 5234
rect 34428 5170 34480 5176
rect 34520 5024 34572 5030
rect 34520 4966 34572 4972
rect 34060 4820 34112 4826
rect 34060 4762 34112 4768
rect 33784 4616 33836 4622
rect 33784 4558 33836 4564
rect 33140 4548 33192 4554
rect 33140 4490 33192 4496
rect 33416 4480 33468 4486
rect 33416 4422 33468 4428
rect 32954 4176 33010 4185
rect 32864 4140 32916 4146
rect 32954 4111 33010 4120
rect 32864 4082 32916 4088
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 32496 3936 32548 3942
rect 32496 3878 32548 3884
rect 32586 3904 32642 3913
rect 32416 3126 32444 3878
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32508 3058 32536 3878
rect 32586 3839 32642 3848
rect 32600 3602 32628 3839
rect 32588 3596 32640 3602
rect 32588 3538 32640 3544
rect 32496 3052 32548 3058
rect 32496 2994 32548 3000
rect 32312 2848 32364 2854
rect 32218 2816 32274 2825
rect 32312 2790 32364 2796
rect 32218 2751 32274 2760
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 31208 2372 31260 2378
rect 31208 2314 31260 2320
rect 32232 800 32260 2751
rect 32968 2446 32996 4111
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 32876 2106 32904 2246
rect 32864 2100 32916 2106
rect 32864 2042 32916 2048
rect 33428 1902 33456 4422
rect 33796 4185 33824 4558
rect 34428 4276 34480 4282
rect 34428 4218 34480 4224
rect 33782 4176 33838 4185
rect 33782 4111 33784 4120
rect 33836 4111 33838 4120
rect 34244 4140 34296 4146
rect 33784 4082 33836 4088
rect 34244 4082 34296 4088
rect 33692 3936 33744 3942
rect 33692 3878 33744 3884
rect 34152 3936 34204 3942
rect 34152 3878 34204 3884
rect 33704 1970 33732 3878
rect 34164 3194 34192 3878
rect 34256 3534 34284 4082
rect 34440 3738 34468 4218
rect 34428 3732 34480 3738
rect 34428 3674 34480 3680
rect 34532 3602 34560 4966
rect 34612 4548 34664 4554
rect 34612 4490 34664 4496
rect 34520 3596 34572 3602
rect 34520 3538 34572 3544
rect 34244 3528 34296 3534
rect 34244 3470 34296 3476
rect 34152 3188 34204 3194
rect 34152 3130 34204 3136
rect 34624 3126 34652 4490
rect 34612 3120 34664 3126
rect 34612 3062 34664 3068
rect 34244 2984 34296 2990
rect 34244 2926 34296 2932
rect 34256 2825 34284 2926
rect 34242 2816 34298 2825
rect 34242 2751 34298 2760
rect 34716 2446 34744 6598
rect 34796 6112 34848 6118
rect 34796 6054 34848 6060
rect 34808 5642 34836 6054
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34796 5636 34848 5642
rect 34796 5578 34848 5584
rect 34808 4468 34836 5578
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34888 4480 34940 4486
rect 34808 4440 34888 4468
rect 34888 4422 34940 4428
rect 34900 3942 34928 4422
rect 34888 3936 34940 3942
rect 34888 3878 34940 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34888 3528 34940 3534
rect 34888 3470 34940 3476
rect 34900 3058 34928 3470
rect 35360 3194 35388 14350
rect 36280 10810 36308 36518
rect 37740 36168 37792 36174
rect 37740 36110 37792 36116
rect 38198 36136 38254 36145
rect 37464 34536 37516 34542
rect 37464 34478 37516 34484
rect 37476 23866 37504 34478
rect 37464 23860 37516 23866
rect 37464 23802 37516 23808
rect 37280 19712 37332 19718
rect 37280 19654 37332 19660
rect 37292 15434 37320 19654
rect 37752 18970 37780 36110
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38304 35834 38332 38111
rect 39316 36922 39344 39200
rect 39304 36916 39356 36922
rect 39304 36858 39356 36864
rect 38292 35828 38344 35834
rect 38292 35770 38344 35776
rect 37924 35692 37976 35698
rect 37924 35634 37976 35640
rect 37936 20602 37964 35634
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 38212 34105 38240 34342
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38292 32360 38344 32366
rect 38292 32302 38344 32308
rect 38304 32065 38332 32302
rect 38290 32056 38346 32065
rect 38290 31991 38292 32000
rect 38344 31991 38346 32000
rect 38292 31962 38344 31968
rect 38292 30184 38344 30190
rect 38292 30126 38344 30132
rect 38304 30025 38332 30126
rect 38290 30016 38346 30025
rect 38290 29951 38346 29960
rect 38304 29850 38332 29951
rect 38292 29844 38344 29850
rect 38292 29786 38344 29792
rect 38016 29164 38068 29170
rect 38016 29106 38068 29112
rect 38028 28422 38056 29106
rect 38200 29028 38252 29034
rect 38200 28970 38252 28976
rect 38212 28665 38240 28970
rect 38198 28656 38254 28665
rect 38198 28591 38254 28600
rect 38016 28416 38068 28422
rect 38016 28358 38068 28364
rect 38016 26920 38068 26926
rect 38016 26862 38068 26868
rect 38292 26920 38344 26926
rect 38292 26862 38344 26868
rect 37924 20596 37976 20602
rect 37924 20538 37976 20544
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37844 19718 37872 20402
rect 37832 19712 37884 19718
rect 37832 19654 37884 19660
rect 38028 19530 38056 26862
rect 38304 26625 38332 26862
rect 38290 26616 38346 26625
rect 38290 26551 38292 26560
rect 38344 26551 38346 26560
rect 38292 26522 38344 26528
rect 38200 24812 38252 24818
rect 38200 24754 38252 24760
rect 38212 24585 38240 24754
rect 38198 24576 38254 24585
rect 38198 24511 38254 24520
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38200 20800 38252 20806
rect 38200 20742 38252 20748
rect 38212 20505 38240 20742
rect 38198 20496 38254 20505
rect 38198 20431 38254 20440
rect 37844 19502 38056 19530
rect 37740 18964 37792 18970
rect 37740 18906 37792 18912
rect 37844 16250 37872 19502
rect 38200 19168 38252 19174
rect 38198 19136 38200 19145
rect 38252 19136 38254 19145
rect 38198 19071 38254 19080
rect 38108 18760 38160 18766
rect 38108 18702 38160 18708
rect 38120 18086 38148 18702
rect 38108 18080 38160 18086
rect 38108 18022 38160 18028
rect 37924 16992 37976 16998
rect 37924 16934 37976 16940
rect 37832 16244 37884 16250
rect 37832 16186 37884 16192
rect 37280 15428 37332 15434
rect 37280 15370 37332 15376
rect 36268 10804 36320 10810
rect 36268 10746 36320 10752
rect 36176 10668 36228 10674
rect 36176 10610 36228 10616
rect 36188 10062 36216 10610
rect 36176 10056 36228 10062
rect 36176 9998 36228 10004
rect 35532 6112 35584 6118
rect 35532 6054 35584 6060
rect 36084 6112 36136 6118
rect 36084 6054 36136 6060
rect 35544 5574 35572 6054
rect 35532 5568 35584 5574
rect 35532 5510 35584 5516
rect 35544 5302 35572 5510
rect 35532 5296 35584 5302
rect 35532 5238 35584 5244
rect 35544 4282 35572 5238
rect 35992 4480 36044 4486
rect 35992 4422 36044 4428
rect 35532 4276 35584 4282
rect 35532 4218 35584 4224
rect 35532 3936 35584 3942
rect 35532 3878 35584 3884
rect 35544 3738 35572 3878
rect 35532 3732 35584 3738
rect 35532 3674 35584 3680
rect 35544 3194 35572 3674
rect 36004 3670 36032 4422
rect 35992 3664 36044 3670
rect 35992 3606 36044 3612
rect 35348 3188 35400 3194
rect 35348 3130 35400 3136
rect 35532 3188 35584 3194
rect 35532 3130 35584 3136
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35544 2650 35572 3130
rect 35532 2644 35584 2650
rect 35532 2586 35584 2592
rect 36096 2446 36124 6054
rect 36188 5914 36216 9998
rect 36176 5908 36228 5914
rect 36176 5850 36228 5856
rect 36452 5296 36504 5302
rect 36452 5238 36504 5244
rect 36464 4826 36492 5238
rect 36544 5024 36596 5030
rect 36544 4966 36596 4972
rect 36452 4820 36504 4826
rect 36452 4762 36504 4768
rect 36556 3058 36584 4966
rect 37188 3936 37240 3942
rect 37188 3878 37240 3884
rect 36636 3392 36688 3398
rect 36636 3334 36688 3340
rect 36544 3052 36596 3058
rect 36544 2994 36596 3000
rect 36648 2961 36676 3334
rect 36634 2952 36690 2961
rect 36634 2887 36690 2896
rect 34428 2440 34480 2446
rect 34428 2382 34480 2388
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 33692 1964 33744 1970
rect 33692 1906 33744 1912
rect 33416 1896 33468 1902
rect 33416 1838 33468 1844
rect 34164 870 34284 898
rect 34164 800 34192 870
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 5170 200 5226 800
rect 7102 200 7158 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 12254 200 12310 800
rect 14186 200 14242 800
rect 16118 200 16174 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 23202 200 23258 800
rect 25134 200 25190 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 34256 762 34284 870
rect 34440 762 34468 2382
rect 34980 2304 35032 2310
rect 34980 2246 35032 2252
rect 34992 2038 35020 2246
rect 34980 2032 35032 2038
rect 34980 1974 35032 1980
rect 36096 800 36124 2382
rect 37200 1465 37228 3878
rect 37292 2582 37320 15370
rect 37740 14272 37792 14278
rect 37740 14214 37792 14220
rect 37752 13938 37780 14214
rect 37740 13932 37792 13938
rect 37740 13874 37792 13880
rect 37752 12646 37780 13874
rect 37740 12640 37792 12646
rect 37740 12582 37792 12588
rect 37464 6112 37516 6118
rect 37464 6054 37516 6060
rect 37280 2576 37332 2582
rect 37280 2518 37332 2524
rect 37476 2514 37504 6054
rect 37752 2514 37780 12582
rect 37832 9172 37884 9178
rect 37832 9114 37884 9120
rect 37844 7954 37872 9114
rect 37832 7948 37884 7954
rect 37832 7890 37884 7896
rect 37844 4622 37872 7890
rect 37936 6866 37964 16934
rect 38016 15496 38068 15502
rect 38016 15438 38068 15444
rect 38028 14074 38056 15438
rect 38016 14068 38068 14074
rect 38016 14010 38068 14016
rect 38016 13320 38068 13326
rect 38016 13262 38068 13268
rect 38028 11626 38056 13262
rect 38016 11620 38068 11626
rect 38016 11562 38068 11568
rect 38120 11082 38148 18022
rect 38292 17196 38344 17202
rect 38292 17138 38344 17144
rect 38304 17105 38332 17138
rect 38290 17096 38346 17105
rect 38290 17031 38346 17040
rect 38200 15360 38252 15366
rect 38200 15302 38252 15308
rect 38212 15065 38240 15302
rect 38198 15056 38254 15065
rect 38198 14991 38254 15000
rect 38200 13184 38252 13190
rect 38200 13126 38252 13132
rect 38212 13025 38240 13126
rect 38198 13016 38254 13025
rect 38198 12951 38254 12960
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38108 11076 38160 11082
rect 38108 11018 38160 11024
rect 38120 9178 38148 11018
rect 38304 10985 38332 11086
rect 38290 10976 38346 10985
rect 38290 10911 38346 10920
rect 38304 10810 38332 10911
rect 38292 10804 38344 10810
rect 38292 10746 38344 10752
rect 38108 9172 38160 9178
rect 38108 9114 38160 9120
rect 38198 8936 38254 8945
rect 38198 8871 38200 8880
rect 38252 8871 38254 8880
rect 38200 8842 38252 8848
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38304 7585 38332 7822
rect 38290 7576 38346 7585
rect 38290 7511 38292 7520
rect 38344 7511 38346 7520
rect 38292 7482 38344 7488
rect 37924 6860 37976 6866
rect 37924 6802 37976 6808
rect 38200 6112 38252 6118
rect 38200 6054 38252 6060
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 38016 4480 38068 4486
rect 38016 4422 38068 4428
rect 38028 4146 38056 4422
rect 38016 4140 38068 4146
rect 38016 4082 38068 4088
rect 38014 3088 38070 3097
rect 38212 3058 38240 6054
rect 38292 5704 38344 5710
rect 38292 5646 38344 5652
rect 38304 5545 38332 5646
rect 38290 5536 38346 5545
rect 38290 5471 38346 5480
rect 38292 5024 38344 5030
rect 38292 4966 38344 4972
rect 38304 3534 38332 4966
rect 38292 3528 38344 3534
rect 38290 3496 38292 3505
rect 38344 3496 38346 3505
rect 38290 3431 38346 3440
rect 38014 3023 38016 3032
rect 38068 3023 38070 3032
rect 38200 3052 38252 3058
rect 38016 2994 38068 3000
rect 38200 2994 38252 3000
rect 39304 3052 39356 3058
rect 39304 2994 39356 3000
rect 37464 2508 37516 2514
rect 37464 2450 37516 2456
rect 37740 2508 37792 2514
rect 37740 2450 37792 2456
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 38028 800 38056 2382
rect 39316 800 39344 2994
rect 34256 734 34468 762
rect 36082 200 36138 800
rect 38014 200 38070 800
rect 39302 200 39358 800
<< via2 >>
rect 2778 38120 2834 38176
rect 1674 36080 1730 36136
rect 1674 34040 1730 34096
rect 1582 32020 1638 32056
rect 1582 32000 1584 32020
rect 1584 32000 1636 32020
rect 1636 32000 1638 32020
rect 1674 30640 1730 30696
rect 1674 28600 1730 28656
rect 1582 26580 1638 26616
rect 1582 26560 1584 26580
rect 1584 26560 1636 26580
rect 1636 26560 1638 26580
rect 1674 24556 1676 24576
rect 1676 24556 1728 24576
rect 1728 24556 1730 24576
rect 1674 24520 1730 24556
rect 1674 22480 1730 22536
rect 1582 20476 1584 20496
rect 1584 20476 1636 20496
rect 1636 20476 1638 20496
rect 1582 20440 1638 20476
rect 1582 19080 1638 19136
rect 1674 17060 1730 17096
rect 1674 17040 1676 17060
rect 1676 17040 1728 17060
rect 1728 17040 1730 17060
rect 1674 15000 1730 15056
rect 1674 12960 1730 13016
rect 1674 10956 1676 10976
rect 1676 10956 1728 10976
rect 1728 10956 1730 10976
rect 1674 10920 1730 10956
rect 1582 9596 1584 9616
rect 1584 9596 1636 9616
rect 1636 9596 1638 9616
rect 1582 9560 1638 9596
rect 1674 7520 1730 7576
rect 1674 5516 1676 5536
rect 1676 5516 1728 5536
rect 1728 5516 1730 5536
rect 1674 5480 1730 5516
rect 1674 3440 1730 3496
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 1582 1400 1638 1456
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 21362 10668 21418 10704
rect 21362 10648 21364 10668
rect 21364 10648 21416 10668
rect 21416 10648 21418 10668
rect 21454 3052 21510 3088
rect 21454 3032 21456 3052
rect 21456 3032 21508 3052
rect 21508 3032 21510 3052
rect 22190 10684 22192 10704
rect 22192 10684 22244 10704
rect 22244 10684 22246 10704
rect 22190 10648 22246 10684
rect 22834 3576 22890 3632
rect 22650 3460 22706 3496
rect 22650 3440 22652 3460
rect 22652 3440 22704 3460
rect 22704 3440 22706 3460
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 26330 23568 26386 23624
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 24950 3596 25006 3632
rect 24950 3576 24952 3596
rect 24952 3576 25004 3596
rect 25004 3576 25006 3596
rect 27250 7112 27306 7168
rect 26514 3440 26570 3496
rect 26882 3440 26938 3496
rect 28906 7112 28962 7168
rect 28906 5072 28962 5128
rect 28538 3168 28594 3224
rect 30654 7520 30710 7576
rect 31022 5072 31078 5128
rect 31114 4140 31170 4176
rect 31114 4120 31116 4140
rect 31116 4120 31168 4140
rect 31168 4120 31170 4140
rect 31206 3440 31262 3496
rect 31206 2896 31262 2952
rect 38290 38120 38346 38176
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 32218 3884 32220 3904
rect 32220 3884 32272 3904
rect 32272 3884 32274 3904
rect 32218 3848 32274 3884
rect 31850 3168 31906 3224
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 32954 4120 33010 4176
rect 32586 3848 32642 3904
rect 32218 2760 32274 2816
rect 33782 4140 33838 4176
rect 33782 4120 33784 4140
rect 33784 4120 33836 4140
rect 33836 4120 33838 4140
rect 34242 2760 34298 2816
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38198 36080 38254 36136
rect 38198 34040 38254 34096
rect 38290 32020 38346 32056
rect 38290 32000 38292 32020
rect 38292 32000 38344 32020
rect 38344 32000 38346 32020
rect 38290 29960 38346 30016
rect 38198 28600 38254 28656
rect 38290 26580 38346 26616
rect 38290 26560 38292 26580
rect 38292 26560 38344 26580
rect 38344 26560 38346 26580
rect 38198 24520 38254 24576
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38198 20440 38254 20496
rect 38198 19116 38200 19136
rect 38200 19116 38252 19136
rect 38252 19116 38254 19136
rect 38198 19080 38254 19116
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36634 2896 36690 2952
rect 38290 17040 38346 17096
rect 38198 15000 38254 15056
rect 38198 12960 38254 13016
rect 38290 10920 38346 10976
rect 38198 8900 38254 8936
rect 38198 8880 38200 8900
rect 38200 8880 38252 8900
rect 38252 8880 38254 8900
rect 38290 7540 38346 7576
rect 38290 7520 38292 7540
rect 38292 7520 38344 7540
rect 38344 7520 38346 7540
rect 38014 3052 38070 3088
rect 38290 5480 38346 5536
rect 38290 3476 38292 3496
rect 38292 3476 38344 3496
rect 38344 3476 38346 3496
rect 38290 3440 38346 3476
rect 38014 3032 38016 3052
rect 38016 3032 38068 3052
rect 38068 3032 38070 3052
rect 37186 1400 37242 1456
<< metal3 >>
rect 200 38178 800 38208
rect 2773 38178 2839 38181
rect 200 38176 2839 38178
rect 200 38120 2778 38176
rect 2834 38120 2839 38176
rect 200 38118 2839 38120
rect 200 38088 800 38118
rect 2773 38115 2839 38118
rect 38285 38178 38351 38181
rect 39200 38178 39800 38208
rect 38285 38176 39800 38178
rect 38285 38120 38290 38176
rect 38346 38120 39800 38176
rect 38285 38118 39800 38120
rect 38285 38115 38351 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1669 36138 1735 36141
rect 200 36136 1735 36138
rect 200 36080 1674 36136
rect 1730 36080 1735 36136
rect 200 36078 1735 36080
rect 200 36048 800 36078
rect 1669 36075 1735 36078
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1669 34098 1735 34101
rect 200 34096 1735 34098
rect 200 34040 1674 34096
rect 1730 34040 1735 34096
rect 200 34038 1735 34040
rect 200 34008 800 34038
rect 1669 34035 1735 34038
rect 38193 34098 38259 34101
rect 39200 34098 39800 34128
rect 38193 34096 39800 34098
rect 38193 34040 38198 34096
rect 38254 34040 39800 34096
rect 38193 34038 39800 34040
rect 38193 34035 38259 34038
rect 39200 34008 39800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1577 32058 1643 32061
rect 200 32056 1643 32058
rect 200 32000 1582 32056
rect 1638 32000 1643 32056
rect 200 31998 1643 32000
rect 200 31968 800 31998
rect 1577 31995 1643 31998
rect 38285 32058 38351 32061
rect 39200 32058 39800 32088
rect 38285 32056 39800 32058
rect 38285 32000 38290 32056
rect 38346 32000 39800 32056
rect 38285 31998 39800 32000
rect 38285 31995 38351 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1669 30698 1735 30701
rect 200 30696 1735 30698
rect 200 30640 1674 30696
rect 1730 30640 1735 30696
rect 200 30638 1735 30640
rect 200 30608 800 30638
rect 1669 30635 1735 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38285 30018 38351 30021
rect 39200 30018 39800 30048
rect 38285 30016 39800 30018
rect 38285 29960 38290 30016
rect 38346 29960 39800 30016
rect 38285 29958 39800 29960
rect 38285 29955 38351 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1669 28658 1735 28661
rect 200 28656 1735 28658
rect 200 28600 1674 28656
rect 1730 28600 1735 28656
rect 200 28598 1735 28600
rect 200 28568 800 28598
rect 1669 28595 1735 28598
rect 38193 28658 38259 28661
rect 39200 28658 39800 28688
rect 38193 28656 39800 28658
rect 38193 28600 38198 28656
rect 38254 28600 39800 28656
rect 38193 28598 39800 28600
rect 38193 28595 38259 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1577 26618 1643 26621
rect 200 26616 1643 26618
rect 200 26560 1582 26616
rect 1638 26560 1643 26616
rect 200 26558 1643 26560
rect 200 26528 800 26558
rect 1577 26555 1643 26558
rect 38285 26618 38351 26621
rect 39200 26618 39800 26648
rect 38285 26616 39800 26618
rect 38285 26560 38290 26616
rect 38346 26560 39800 26616
rect 38285 26558 39800 26560
rect 38285 26555 38351 26558
rect 39200 26528 39800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 200 24578 800 24608
rect 1669 24578 1735 24581
rect 200 24576 1735 24578
rect 200 24520 1674 24576
rect 1730 24520 1735 24576
rect 200 24518 1735 24520
rect 200 24488 800 24518
rect 1669 24515 1735 24518
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 26325 23628 26391 23629
rect 26325 23626 26372 23628
rect 26280 23624 26372 23626
rect 26280 23568 26330 23624
rect 26280 23566 26372 23568
rect 26325 23564 26372 23566
rect 26436 23564 26442 23628
rect 26325 23563 26391 23564
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1669 22538 1735 22541
rect 200 22536 1735 22538
rect 200 22480 1674 22536
rect 1730 22480 1735 22536
rect 200 22478 1735 22480
rect 200 22448 800 22478
rect 1669 22475 1735 22478
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1577 20498 1643 20501
rect 200 20496 1643 20498
rect 200 20440 1582 20496
rect 1638 20440 1643 20496
rect 200 20438 1643 20440
rect 200 20408 800 20438
rect 1577 20435 1643 20438
rect 38193 20498 38259 20501
rect 39200 20498 39800 20528
rect 38193 20496 39800 20498
rect 38193 20440 38198 20496
rect 38254 20440 39800 20496
rect 38193 20438 39800 20440
rect 38193 20435 38259 20438
rect 39200 20408 39800 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 19138 800 19168
rect 1577 19138 1643 19141
rect 200 19136 1643 19138
rect 200 19080 1582 19136
rect 1638 19080 1643 19136
rect 200 19078 1643 19080
rect 200 19048 800 19078
rect 1577 19075 1643 19078
rect 38193 19138 38259 19141
rect 39200 19138 39800 19168
rect 38193 19136 39800 19138
rect 38193 19080 38198 19136
rect 38254 19080 39800 19136
rect 38193 19078 39800 19080
rect 38193 19075 38259 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 200 17098 800 17128
rect 1669 17098 1735 17101
rect 200 17096 1735 17098
rect 200 17040 1674 17096
rect 1730 17040 1735 17096
rect 200 17038 1735 17040
rect 200 17008 800 17038
rect 1669 17035 1735 17038
rect 38285 17098 38351 17101
rect 39200 17098 39800 17128
rect 38285 17096 39800 17098
rect 38285 17040 38290 17096
rect 38346 17040 39800 17096
rect 38285 17038 39800 17040
rect 38285 17035 38351 17038
rect 39200 17008 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 200 15058 800 15088
rect 1669 15058 1735 15061
rect 200 15056 1735 15058
rect 200 15000 1674 15056
rect 1730 15000 1735 15056
rect 200 14998 1735 15000
rect 200 14968 800 14998
rect 1669 14995 1735 14998
rect 38193 15058 38259 15061
rect 39200 15058 39800 15088
rect 38193 15056 39800 15058
rect 38193 15000 38198 15056
rect 38254 15000 39800 15056
rect 38193 14998 39800 15000
rect 38193 14995 38259 14998
rect 39200 14968 39800 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 200 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 1669 13018 1735 13021
rect 200 13016 1735 13018
rect 200 12960 1674 13016
rect 1730 12960 1735 13016
rect 200 12958 1735 12960
rect 200 12928 800 12958
rect 1669 12955 1735 12958
rect 38193 13018 38259 13021
rect 39200 13018 39800 13048
rect 38193 13016 39800 13018
rect 38193 12960 38198 13016
rect 38254 12960 39800 13016
rect 38193 12958 39800 12960
rect 38193 12955 38259 12958
rect 39200 12928 39800 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 200 10978 800 11008
rect 1669 10978 1735 10981
rect 200 10976 1735 10978
rect 200 10920 1674 10976
rect 1730 10920 1735 10976
rect 200 10918 1735 10920
rect 200 10888 800 10918
rect 1669 10915 1735 10918
rect 38285 10978 38351 10981
rect 39200 10978 39800 11008
rect 38285 10976 39800 10978
rect 38285 10920 38290 10976
rect 38346 10920 39800 10976
rect 38285 10918 39800 10920
rect 38285 10915 38351 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 21357 10706 21423 10709
rect 22185 10706 22251 10709
rect 21357 10704 22251 10706
rect 21357 10648 21362 10704
rect 21418 10648 22190 10704
rect 22246 10648 22251 10704
rect 21357 10646 22251 10648
rect 21357 10643 21423 10646
rect 22185 10643 22251 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9648
rect 1577 9618 1643 9621
rect 200 9616 1643 9618
rect 200 9560 1582 9616
rect 1638 9560 1643 9616
rect 200 9558 1643 9560
rect 200 9528 800 9558
rect 1577 9555 1643 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1669 7578 1735 7581
rect 200 7576 1735 7578
rect 200 7520 1674 7576
rect 1730 7520 1735 7576
rect 200 7518 1735 7520
rect 200 7488 800 7518
rect 1669 7515 1735 7518
rect 26366 7516 26372 7580
rect 26436 7578 26442 7580
rect 30649 7578 30715 7581
rect 26436 7576 30715 7578
rect 26436 7520 30654 7576
rect 30710 7520 30715 7576
rect 26436 7518 30715 7520
rect 26436 7516 26442 7518
rect 30649 7515 30715 7518
rect 38285 7578 38351 7581
rect 39200 7578 39800 7608
rect 38285 7576 39800 7578
rect 38285 7520 38290 7576
rect 38346 7520 39800 7576
rect 38285 7518 39800 7520
rect 38285 7515 38351 7518
rect 39200 7488 39800 7518
rect 27245 7170 27311 7173
rect 28901 7170 28967 7173
rect 27245 7168 28967 7170
rect 27245 7112 27250 7168
rect 27306 7112 28906 7168
rect 28962 7112 28967 7168
rect 27245 7110 28967 7112
rect 27245 7107 27311 7110
rect 28901 7107 28967 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5538 800 5568
rect 1669 5538 1735 5541
rect 200 5536 1735 5538
rect 200 5480 1674 5536
rect 1730 5480 1735 5536
rect 200 5478 1735 5480
rect 200 5448 800 5478
rect 1669 5475 1735 5478
rect 38285 5538 38351 5541
rect 39200 5538 39800 5568
rect 38285 5536 39800 5538
rect 38285 5480 38290 5536
rect 38346 5480 39800 5536
rect 38285 5478 39800 5480
rect 38285 5475 38351 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 28901 5130 28967 5133
rect 31017 5130 31083 5133
rect 28901 5128 31083 5130
rect 28901 5072 28906 5128
rect 28962 5072 31022 5128
rect 31078 5072 31083 5128
rect 28901 5070 31083 5072
rect 28901 5067 28967 5070
rect 31017 5067 31083 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 31109 4178 31175 4181
rect 32949 4178 33015 4181
rect 33777 4178 33843 4181
rect 31109 4176 33843 4178
rect 31109 4120 31114 4176
rect 31170 4120 32954 4176
rect 33010 4120 33782 4176
rect 33838 4120 33843 4176
rect 31109 4118 33843 4120
rect 31109 4115 31175 4118
rect 32949 4115 33015 4118
rect 33777 4115 33843 4118
rect 32213 3906 32279 3909
rect 32581 3906 32647 3909
rect 32213 3904 32647 3906
rect 32213 3848 32218 3904
rect 32274 3848 32586 3904
rect 32642 3848 32647 3904
rect 32213 3846 32647 3848
rect 32213 3843 32279 3846
rect 32581 3843 32647 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 22829 3634 22895 3637
rect 24945 3634 25011 3637
rect 22829 3632 25011 3634
rect 22829 3576 22834 3632
rect 22890 3576 24950 3632
rect 25006 3576 25011 3632
rect 22829 3574 25011 3576
rect 22829 3571 22895 3574
rect 24945 3571 25011 3574
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 22645 3498 22711 3501
rect 26509 3498 26575 3501
rect 22645 3496 26575 3498
rect 22645 3440 22650 3496
rect 22706 3440 26514 3496
rect 26570 3440 26575 3496
rect 22645 3438 26575 3440
rect 22645 3435 22711 3438
rect 26509 3435 26575 3438
rect 26877 3498 26943 3501
rect 31201 3498 31267 3501
rect 26877 3496 31267 3498
rect 26877 3440 26882 3496
rect 26938 3440 31206 3496
rect 31262 3440 31267 3496
rect 26877 3438 31267 3440
rect 26877 3435 26943 3438
rect 31201 3435 31267 3438
rect 38285 3498 38351 3501
rect 39200 3498 39800 3528
rect 38285 3496 39800 3498
rect 38285 3440 38290 3496
rect 38346 3440 39800 3496
rect 38285 3438 39800 3440
rect 38285 3435 38351 3438
rect 39200 3408 39800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 28533 3226 28599 3229
rect 31845 3226 31911 3229
rect 28533 3224 31911 3226
rect 28533 3168 28538 3224
rect 28594 3168 31850 3224
rect 31906 3168 31911 3224
rect 28533 3166 31911 3168
rect 28533 3163 28599 3166
rect 31845 3163 31911 3166
rect 21449 3090 21515 3093
rect 38009 3090 38075 3093
rect 21449 3088 38075 3090
rect 21449 3032 21454 3088
rect 21510 3032 38014 3088
rect 38070 3032 38075 3088
rect 21449 3030 38075 3032
rect 21449 3027 21515 3030
rect 38009 3027 38075 3030
rect 31201 2954 31267 2957
rect 36629 2954 36695 2957
rect 31201 2952 36695 2954
rect 31201 2896 31206 2952
rect 31262 2896 36634 2952
rect 36690 2896 36695 2952
rect 31201 2894 36695 2896
rect 31201 2891 31267 2894
rect 36629 2891 36695 2894
rect 32213 2818 32279 2821
rect 34237 2818 34303 2821
rect 32213 2816 34303 2818
rect 32213 2760 32218 2816
rect 32274 2760 34242 2816
rect 34298 2760 34303 2816
rect 32213 2758 34303 2760
rect 32213 2755 32279 2758
rect 34237 2755 34303 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 1577 1458 1643 1461
rect 200 1456 1643 1458
rect 200 1400 1582 1456
rect 1638 1400 1643 1456
rect 200 1398 1643 1400
rect 200 1368 800 1398
rect 1577 1395 1643 1398
rect 37181 1458 37247 1461
rect 39200 1458 39800 1488
rect 37181 1456 39800 1458
rect 37181 1400 37186 1456
rect 37242 1400 39800 1456
rect 37181 1398 39800 1400
rect 37181 1395 37247 1398
rect 39200 1368 39800 1398
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 26372 23624 26436 23628
rect 26372 23568 26386 23624
rect 26386 23568 26436 23624
rect 26372 23564 26436 23568
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 26372 7516 26436 7580
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 26371 23628 26437 23629
rect 26371 23564 26372 23628
rect 26436 23564 26437 23628
rect 26371 23563 26437 23564
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 26374 7581 26434 23563
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 26371 7580 26437 7581
rect 26371 7516 26372 7580
rect 26436 7516 26437 7580
rect 26371 7515 26437 7516
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 27324 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1667941163
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1667941163
transform -1 0 25760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1667941163
transform 1 0 25944 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A
timestamp 1667941163
transform 1 0 27140 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1667941163
transform 1 0 22632 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1667941163
transform 1 0 23920 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1667941163
transform -1 0 21896 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1667941163
transform -1 0 22080 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1667941163
transform -1 0 28612 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1667941163
transform -1 0 27232 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1667941163
transform -1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1667941163
transform 1 0 20792 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1667941163
transform 1 0 21344 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1667941163
transform -1 0 27968 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1667941163
transform -1 0 26680 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1667941163
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1667941163
transform -1 0 28244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1667941163
transform -1 0 27784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1667941163
transform -1 0 20700 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1667941163
transform -1 0 21252 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1667941163
transform -1 0 21252 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 1667941163
transform 1 0 17756 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1667941163
transform 1 0 20056 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1667941163
transform 1 0 20976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1667941163
transform -1 0 17940 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A
timestamp 1667941163
transform 1 0 29072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1667941163
transform -1 0 19964 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1667941163
transform -1 0 24932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1667941163
transform -1 0 26312 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1667941163
transform 1 0 28060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A
timestamp 1667941163
transform -1 0 23552 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1667941163
transform 1 0 28704 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 1667941163
transform 1 0 27324 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1667941163
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A
timestamp 1667941163
transform -1 0 22448 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1667941163
transform -1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A
timestamp 1667941163
transform -1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1667941163
transform -1 0 12880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A
timestamp 1667941163
transform -1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1667941163
transform -1 0 30820 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1667941163
transform -1 0 17388 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1667941163
transform 1 0 27784 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 1667941163
transform -1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1667941163
transform 1 0 4048 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A
timestamp 1667941163
transform -1 0 23184 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1667941163
transform -1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1667941163
transform 1 0 25944 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1667941163
transform 1 0 23092 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1667941163
transform -1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1667941163
transform -1 0 22264 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1667941163
transform 1 0 27876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1667941163
transform -1 0 10948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1667941163
transform 1 0 35512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1667941163
transform 1 0 35880 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1667941163
transform 1 0 36064 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1667941163
transform -1 0 36708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1667941163
transform 1 0 36432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1667941163
transform 1 0 35328 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A
timestamp 1667941163
transform 1 0 33580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1667941163
transform -1 0 36156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__CLK
timestamp 1667941163
transform -1 0 29900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__CLK
timestamp 1667941163
transform 1 0 29072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__CLK
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__CLK
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__CLK
timestamp 1667941163
transform 1 0 28520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__D
timestamp 1667941163
transform 1 0 27508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__CLK
timestamp 1667941163
transform 1 0 27692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__D
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__CLK
timestamp 1667941163
transform 1 0 32292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__CLK
timestamp 1667941163
transform 1 0 35420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__CLK
timestamp 1667941163
transform 1 0 26496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__CLK
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__CLK
timestamp 1667941163
transform 1 0 25668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__CLK
timestamp 1667941163
transform 1 0 30360 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__CLK
timestamp 1667941163
transform 1 0 25668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__CLK
timestamp 1667941163
transform 1 0 27140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__CLK
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__CLK
timestamp 1667941163
transform 1 0 25760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__CLK
timestamp 1667941163
transform 1 0 26312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__CLK
timestamp 1667941163
transform -1 0 27416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__CLK
timestamp 1667941163
transform -1 0 37628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__D
timestamp 1667941163
transform -1 0 37260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__CLK
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__CLK
timestamp 1667941163
transform 1 0 35512 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__D
timestamp 1667941163
transform 1 0 22264 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__CLK
timestamp 1667941163
transform 1 0 22816 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__D
timestamp 1667941163
transform 1 0 22816 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__CLK
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__D
timestamp 1667941163
transform 1 0 26496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__CLK
timestamp 1667941163
transform 1 0 28980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__CLK
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__D
timestamp 1667941163
transform 1 0 30728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__CLK
timestamp 1667941163
transform 1 0 36064 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__D
timestamp 1667941163
transform -1 0 36800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__CLK
timestamp 1667941163
transform 1 0 27692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__D
timestamp 1667941163
transform 1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__CLK
timestamp 1667941163
transform 1 0 27140 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__D
timestamp 1667941163
transform 1 0 26404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__CLK
timestamp 1667941163
transform 1 0 23368 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__D
timestamp 1667941163
transform 1 0 29072 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__CLK
timestamp 1667941163
transform 1 0 36340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__D
timestamp 1667941163
transform -1 0 36156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__CLK
timestamp 1667941163
transform 1 0 34868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__CLK
timestamp 1667941163
transform 1 0 36616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__CLK
timestamp 1667941163
transform 1 0 34868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__CLK
timestamp 1667941163
transform 1 0 25852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__CLK
timestamp 1667941163
transform 1 0 35604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__CLK
timestamp 1667941163
transform 1 0 34868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A
timestamp 1667941163
transform -1 0 38272 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 1667941163
transform -1 0 23828 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 1667941163
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A
timestamp 1667941163
transform 1 0 21252 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A
timestamp 1667941163
transform -1 0 20516 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A
timestamp 1667941163
transform 1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1667941163
transform 1 0 23368 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 1667941163
transform -1 0 2852 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A
timestamp 1667941163
transform -1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1667941163
transform -1 0 10028 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A
timestamp 1667941163
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A
timestamp 1667941163
transform 1 0 2392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 1667941163
transform -1 0 29348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A
timestamp 1667941163
transform -1 0 2668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1667941163
transform 1 0 38088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A
timestamp 1667941163
transform 1 0 20608 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A
timestamp 1667941163
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 1667941163
transform -1 0 24840 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A
timestamp 1667941163
transform -1 0 20608 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1667941163
transform -1 0 16836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A
timestamp 1667941163
transform -1 0 24472 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1667941163
transform 1 0 14628 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1667941163
transform -1 0 20884 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A
timestamp 1667941163
transform -1 0 22264 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1667941163
transform 1 0 17940 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1667941163
transform 1 0 25760 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1667941163
transform -1 0 30912 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A
timestamp 1667941163
transform -1 0 8096 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1667941163
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1667941163
transform -1 0 7728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 37720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 1748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 1748 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 37720 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 37628 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 19688 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 1748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 36156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 24748 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 35052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform 1 0 34224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 37628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 11868 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 36708 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 22172 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 2484 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 37812 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 11960 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 37628 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 35972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 1748 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform 1 0 16192 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 9936 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1667941163
transform 1 0 37444 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output42_A
timestamp 1667941163
transform -1 0 8096 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output47_A
timestamp 1667941163
transform -1 0 2484 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1667941163
transform -1 0 2484 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1667941163
transform -1 0 3220 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output59_A
timestamp 1667941163
transform 1 0 2300 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1667941163
transform -1 0 36708 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1667941163
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output67_A
timestamp 1667941163
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1667941163
transform 1 0 7912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1667941163
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1667941163
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1667941163
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76
timestamp 1667941163
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99
timestamp 1667941163
transform 1 0 10212 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1667941163
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_126
timestamp 1667941163
transform 1 0 12696 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1667941163
transform 1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1667941163
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1667941163
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1667941163
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_203
timestamp 1667941163
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 1667941163
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_217
timestamp 1667941163
transform 1 0 21068 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1667941163
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1667941163
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1667941163
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1667941163
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_354
timestamp 1667941163
transform 1 0 33672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1667941163
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_25
timestamp 1667941163
transform 1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1667941163
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_43
timestamp 1667941163
transform 1 0 5060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_175
timestamp 1667941163
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1667941163
transform 1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_185
timestamp 1667941163
transform 1 0 18124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1667941163
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1667941163
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1667941163
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1667941163
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_264
timestamp 1667941163
transform 1 0 25392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_272
timestamp 1667941163
transform 1 0 26128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_285
timestamp 1667941163
transform 1 0 27324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_291
timestamp 1667941163
transform 1 0 27876 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1667941163
transform 1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_323
timestamp 1667941163
transform 1 0 30820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1667941163
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_359
timestamp 1667941163
transform 1 0 34132 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_366
timestamp 1667941163
transform 1 0 34776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_379
timestamp 1667941163
transform 1 0 35972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1667941163
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1667941163
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1667941163
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1667941163
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_229
timestamp 1667941163
transform 1 0 22172 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_276
timestamp 1667941163
transform 1 0 26496 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_300
timestamp 1667941163
transform 1 0 28704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1667941163
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_331
timestamp 1667941163
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_355
timestamp 1667941163
transform 1 0 33764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1667941163
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_370
timestamp 1667941163
transform 1 0 35144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_376
timestamp 1667941163
transform 1 0 35696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_382
timestamp 1667941163
transform 1 0 36248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_388
timestamp 1667941163
transform 1 0 36800 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_394
timestamp 1667941163
transform 1 0 37352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7
timestamp 1667941163
transform 1 0 1748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_19
timestamp 1667941163
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_31
timestamp 1667941163
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_43
timestamp 1667941163
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_211
timestamp 1667941163
transform 1 0 20516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1667941163
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1667941163
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1667941163
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_238
timestamp 1667941163
transform 1 0 23000 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1667941163
transform 1 0 25484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1667941163
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1667941163
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_285
timestamp 1667941163
transform 1 0 27324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_291
timestamp 1667941163
transform 1 0 27876 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_295
timestamp 1667941163
transform 1 0 28244 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_323
timestamp 1667941163
transform 1 0 30820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_327
timestamp 1667941163
transform 1 0 31188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1667941163
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_342
timestamp 1667941163
transform 1 0 32568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_356
timestamp 1667941163
transform 1 0 33856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_363
timestamp 1667941163
transform 1 0 34500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_369
timestamp 1667941163
transform 1 0 35052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_375
timestamp 1667941163
transform 1 0 35604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_381
timestamp 1667941163
transform 1 0 36156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1667941163
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_397
timestamp 1667941163
transform 1 0 37628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_213
timestamp 1667941163
transform 1 0 20700 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_231
timestamp 1667941163
transform 1 0 22356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_235
timestamp 1667941163
transform 1 0 22724 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_238
timestamp 1667941163
transform 1 0 23000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_244
timestamp 1667941163
transform 1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1667941163
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_275
timestamp 1667941163
transform 1 0 26404 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_299
timestamp 1667941163
transform 1 0 28612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1667941163
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1667941163
transform 1 0 31556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1667941163
transform 1 0 31924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_339
timestamp 1667941163
transform 1 0 32292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_346
timestamp 1667941163
transform 1 0 32936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_353
timestamp 1667941163
transform 1 0 33580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1667941163
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_369
timestamp 1667941163
transform 1 0 35052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_375
timestamp 1667941163
transform 1 0 35604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_381
timestamp 1667941163
transform 1 0 36156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_387
timestamp 1667941163
transform 1 0 36708 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_393
timestamp 1667941163
transform 1 0 37260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_402
timestamp 1667941163
transform 1 0 38088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1667941163
transform 1 0 38456 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_201
timestamp 1667941163
transform 1 0 19596 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_212
timestamp 1667941163
transform 1 0 20608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1667941163
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_230
timestamp 1667941163
transform 1 0 22264 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_241
timestamp 1667941163
transform 1 0 23276 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_263
timestamp 1667941163
transform 1 0 25300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_269
timestamp 1667941163
transform 1 0 25852 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_275
timestamp 1667941163
transform 1 0 26404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1667941163
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_285
timestamp 1667941163
transform 1 0 27324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_291
timestamp 1667941163
transform 1 0 27876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_295
timestamp 1667941163
transform 1 0 28244 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_316
timestamp 1667941163
transform 1 0 30176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_327
timestamp 1667941163
transform 1 0 31188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1667941163
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_341
timestamp 1667941163
transform 1 0 32476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_351
timestamp 1667941163
transform 1 0 33396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_368
timestamp 1667941163
transform 1 0 34960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_374
timestamp 1667941163
transform 1 0 35512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_380
timestamp 1667941163
transform 1 0 36064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_386
timestamp 1667941163
transform 1 0 36616 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_397
timestamp 1667941163
transform 1 0 37628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_9
timestamp 1667941163
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1667941163
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_44
timestamp 1667941163
transform 1 0 5152 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_50
timestamp 1667941163
transform 1 0 5704 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_62
timestamp 1667941163
transform 1 0 6808 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_74
timestamp 1667941163
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1667941163
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_226
timestamp 1667941163
transform 1 0 21896 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_232
timestamp 1667941163
transform 1 0 22448 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 1667941163
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_257
timestamp 1667941163
transform 1 0 24748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_261
timestamp 1667941163
transform 1 0 25116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_282
timestamp 1667941163
transform 1 0 27048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1667941163
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_331
timestamp 1667941163
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_338
timestamp 1667941163
transform 1 0 32200 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_344
timestamp 1667941163
transform 1 0 32752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_351
timestamp 1667941163
transform 1 0 33396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_358
timestamp 1667941163
transform 1 0 34040 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_370
timestamp 1667941163
transform 1 0 35144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_376
timestamp 1667941163
transform 1 0 35696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_382
timestamp 1667941163
transform 1 0 36248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_388
timestamp 1667941163
transform 1 0 36800 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_398
timestamp 1667941163
transform 1 0 37720 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_236
timestamp 1667941163
transform 1 0 22816 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_242
timestamp 1667941163
transform 1 0 23368 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_264
timestamp 1667941163
transform 1 0 25392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_270
timestamp 1667941163
transform 1 0 25944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1667941163
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_285
timestamp 1667941163
transform 1 0 27324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_314
timestamp 1667941163
transform 1 0 29992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1667941163
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_327
timestamp 1667941163
transform 1 0 31188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1667941163
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_342
timestamp 1667941163
transform 1 0 32568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_356
timestamp 1667941163
transform 1 0 33856 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_363
timestamp 1667941163
transform 1 0 34500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_369
timestamp 1667941163
transform 1 0 35052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_375
timestamp 1667941163
transform 1 0 35604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_381
timestamp 1667941163
transform 1 0 36156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_389
timestamp 1667941163
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_399
timestamp 1667941163
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_205
timestamp 1667941163
transform 1 0 19964 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_217
timestamp 1667941163
transform 1 0 21068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_229
timestamp 1667941163
transform 1 0 22172 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_276
timestamp 1667941163
transform 1 0 26496 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_332
timestamp 1667941163
transform 1 0 31648 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_339
timestamp 1667941163
transform 1 0 32292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_346
timestamp 1667941163
transform 1 0 32936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_353
timestamp 1667941163
transform 1 0 33580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1667941163
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_369
timestamp 1667941163
transform 1 0 35052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_381
timestamp 1667941163
transform 1 0 36156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_393
timestamp 1667941163
transform 1 0 37260 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_405
timestamp 1667941163
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1667941163
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_144
timestamp 1667941163
transform 1 0 14352 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_150
timestamp 1667941163
transform 1 0 14904 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1667941163
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_234
timestamp 1667941163
transform 1 0 22632 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_263
timestamp 1667941163
transform 1 0 25300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_269
timestamp 1667941163
transform 1 0 25852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1667941163
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_289
timestamp 1667941163
transform 1 0 27692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1667941163
transform 1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_322
timestamp 1667941163
transform 1 0 30728 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_330
timestamp 1667941163
transform 1 0 31464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1667941163
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_342
timestamp 1667941163
transform 1 0 32568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_355
timestamp 1667941163
transform 1 0 33764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_367
timestamp 1667941163
transform 1 0 34868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_379
timestamp 1667941163
transform 1 0 35972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_401
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_9
timestamp 1667941163
transform 1 0 1932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1667941163
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_226
timestamp 1667941163
transform 1 0 21896 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1667941163
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_285
timestamp 1667941163
transform 1 0 27324 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_291
timestamp 1667941163
transform 1 0 27876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_297
timestamp 1667941163
transform 1 0 28428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_300
timestamp 1667941163
transform 1 0 28704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1667941163
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_331
timestamp 1667941163
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_338
timestamp 1667941163
transform 1 0 32200 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1667941163
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_232
timestamp 1667941163
transform 1 0 22448 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_238
timestamp 1667941163
transform 1 0 23000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_259
timestamp 1667941163
transform 1 0 24932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_266
timestamp 1667941163
transform 1 0 25576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_285
timestamp 1667941163
transform 1 0 27324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_307
timestamp 1667941163
transform 1 0 29348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_331
timestamp 1667941163
transform 1 0 31556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1667941163
transform 1 0 20700 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_217
timestamp 1667941163
transform 1 0 21068 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_230
timestamp 1667941163
transform 1 0 22264 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_262
timestamp 1667941163
transform 1 0 25208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_269
timestamp 1667941163
transform 1 0 25852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_276
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_286
timestamp 1667941163
transform 1 0 27416 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_298
timestamp 1667941163
transform 1 0 28520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1667941163
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_313
timestamp 1667941163
transform 1 0 29900 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_324
timestamp 1667941163
transform 1 0 30912 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_336
timestamp 1667941163
transform 1 0 32016 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_348
timestamp 1667941163
transform 1 0 33120 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1667941163
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_397
timestamp 1667941163
transform 1 0 37628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_7
timestamp 1667941163
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_19
timestamp 1667941163
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1667941163
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_43
timestamp 1667941163
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_232
timestamp 1667941163
transform 1 0 22448 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_244
timestamp 1667941163
transform 1 0 23552 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_259
timestamp 1667941163
transform 1 0 24932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1667941163
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_146
timestamp 1667941163
transform 1 0 14536 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_158
timestamp 1667941163
transform 1 0 15640 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_170
timestamp 1667941163
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_183
timestamp 1667941163
transform 1 0 17940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_238
timestamp 1667941163
transform 1 0 23000 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_244
timestamp 1667941163
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_279
timestamp 1667941163
transform 1 0 26772 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_286
timestamp 1667941163
transform 1 0 27416 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_298
timestamp 1667941163
transform 1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1667941163
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_351
timestamp 1667941163
transform 1 0 33396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_355
timestamp 1667941163
transform 1 0 33764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1667941163
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1667941163
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1667941163
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1667941163
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_236
timestamp 1667941163
transform 1 0 22816 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_243
timestamp 1667941163
transform 1 0 23460 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_253
timestamp 1667941163
transform 1 0 24380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1667941163
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_301
timestamp 1667941163
transform 1 0 28796 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_307
timestamp 1667941163
transform 1 0 29348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_319
timestamp 1667941163
transform 1 0 30452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 1667941163
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_379
timestamp 1667941163
transform 1 0 35972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_384
timestamp 1667941163
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_401
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_9
timestamp 1667941163
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1667941163
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_162
timestamp 1667941163
transform 1 0 16008 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_168
timestamp 1667941163
transform 1 0 16560 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_180
timestamp 1667941163
transform 1 0 17664 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1667941163
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_215
timestamp 1667941163
transform 1 0 20884 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1667941163
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_226
timestamp 1667941163
transform 1 0 21896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_240
timestamp 1667941163
transform 1 0 23184 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1667941163
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_268
timestamp 1667941163
transform 1 0 25760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_281
timestamp 1667941163
transform 1 0 26956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_287
timestamp 1667941163
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_293
timestamp 1667941163
transform 1 0 28060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1667941163
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_215
timestamp 1667941163
transform 1 0 20884 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_244
timestamp 1667941163
transform 1 0 23552 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_252
timestamp 1667941163
transform 1 0 24288 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_266
timestamp 1667941163
transform 1 0 25576 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1667941163
transform 1 0 27416 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_33
timestamp 1667941163
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_37
timestamp 1667941163
transform 1 0 4508 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_43
timestamp 1667941163
transform 1 0 5060 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_55
timestamp 1667941163
transform 1 0 6164 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_67
timestamp 1667941163
transform 1 0 7268 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp 1667941163
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_183
timestamp 1667941163
transform 1 0 17940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_205
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1667941163
transform 1 0 20240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1667941163
transform 1 0 20884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_222
timestamp 1667941163
transform 1 0 21528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_235
timestamp 1667941163
transform 1 0 22724 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1667941163
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_272
timestamp 1667941163
transform 1 0 26128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_285
timestamp 1667941163
transform 1 0 27324 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_292
timestamp 1667941163
transform 1 0 27968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_299
timestamp 1667941163
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1667941163
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1667941163
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1667941163
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_231
timestamp 1667941163
transform 1 0 22356 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_236
timestamp 1667941163
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_262
timestamp 1667941163
transform 1 0 25208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_269
timestamp 1667941163
transform 1 0 25852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1667941163
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1667941163
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_300
timestamp 1667941163
transform 1 0 28704 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_306
timestamp 1667941163
transform 1 0 29256 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_318
timestamp 1667941163
transform 1 0 30360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_330
timestamp 1667941163
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_9
timestamp 1667941163
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1667941163
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_101
timestamp 1667941163
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_105
timestamp 1667941163
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_111
timestamp 1667941163
transform 1 0 11316 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_123
timestamp 1667941163
transform 1 0 12420 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1667941163
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1667941163
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_226
timestamp 1667941163
transform 1 0 21896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_239
timestamp 1667941163
transform 1 0 23092 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1667941163
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_264
timestamp 1667941163
transform 1 0 25392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp 1667941163
transform 1 0 26496 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_283
timestamp 1667941163
transform 1 0 27140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_295
timestamp 1667941163
transform 1 0 28244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_199
timestamp 1667941163
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_231
timestamp 1667941163
transform 1 0 22356 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_239
timestamp 1667941163
transform 1 0 23092 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_243
timestamp 1667941163
transform 1 0 23460 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_250
timestamp 1667941163
transform 1 0 24104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_263
timestamp 1667941163
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_267
timestamp 1667941163
transform 1 0 25668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1667941163
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_286
timestamp 1667941163
transform 1 0 27416 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_298
timestamp 1667941163
transform 1 0 28520 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_310
timestamp 1667941163
transform 1 0 29624 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_322
timestamp 1667941163
transform 1 0 30728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1667941163
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_402
timestamp 1667941163
transform 1 0 38088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_406
timestamp 1667941163
transform 1 0 38456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1667941163
transform 1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_17
timestamp 1667941163
transform 1 0 2668 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1667941163
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_117
timestamp 1667941163
transform 1 0 11868 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_122
timestamp 1667941163
transform 1 0 12328 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_128
timestamp 1667941163
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_236
timestamp 1667941163
transform 1 0 22816 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1667941163
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_271
timestamp 1667941163
transform 1 0 26036 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1667941163
transform 1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_294
timestamp 1667941163
transform 1 0 28152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1667941163
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_373
timestamp 1667941163
transform 1 0 35420 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_404
timestamp 1667941163
transform 1 0 38272 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1667941163
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1667941163
transform 1 0 12420 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_129
timestamp 1667941163
transform 1 0 12972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_141
timestamp 1667941163
transform 1 0 14076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_153
timestamp 1667941163
transform 1 0 15180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1667941163
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_250
timestamp 1667941163
transform 1 0 24104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_263
timestamp 1667941163
transform 1 0 25300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_270
timestamp 1667941163
transform 1 0 25944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1667941163
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_291
timestamp 1667941163
transform 1 0 27876 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_298
timestamp 1667941163
transform 1 0 28520 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_310
timestamp 1667941163
transform 1 0 29624 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_322
timestamp 1667941163
transform 1 0 30728 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1667941163
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_9
timestamp 1667941163
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1667941163
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_61
timestamp 1667941163
transform 1 0 6716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_66
timestamp 1667941163
transform 1 0 7176 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_72
timestamp 1667941163
transform 1 0 7728 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_223
timestamp 1667941163
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_231
timestamp 1667941163
transform 1 0 22356 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_244
timestamp 1667941163
transform 1 0 23552 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_263
timestamp 1667941163
transform 1 0 25300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_275
timestamp 1667941163
transform 1 0 26404 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_282
timestamp 1667941163
transform 1 0 27048 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_296
timestamp 1667941163
transform 1 0 28336 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1667941163
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_205
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_209
timestamp 1667941163
transform 1 0 20332 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_212
timestamp 1667941163
transform 1 0 20608 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_218
timestamp 1667941163
transform 1 0 21160 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_229
timestamp 1667941163
transform 1 0 22172 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_238
timestamp 1667941163
transform 1 0 23000 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1667941163
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_263
timestamp 1667941163
transform 1 0 25300 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1667941163
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_286
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_292
timestamp 1667941163
transform 1 0 27968 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_304
timestamp 1667941163
transform 1 0 29072 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_316
timestamp 1667941163
transform 1 0 30176 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_328
timestamp 1667941163
transform 1 0 31280 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_10
timestamp 1667941163
transform 1 0 2024 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_16
timestamp 1667941163
transform 1 0 2576 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1667941163
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_107
timestamp 1667941163
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_119
timestamp 1667941163
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_131
timestamp 1667941163
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 1667941163
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_210
timestamp 1667941163
transform 1 0 20424 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_228
timestamp 1667941163
transform 1 0 22080 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1667941163
transform 1 0 23276 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1667941163
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_258
timestamp 1667941163
transform 1 0 24840 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_275
timestamp 1667941163
transform 1 0 26404 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_282
timestamp 1667941163
transform 1 0 27048 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_295
timestamp 1667941163
transform 1 0 28244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1667941163
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1667941163
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1667941163
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1667941163
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1667941163
transform 1 0 20700 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_216
timestamp 1667941163
transform 1 0 20976 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_234
timestamp 1667941163
transform 1 0 22632 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_247
timestamp 1667941163
transform 1 0 23828 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_254
timestamp 1667941163
transform 1 0 24472 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_260
timestamp 1667941163
transform 1 0 25024 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1667941163
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_299
timestamp 1667941163
transform 1 0 28612 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_311
timestamp 1667941163
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_323
timestamp 1667941163
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_398
timestamp 1667941163
transform 1 0 37720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_213
timestamp 1667941163
transform 1 0 20700 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1667941163
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_226
timestamp 1667941163
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1667941163
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_263
timestamp 1667941163
transform 1 0 25300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_275
timestamp 1667941163
transform 1 0 26404 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_282
timestamp 1667941163
transform 1 0 27048 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_295
timestamp 1667941163
transform 1 0 28244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_314
timestamp 1667941163
transform 1 0 29992 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_326
timestamp 1667941163
transform 1 0 31096 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_338
timestamp 1667941163
transform 1 0 32200 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_350
timestamp 1667941163
transform 1 0 33304 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1667941163
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1667941163
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1667941163
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_229
timestamp 1667941163
transform 1 0 22172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_242
timestamp 1667941163
transform 1 0 23368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_254
timestamp 1667941163
transform 1 0 24472 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_262
timestamp 1667941163
transform 1 0 25208 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1667941163
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_285
timestamp 1667941163
transform 1 0 27324 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_297
timestamp 1667941163
transform 1 0 28428 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_309
timestamp 1667941163
transform 1 0 29532 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_321
timestamp 1667941163
transform 1 0 30636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1667941163
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_401
timestamp 1667941163
transform 1 0 37996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_404
timestamp 1667941163
transform 1 0 38272 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_7
timestamp 1667941163
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_19
timestamp 1667941163
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_102
timestamp 1667941163
transform 1 0 10488 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_108
timestamp 1667941163
transform 1 0 11040 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_120
timestamp 1667941163
transform 1 0 12144 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1667941163
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1667941163
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_231
timestamp 1667941163
transform 1 0 22356 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_237
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1667941163
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1667941163
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_272
timestamp 1667941163
transform 1 0 26128 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_278
timestamp 1667941163
transform 1 0 26680 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1667941163
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_290
timestamp 1667941163
transform 1 0 27784 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1667941163
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_397
timestamp 1667941163
transform 1 0 37628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_402
timestamp 1667941163
transform 1 0 38088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1667941163
transform 1 0 38456 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1667941163
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_243
timestamp 1667941163
transform 1 0 23460 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_264
timestamp 1667941163
transform 1 0 25392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1667941163
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_91
timestamp 1667941163
transform 1 0 9476 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_171
timestamp 1667941163
transform 1 0 16836 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_225
timestamp 1667941163
transform 1 0 21804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1667941163
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_240
timestamp 1667941163
transform 1 0 23184 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_260
timestamp 1667941163
transform 1 0 25024 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_266
timestamp 1667941163
transform 1 0 25576 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_272
timestamp 1667941163
transform 1 0 26128 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_284
timestamp 1667941163
transform 1 0 27232 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_296
timestamp 1667941163
transform 1 0 28336 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_399
timestamp 1667941163
transform 1 0 37812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_7
timestamp 1667941163
transform 1 0 1748 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_19
timestamp 1667941163
transform 1 0 2852 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_31
timestamp 1667941163
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_43
timestamp 1667941163
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_250
timestamp 1667941163
transform 1 0 24104 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_256
timestamp 1667941163
transform 1 0 24656 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_266
timestamp 1667941163
transform 1 0 25576 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_286
timestamp 1667941163
transform 1 0 27416 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_292
timestamp 1667941163
transform 1 0 27968 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_304
timestamp 1667941163
transform 1 0 29072 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_316
timestamp 1667941163
transform 1 0 30176 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_328
timestamp 1667941163
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_402
timestamp 1667941163
transform 1 0 38088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_406
timestamp 1667941163
transform 1 0 38456 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_9
timestamp 1667941163
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1667941163
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_205
timestamp 1667941163
transform 1 0 19964 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_211
timestamp 1667941163
transform 1 0 20516 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_223
timestamp 1667941163
transform 1 0 21620 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_231
timestamp 1667941163
transform 1 0 22356 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_236
timestamp 1667941163
transform 1 0 22816 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_240
timestamp 1667941163
transform 1 0 23184 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_244
timestamp 1667941163
transform 1 0 23552 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1667941163
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_257
timestamp 1667941163
transform 1 0 24748 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_269
timestamp 1667941163
transform 1 0 25852 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_281
timestamp 1667941163
transform 1 0 26956 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_293
timestamp 1667941163
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1667941163
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_318
timestamp 1667941163
transform 1 0 30360 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_324
timestamp 1667941163
transform 1 0 30912 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_336
timestamp 1667941163
transform 1 0 32016 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_348
timestamp 1667941163
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1667941163
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_234
timestamp 1667941163
transform 1 0 22632 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_241
timestamp 1667941163
transform 1 0 23276 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1667941163
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_259
timestamp 1667941163
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_271
timestamp 1667941163
transform 1 0 26036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1667941163
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1667941163
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_19
timestamp 1667941163
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_226
timestamp 1667941163
transform 1 0 21896 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_262
timestamp 1667941163
transform 1 0 25208 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_268
timestamp 1667941163
transform 1 0 25760 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_280
timestamp 1667941163
transform 1 0 26864 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_292
timestamp 1667941163
transform 1 0 27968 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1667941163
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_9
timestamp 1667941163
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_21
timestamp 1667941163
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1667941163
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1667941163
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1667941163
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_241
timestamp 1667941163
transform 1 0 23276 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_253
timestamp 1667941163
transform 1 0 24380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_257
timestamp 1667941163
transform 1 0 24748 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_267
timestamp 1667941163
transform 1 0 25668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_7
timestamp 1667941163
transform 1 0 1748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_19
timestamp 1667941163
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_70
timestamp 1667941163
transform 1 0 7544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1667941163
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_242
timestamp 1667941163
transform 1 0 23368 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_261
timestamp 1667941163
transform 1 0 25116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_266
timestamp 1667941163
transform 1 0 25576 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_272
timestamp 1667941163
transform 1 0 26128 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_284
timestamp 1667941163
transform 1 0 27232 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_296
timestamp 1667941163
transform 1 0 28336 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_239
timestamp 1667941163
transform 1 0 23092 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_260
timestamp 1667941163
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_268
timestamp 1667941163
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_285
timestamp 1667941163
transform 1 0 27324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_297
timestamp 1667941163
transform 1 0 28428 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_301
timestamp 1667941163
transform 1 0 28796 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_307
timestamp 1667941163
transform 1 0 29348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_319
timestamp 1667941163
transform 1 0 30452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1667941163
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_270
timestamp 1667941163
transform 1 0 25944 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_282
timestamp 1667941163
transform 1 0 27048 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_294
timestamp 1667941163
transform 1 0 28152 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1667941163
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_21
timestamp 1667941163
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_33
timestamp 1667941163
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1667941163
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_397
timestamp 1667941163
transform 1 0 37628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1667941163
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_7
timestamp 1667941163
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1667941163
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_161
timestamp 1667941163
transform 1 0 15916 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_171
timestamp 1667941163
transform 1 0 16836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_183
timestamp 1667941163
transform 1 0 17940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_229
timestamp 1667941163
transform 1 0 22172 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_235
timestamp 1667941163
transform 1 0 22724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_241
timestamp 1667941163
transform 1 0 23276 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1667941163
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_234
timestamp 1667941163
transform 1 0 22632 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_240
timestamp 1667941163
transform 1 0 23184 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_252
timestamp 1667941163
transform 1 0 24288 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_264
timestamp 1667941163
transform 1 0 25392 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_268
timestamp 1667941163
transform 1 0 25760 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1667941163
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_237
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_241
timestamp 1667941163
transform 1 0 23276 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_247
timestamp 1667941163
transform 1 0 23828 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_9
timestamp 1667941163
transform 1 0 1932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_21
timestamp 1667941163
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_33
timestamp 1667941163
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1667941163
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_143
timestamp 1667941163
transform 1 0 14260 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_233
timestamp 1667941163
transform 1 0 22540 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_238
timestamp 1667941163
transform 1 0 23000 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_244
timestamp 1667941163
transform 1 0 23552 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_256
timestamp 1667941163
transform 1 0 24656 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_268
timestamp 1667941163
transform 1 0 25760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_189
timestamp 1667941163
transform 1 0 18492 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_195
timestamp 1667941163
transform 1 0 19044 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_207
timestamp 1667941163
transform 1 0 20148 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_219
timestamp 1667941163
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_105
timestamp 1667941163
transform 1 0 10764 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_113
timestamp 1667941163
transform 1 0 11500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_125
timestamp 1667941163
transform 1 0 12604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 1667941163
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_240
timestamp 1667941163
transform 1 0 23184 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_248
timestamp 1667941163
transform 1 0 23920 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_254
timestamp 1667941163
transform 1 0 24472 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_262
timestamp 1667941163
transform 1 0 25208 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_266
timestamp 1667941163
transform 1 0 25576 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1667941163
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_7
timestamp 1667941163
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1667941163
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_267
timestamp 1667941163
transform 1 0 25668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_397
timestamp 1667941163
transform 1 0 37628 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_7
timestamp 1667941163
transform 1 0 1748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_11
timestamp 1667941163
transform 1 0 2116 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_17
timestamp 1667941163
transform 1 0 2668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_29
timestamp 1667941163
transform 1 0 3772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_41
timestamp 1667941163
transform 1 0 4876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1667941163
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_23
timestamp 1667941163
transform 1 0 3220 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_28
timestamp 1667941163
transform 1 0 3680 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_34
timestamp 1667941163
transform 1 0 4232 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_46
timestamp 1667941163
transform 1 0 5336 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_117
timestamp 1667941163
transform 1 0 11868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_129
timestamp 1667941163
transform 1 0 12972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_141
timestamp 1667941163
transform 1 0 14076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_153
timestamp 1667941163
transform 1 0 15180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_165
timestamp 1667941163
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_177
timestamp 1667941163
transform 1 0 17388 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_183
timestamp 1667941163
transform 1 0 17940 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_195
timestamp 1667941163
transform 1 0 19044 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_207
timestamp 1667941163
transform 1 0 20148 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_211
timestamp 1667941163
transform 1 0 20516 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_214
timestamp 1667941163
transform 1 0 20792 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 1667941163
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_252
timestamp 1667941163
transform 1 0 24288 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_258
timestamp 1667941163
transform 1 0 24840 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_266
timestamp 1667941163
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_298
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_310
timestamp 1667941163
transform 1 0 29624 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_323
timestamp 1667941163
transform 1 0 30820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_387
timestamp 1667941163
transform 1 0 36708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_17
timestamp 1667941163
transform 1 0 2668 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_43
timestamp 1667941163
transform 1 0 5060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_49
timestamp 1667941163
transform 1 0 5612 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1667941163
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_65
timestamp 1667941163
transform 1 0 7084 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_70
timestamp 1667941163
transform 1 0 7544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1667941163
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_96
timestamp 1667941163
transform 1 0 9936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_118
timestamp 1667941163
transform 1 0 11960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1667941163
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1667941163
transform 1 0 15732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_163
timestamp 1667941163
transform 1 0 16100 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_202
timestamp 1667941163
transform 1 0 19688 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_216
timestamp 1667941163
transform 1 0 20976 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_239
timestamp 1667941163
transform 1 0 23092 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1667941163
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_257
timestamp 1667941163
transform 1 0 24748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_261
timestamp 1667941163
transform 1 0 25116 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_274
timestamp 1667941163
transform 1 0 26312 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_323
timestamp 1667941163
transform 1 0 30820 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1667941163
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_355
timestamp 1667941163
transform 1 0 33764 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_359
timestamp 1667941163
transform 1 0 34132 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _115_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 25576 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1667941163
transform -1 0 27140 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1667941163
transform 1 0 27784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1667941163
transform -1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1667941163
transform -1 0 27416 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 1667941163
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1667941163
transform -1 0 27416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1667941163
transform -1 0 24104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1667941163
transform -1 0 24104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1667941163
transform -1 0 27048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1667941163
transform -1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _126_
timestamp 1667941163
transform 1 0 24932 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1667941163
transform 1 0 24748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _128_
timestamp 1667941163
transform -1 0 26404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1667941163
transform 1 0 22356 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _130_
timestamp 1667941163
transform -1 0 23276 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 1667941163
transform 1 0 22264 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _132_
timestamp 1667941163
transform -1 0 21528 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _133_
timestamp 1667941163
transform -1 0 23460 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _134_
timestamp 1667941163
transform 1 0 24196 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1667941163
transform -1 0 25484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1667941163
transform -1 0 28520 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1667941163
transform 1 0 22632 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1667941163
transform 1 0 22356 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 1667941163
transform -1 0 22356 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1667941163
transform -1 0 27692 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1667941163
transform -1 0 24840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1667941163
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1667941163
transform 1 0 21160 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1667941163
transform -1 0 27692 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1667941163
transform 1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp 1667941163
transform -1 0 22540 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1667941163
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1667941163
transform -1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _150_
timestamp 1667941163
transform -1 0 23460 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1667941163
transform 1 0 24104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152_
timestamp 1667941163
transform -1 0 21528 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _153_
timestamp 1667941163
transform -1 0 21160 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1667941163
transform -1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1667941163
transform -1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1667941163
transform -1 0 21528 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 1667941163
transform -1 0 23184 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1667941163
transform -1 0 22448 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1667941163
transform -1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1667941163
transform -1 0 28060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1667941163
transform -1 0 23460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1667941163
transform 1 0 26772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1667941163
transform -1 0 28612 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1667941163
transform 1 0 25576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1667941163
transform -1 0 27692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1667941163
transform -1 0 27416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1667941163
transform -1 0 27048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1667941163
transform -1 0 25944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1667941163
transform 1 0 27784 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1667941163
transform -1 0 23644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1667941163
transform 1 0 21620 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1667941163
transform -1 0 26220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1667941163
transform -1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1667941163
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1667941163
transform 1 0 20608 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1667941163
transform -1 0 27968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1667941163
transform -1 0 22540 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1667941163
transform 1 0 29072 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1667941163
transform -1 0 21528 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1667941163
transform -1 0 26496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1667941163
transform 1 0 22172 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _184_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21528 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1667941163
transform 1 0 17112 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1667941163
transform -1 0 2116 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1667941163
transform -1 0 28704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1667941163
transform 1 0 19136 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1667941163
transform -1 0 25576 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1667941163
transform 1 0 20792 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1667941163
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1667941163
transform -1 0 33764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1667941163
transform 1 0 24104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1667941163
transform 1 0 25484 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _196_
timestamp 1667941163
transform -1 0 24012 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1667941163
transform 1 0 22724 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1667941163
transform -1 0 28336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1667941163
transform -1 0 26220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1667941163
transform -1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1667941163
transform -1 0 21528 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1667941163
transform -1 0 22264 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _203_
timestamp 1667941163
transform 1 0 22448 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1667941163
transform 1 0 10488 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1667941163
transform 1 0 12052 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1667941163
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1667941163
transform 1 0 29992 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1667941163
transform 1 0 22908 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1667941163
transform 1 0 18768 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1667941163
transform 1 0 16560 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1667941163
transform -1 0 27416 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1667941163
transform -1 0 23552 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _213_
timestamp 1667941163
transform 1 0 21988 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _214_
timestamp 1667941163
transform -1 0 3680 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1667941163
transform -1 0 22632 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1667941163
transform 1 0 10212 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform -1 0 25576 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform 1 0 22448 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform -1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform 1 0 22632 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform -1 0 27416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform -1 0 25208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform 1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _224_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _225_
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform -1 0 32936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform -1 0 32292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform -1 0 31832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform -1 0 33580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform -1 0 32568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform -1 0 32568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1667941163
transform -1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1667941163
transform 1 0 33580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform -1 0 32200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform -1 0 31832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _236_
timestamp 1667941163
transform 1 0 32844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform -1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform -1 0 34500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform -1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform -1 0 32200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform -1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform -1 0 31832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform -1 0 34040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform -1 0 33212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform -1 0 34960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform 1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _247_
timestamp 1667941163
transform -1 0 34316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform -1 0 34408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform -1 0 33856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform -1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform -1 0 33672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform -1 0 34224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform -1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform -1 0 34776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform 1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform -1 0 34500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform -1 0 31188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform -1 0 32936 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform 1 0 32292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform -1 0 31188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform -1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform -1 0 33580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 31832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _264_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 31556 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _265_
timestamp 1667941163
transform 1 0 29716 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _266_
timestamp 1667941163
transform 1 0 23092 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _267_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 27324 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _268_
timestamp 1667941163
transform 1 0 29716 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _269_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 29992 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _270_
timestamp 1667941163
transform 1 0 28336 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _271_
timestamp 1667941163
transform 1 0 29716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _272_
timestamp 1667941163
transform 1 0 27416 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _273_
timestamp 1667941163
transform 1 0 24564 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _274_
timestamp 1667941163
transform 1 0 23368 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _275_
timestamp 1667941163
transform -1 0 28796 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _276_
timestamp 1667941163
transform 1 0 22264 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _277_
timestamp 1667941163
transform 1 0 25208 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _278_
timestamp 1667941163
transform 1 0 22264 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _279_
timestamp 1667941163
transform -1 0 25300 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _280_
timestamp 1667941163
transform -1 0 25392 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _281_
timestamp 1667941163
transform -1 0 29348 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _282_
timestamp 1667941163
transform 1 0 31924 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _283_
timestamp 1667941163
transform 1 0 29716 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _284_
timestamp 1667941163
transform 1 0 26864 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _285_
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _286_
timestamp 1667941163
transform 1 0 22172 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _287_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _288_
timestamp 1667941163
transform 1 0 28612 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _289_
timestamp 1667941163
transform -1 0 31556 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _290_
timestamp 1667941163
transform 1 0 24564 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _291_
timestamp 1667941163
transform 1 0 23368 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _292_
timestamp 1667941163
transform 1 0 23276 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _293_
timestamp 1667941163
transform -1 0 30820 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _294_
timestamp 1667941163
transform -1 0 31556 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _295_
timestamp 1667941163
transform -1 0 34132 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _296_
timestamp 1667941163
transform 1 0 26772 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _297_
timestamp 1667941163
transform 1 0 22264 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _298_
timestamp 1667941163
transform -1 0 29072 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _299_
timestamp 1667941163
transform -1 0 30268 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _306_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1667941163
transform -1 0 23276 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1667941163
transform 1 0 12144 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1667941163
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _310_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19964 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1667941163
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1667941163
transform -1 0 23552 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1667941163
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1667941163
transform -1 0 17940 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1667941163
transform -1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _316_
timestamp 1667941163
transform -1 0 9476 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1667941163
transform -1 0 26220 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _318_
timestamp 1667941163
transform 1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1667941163
transform 1 0 1748 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1667941163
transform -1 0 28796 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _321_
timestamp 1667941163
transform 1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1667941163
transform -1 0 38088 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1667941163
transform -1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _324_
timestamp 1667941163
transform -1 0 25668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp 1667941163
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1667941163
transform -1 0 24288 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1667941163
transform -1 0 27416 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1667941163
transform 1 0 20608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _329_
timestamp 1667941163
transform -1 0 20424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1667941163
transform 1 0 16008 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _331_
timestamp 1667941163
transform 1 0 36064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1667941163
transform -1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1667941163
transform -1 0 14260 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1667941163
transform 1 0 21252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1667941163
transform -1 0 35788 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1667941163
transform 1 0 21804 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1667941163
transform 1 0 17296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _338_
timestamp 1667941163
transform -1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1667941163
transform -1 0 30360 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1667941163
transform 1 0 7268 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1667941163
transform -1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1667941163
transform -1 0 38088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1667941163
transform 1 0 6900 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _344_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22172 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _345_
timestamp 1667941163
transform -1 0 25300 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _346_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _347_
timestamp 1667941163
transform -1 0 31464 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _348__86 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 21528 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _348_
timestamp 1667941163
transform 1 0 21896 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _349_
timestamp 1667941163
transform -1 0 27324 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _350_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26128 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _351_
timestamp 1667941163
transform -1 0 26772 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _352_
timestamp 1667941163
transform 1 0 22264 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _353_
timestamp 1667941163
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _354_
timestamp 1667941163
transform 1 0 20608 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _355_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _356_
timestamp 1667941163
transform 1 0 25852 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _357__87
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _357_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26404 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _358_
timestamp 1667941163
transform 1 0 25760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _359_
timestamp 1667941163
transform 1 0 25760 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _360_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _361_
timestamp 1667941163
transform -1 0 25484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _362_
timestamp 1667941163
transform 1 0 25668 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _363_
timestamp 1667941163
transform -1 0 23000 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _364_
timestamp 1667941163
transform -1 0 28152 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _365_
timestamp 1667941163
transform 1 0 24564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _366_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _367_
timestamp 1667941163
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _368_
timestamp 1667941163
transform -1 0 21896 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _369_
timestamp 1667941163
transform -1 0 21068 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _370_
timestamp 1667941163
transform -1 0 20608 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _371__88
timestamp 1667941163
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _371_
timestamp 1667941163
transform -1 0 22356 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _372_
timestamp 1667941163
transform -1 0 24012 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _373_
timestamp 1667941163
transform 1 0 21988 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _374_
timestamp 1667941163
transform -1 0 25392 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _375_
timestamp 1667941163
transform 1 0 23092 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _376_
timestamp 1667941163
transform -1 0 22264 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _377_
timestamp 1667941163
transform -1 0 20884 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _378_
timestamp 1667941163
transform 1 0 22080 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _379_
timestamp 1667941163
transform -1 0 24932 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _380_
timestamp 1667941163
transform 1 0 25300 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _381_
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _382_
timestamp 1667941163
transform 1 0 22448 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _383__89
timestamp 1667941163
transform -1 0 21160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _383_
timestamp 1667941163
transform 1 0 22540 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _384_
timestamp 1667941163
transform 1 0 21528 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _385_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _386_
timestamp 1667941163
transform 1 0 21988 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _387_
timestamp 1667941163
transform 1 0 23000 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _388_
timestamp 1667941163
transform 1 0 25208 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _389_
timestamp 1667941163
transform 1 0 23000 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _390_
timestamp 1667941163
transform -1 0 26588 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _391_
timestamp 1667941163
transform 1 0 22724 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _392_
timestamp 1667941163
transform 1 0 22908 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _393_
timestamp 1667941163
transform -1 0 25024 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _394_
timestamp 1667941163
transform 1 0 22632 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _395__90
timestamp 1667941163
transform 1 0 23000 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _395_
timestamp 1667941163
transform 1 0 22908 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _396_
timestamp 1667941163
transform 1 0 23736 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _397_
timestamp 1667941163
transform 1 0 24564 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _398_
timestamp 1667941163
transform -1 0 25576 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _399_
timestamp 1667941163
transform -1 0 25668 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _400_
timestamp 1667941163
transform -1 0 25392 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _401_
timestamp 1667941163
transform 1 0 22356 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _402_
timestamp 1667941163
transform 1 0 22448 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _403_
timestamp 1667941163
transform 1 0 23276 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _404_
timestamp 1667941163
transform 1 0 24380 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _405_
timestamp 1667941163
transform -1 0 26496 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _405__91
timestamp 1667941163
transform -1 0 26496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _406_
timestamp 1667941163
transform 1 0 23368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _407_
timestamp 1667941163
transform 1 0 23276 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _408_
timestamp 1667941163
transform 1 0 24472 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _409_
timestamp 1667941163
transform -1 0 26956 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _410_
timestamp 1667941163
transform 1 0 25208 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _411_
timestamp 1667941163
transform -1 0 25208 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _412_
timestamp 1667941163
transform -1 0 26956 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 38088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 38088 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform -1 0 38364 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38364 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1667941163
transform -1 0 38364 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1667941163
transform -1 0 38364 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1667941163
transform -1 0 24104 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1667941163
transform -1 0 38364 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform -1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform -1 0 35236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform -1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform -1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1667941163
transform -1 0 38364 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1667941163
transform -1 0 11224 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1667941163
transform -1 0 11224 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform -1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1667941163
transform -1 0 38364 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1667941163
transform -1 0 38364 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1667941163
transform -1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform -1 0 38364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform -1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1667941163
transform 1 0 1564 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1667941163
transform 1 0 18032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform -1 0 9384 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform -1 0 7544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform -1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform -1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform -1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform -1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 2300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform -1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform -1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform -1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform -1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 25208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform -1 0 36524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform -1 0 1932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform -1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform -1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 30452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform -1 0 5612 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform -1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform -1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform -1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 21160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform -1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform -1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform -1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 406 592
<< labels >>
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal2 s 14186 200 14242 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_bottom_in[10]
port 3 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chany_bottom_in[11]
port 4 nsew signal input
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chany_bottom_in[12]
port 5 nsew signal input
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 6 nsew signal input
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 chany_bottom_in[14]
port 7 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 8 nsew signal input
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 9 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_bottom_in[17]
port 10 nsew signal input
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chany_bottom_in[18]
port 11 nsew signal input
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 12 nsew signal input
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 13 nsew signal input
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 14 nsew signal input
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 15 nsew signal input
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 16 nsew signal input
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 17 nsew signal input
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 18 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 19 nsew signal input
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 20 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 21 nsew signal tristate
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 22 nsew signal tristate
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 23 nsew signal tristate
flabel metal3 s 39200 12928 39800 13048 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 24 nsew signal tristate
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 chany_bottom_out[13]
port 25 nsew signal tristate
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 26 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_bottom_out[15]
port 27 nsew signal tristate
flabel metal3 s 200 14968 800 15088 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 28 nsew signal tristate
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chany_bottom_out[17]
port 29 nsew signal tristate
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chany_bottom_out[18]
port 30 nsew signal tristate
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 31 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 32 nsew signal tristate
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 33 nsew signal tristate
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 34 nsew signal tristate
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 35 nsew signal tristate
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 36 nsew signal tristate
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 37 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 38 nsew signal tristate
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 39 nsew signal tristate
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal2 s 14186 39200 14242 39800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal2 s 12254 200 12310 800 0 FreeSans 224 90 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 78 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 79 nsew signal tristate
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 80 nsew signal tristate
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 pReset
port 81 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 prog_clk
port 82 nsew signal input
flabel metal3 s 200 12928 800 13048 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
port 83 nsew signal tristate
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 84 nsew signal tristate
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 85 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 86 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 86 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 87 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal2 30130 7650 30130 7650 0 _000_
rlabel metal1 32108 6766 32108 6766 0 _001_
rlabel metal2 27462 7888 27462 7888 0 _002_
rlabel metal1 32062 6664 32062 6664 0 _003_
rlabel metal1 32200 6426 32200 6426 0 _004_
rlabel metal1 29447 6358 29447 6358 0 _005_
rlabel metal2 31050 5678 31050 5678 0 _006_
rlabel metal2 32062 5304 32062 5304 0 _007_
rlabel metal1 28842 5719 28842 5719 0 _008_
rlabel metal1 29440 6426 29440 6426 0 _009_
rlabel metal2 30774 6358 30774 6358 0 _010_
rlabel metal1 28205 6698 28205 6698 0 _011_
rlabel metal2 32154 6528 32154 6528 0 _012_
rlabel metal1 27055 5610 27055 5610 0 _013_
rlabel metal1 23690 6807 23690 6807 0 _014_
rlabel metal1 30360 4998 30360 4998 0 _015_
rlabel metal2 24610 6120 24610 6120 0 _016_
rlabel metal2 30498 7616 30498 7616 0 _017_
rlabel metal1 33350 3543 33350 3543 0 _018_
rlabel metal1 32982 5678 32982 5678 0 _019_
rlabel metal1 28290 3543 28290 3543 0 _020_
rlabel metal1 25990 2455 25990 2455 0 _021_
rlabel metal1 24157 2346 24157 2346 0 _022_
rlabel metal1 32108 2618 32108 2618 0 _023_
rlabel metal2 34086 6052 34086 6052 0 _024_
rlabel metal1 30965 2346 30965 2346 0 _025_
rlabel metal2 34638 3808 34638 3808 0 _026_
rlabel metal1 34730 3706 34730 3706 0 _027_
rlabel via1 30314 4029 30314 4029 0 _028_
rlabel metal1 30137 3094 30137 3094 0 _029_
rlabel metal1 30965 5610 30965 5610 0 _030_
rlabel metal2 32430 3502 32430 3502 0 _031_
rlabel metal1 28757 4590 28757 4590 0 _032_
rlabel metal1 24295 3434 24295 3434 0 _033_
rlabel metal2 28290 2108 28290 2108 0 _034_
rlabel metal1 30597 4182 30597 4182 0 _035_
rlabel metal1 22494 30634 22494 30634 0 _036_
rlabel metal1 32154 7378 32154 7378 0 _037_
rlabel metal1 32476 7854 32476 7854 0 _038_
rlabel via2 33810 4131 33810 4131 0 _039_
rlabel metal1 22356 9690 22356 9690 0 _040_
rlabel metal2 26358 13498 26358 13498 0 _041_
rlabel via2 22218 10693 22218 10693 0 _042_
rlabel metal1 30222 10710 30222 10710 0 _043_
rlabel metal2 22402 11730 22402 11730 0 _044_
rlabel metal1 27094 12104 27094 12104 0 _045_
rlabel metal2 25714 10608 25714 10608 0 _046_
rlabel metal1 26312 8602 26312 8602 0 _047_
rlabel metal1 22494 13192 22494 13192 0 _048_
rlabel metal2 17250 10472 17250 10472 0 _049_
rlabel metal1 20792 12410 20792 12410 0 _050_
rlabel metal1 24012 9146 24012 9146 0 _051_
rlabel metal1 27186 14042 27186 14042 0 _052_
rlabel metal1 26864 15538 26864 15538 0 _053_
rlabel metal1 25852 12954 25852 12954 0 _054_
rlabel metal1 27232 13974 27232 13974 0 _055_
rlabel metal1 27324 14994 27324 14994 0 _056_
rlabel metal1 25806 14450 25806 14450 0 _057_
rlabel metal1 26910 17306 26910 17306 0 _058_
rlabel metal1 24840 15130 24840 15130 0 _059_
rlabel metal2 27922 13634 27922 13634 0 _060_
rlabel metal2 24794 16252 24794 16252 0 _061_
rlabel metal1 24840 15538 24840 15538 0 _062_
rlabel metal1 23460 14042 23460 14042 0 _063_
rlabel metal2 21390 7650 21390 7650 0 _064_
rlabel metal1 21114 6426 21114 6426 0 _065_
rlabel metal1 20746 5202 20746 5202 0 _066_
rlabel metal2 22126 4828 22126 4828 0 _067_
rlabel metal1 23736 11322 23736 11322 0 _068_
rlabel metal2 22218 7446 22218 7446 0 _069_
rlabel metal1 24978 13226 24978 13226 0 _070_
rlabel metal2 23322 11458 23322 11458 0 _071_
rlabel metal1 22034 8840 22034 8840 0 _072_
rlabel metal2 20654 3740 20654 3740 0 _073_
rlabel metal2 23046 11560 23046 11560 0 _074_
rlabel metal2 24702 9758 24702 9758 0 _075_
rlabel metal1 26956 17850 26956 17850 0 _076_
rlabel metal1 27508 15674 27508 15674 0 _077_
rlabel metal1 21689 16490 21689 16490 0 _078_
rlabel metal1 21735 18394 21735 18394 0 _079_
rlabel metal2 21758 18258 21758 18258 0 _080_
rlabel metal1 22310 17850 22310 17850 0 _081_
rlabel metal2 22218 14178 22218 14178 0 _082_
rlabel metal1 22862 17238 22862 17238 0 _083_
rlabel metal1 27876 15130 27876 15130 0 _084_
rlabel metal1 23230 18632 23230 18632 0 _085_
rlabel metal1 26174 18938 26174 18938 0 _086_
rlabel metal1 22862 15130 22862 15130 0 _087_
rlabel metal2 22678 16864 22678 16864 0 _088_
rlabel metal1 25530 23766 25530 23766 0 _089_
rlabel metal1 22632 22202 22632 22202 0 _090_
rlabel metal2 23138 21828 23138 21828 0 _091_
rlabel metal1 24380 18258 24380 18258 0 _092_
rlabel metal1 24564 17306 24564 17306 0 _093_
rlabel metal1 25116 20026 25116 20026 0 _094_
rlabel metal1 25254 22202 25254 22202 0 _095_
rlabel metal2 26910 18632 26910 18632 0 _096_
rlabel metal1 22540 21658 22540 21658 0 _097_
rlabel metal2 23322 19652 23322 19652 0 _098_
rlabel metal2 23690 20264 23690 20264 0 _099_
rlabel metal1 24656 8058 24656 8058 0 _100_
rlabel metal2 26266 9758 26266 9758 0 _101_
rlabel metal2 23966 15096 23966 15096 0 _102_
rlabel metal1 23736 13498 23736 13498 0 _103_
rlabel metal1 25576 15062 25576 15062 0 _104_
rlabel metal2 26726 11322 26726 11322 0 _105_
rlabel metal2 25438 9656 25438 9656 0 _106_
rlabel metal1 26128 12886 26128 12886 0 _107_
rlabel metal1 26864 13498 26864 13498 0 _108_
rlabel metal2 38318 17119 38318 17119 0 ccff_head
rlabel metal2 38226 34221 38226 34221 0 ccff_tail
rlabel metal1 14306 2346 14306 2346 0 chany_bottom_in[0]
rlabel via2 1610 20485 1610 20485 0 chany_bottom_in[10]
rlabel metal2 1702 22559 1702 22559 0 chany_bottom_in[11]
rlabel metal2 38318 5593 38318 5593 0 chany_bottom_in[12]
rlabel metal2 38226 24667 38226 24667 0 chany_bottom_in[13]
rlabel via2 38318 26571 38318 26571 0 chany_bottom_in[14]
rlabel metal1 38272 3026 38272 3026 0 chany_bottom_in[15]
rlabel metal1 20056 37298 20056 37298 0 chany_bottom_in[16]
rlabel via2 1610 32011 1610 32011 0 chany_bottom_in[17]
rlabel metal2 1610 19023 1610 19023 0 chany_bottom_in[18]
rlabel metal1 36202 2414 36202 2414 0 chany_bottom_in[1]
rlabel via2 38318 7531 38318 7531 0 chany_bottom_in[2]
rlabel metal1 9154 2346 9154 2346 0 chany_bottom_in[3]
rlabel metal1 23644 37298 23644 37298 0 chany_bottom_in[4]
rlabel metal2 38318 29903 38318 29903 0 chany_bottom_in[5]
rlabel metal1 34914 2414 34914 2414 0 chany_bottom_in[6]
rlabel metal1 34224 37434 34224 37434 0 chany_bottom_in[7]
rlabel metal1 35880 3026 35880 3026 0 chany_bottom_in[8]
rlabel metal1 26864 37434 26864 37434 0 chany_bottom_in[9]
rlabel metal1 7222 37094 7222 37094 0 chany_bottom_out[0]
rlabel metal1 18216 37094 18216 37094 0 chany_bottom_out[10]
rlabel metal3 1188 24548 1188 24548 0 chany_bottom_out[11]
rlabel metal2 38226 13073 38226 13073 0 chany_bottom_out[12]
rlabel metal3 1188 7548 1188 7548 0 chany_bottom_out[13]
rlabel metal3 1188 30668 1188 30668 0 chany_bottom_out[14]
rlabel metal3 1188 3468 1188 3468 0 chany_bottom_out[15]
rlabel metal3 1188 15028 1188 15028 0 chany_bottom_out[16]
rlabel metal2 38226 28815 38226 28815 0 chany_bottom_out[17]
rlabel metal2 38226 15181 38226 15181 0 chany_bottom_out[18]
rlabel metal1 21758 37094 21758 37094 0 chany_bottom_out[1]
rlabel metal2 38226 36057 38226 36057 0 chany_bottom_out[2]
rlabel metal1 2668 37094 2668 37094 0 chany_bottom_out[3]
rlabel metal1 29486 37094 29486 37094 0 chany_bottom_out[4]
rlabel metal3 1188 10948 1188 10948 0 chany_bottom_out[5]
rlabel metal1 1518 37094 1518 37094 0 chany_bottom_out[6]
rlabel metal1 38134 37094 38134 37094 0 chany_bottom_out[7]
rlabel metal3 1188 34068 1188 34068 0 chany_bottom_out[8]
rlabel metal1 25576 2822 25576 2822 0 chany_bottom_out[9]
rlabel via2 38318 32011 38318 32011 0 chany_top_in[0]
rlabel metal1 10764 37298 10764 37298 0 chany_top_in[10]
rlabel metal1 3680 2346 3680 2346 0 chany_top_in[11]
rlabel metal1 10764 2482 10764 2482 0 chany_top_in[12]
rlabel metal2 32522 3468 32522 3468 0 chany_top_in[13]
rlabel metal2 38318 10863 38318 10863 0 chany_top_in[14]
rlabel via2 38318 3485 38318 3485 0 chany_top_in[15]
rlabel metal1 22908 3026 22908 3026 0 chany_top_in[16]
rlabel metal1 874 36822 874 36822 0 chany_top_in[17]
rlabel metal2 38042 1588 38042 1588 0 chany_top_in[18]
rlabel metal1 12328 37298 12328 37298 0 chany_top_in[1]
rlabel via2 38226 8891 38226 8891 0 chany_top_in[2]
rlabel metal2 1610 1921 1610 1921 0 chany_top_in[3]
rlabel metal2 29026 1435 29026 1435 0 chany_top_in[4]
rlabel via2 1610 26571 1610 26571 0 chany_top_in[5]
rlabel via2 1610 9605 1610 9605 0 chany_top_in[6]
rlabel metal1 16721 37298 16721 37298 0 chany_top_in[7]
rlabel metal1 18170 2414 18170 2414 0 chany_top_in[8]
rlabel metal1 828 2958 828 2958 0 chany_top_in[9]
rlabel metal3 1188 17068 1188 17068 0 chany_top_out[0]
rlabel metal1 14352 37094 14352 37094 0 chany_top_out[10]
rlabel metal1 25300 37094 25300 37094 0 chany_top_out[11]
rlabel metal1 36202 37094 36202 37094 0 chany_top_out[12]
rlabel metal3 1188 28628 1188 28628 0 chany_top_out[13]
rlabel metal2 5198 1520 5198 1520 0 chany_top_out[14]
rlabel metal2 1334 1520 1334 1520 0 chany_top_out[15]
rlabel metal1 38778 36890 38778 36890 0 chany_top_out[16]
rlabel metal1 30544 37094 30544 37094 0 chany_top_out[17]
rlabel metal2 16146 1520 16146 1520 0 chany_top_out[18]
rlabel metal3 38786 38148 38786 38148 0 chany_top_out[1]
rlabel metal3 38234 1428 38234 1428 0 chany_top_out[2]
rlabel metal1 5290 37094 5290 37094 0 chany_top_out[3]
rlabel metal2 38226 20621 38226 20621 0 chany_top_out[4]
rlabel metal2 7130 1520 7130 1520 0 chany_top_out[5]
rlabel metal2 12282 1520 12282 1520 0 chany_top_out[6]
rlabel metal2 19366 1520 19366 1520 0 chany_top_out[7]
rlabel via2 38226 22491 38226 22491 0 chany_top_out[8]
rlabel metal2 21298 1520 21298 1520 0 chany_top_out[9]
rlabel metal3 1188 5508 1188 5508 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
rlabel metal1 32384 37094 32384 37094 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
rlabel metal1 3726 37094 3726 37094 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
rlabel metal1 20746 12206 20746 12206 0 mem_left_ipin_0.DFFR_0_.Q
rlabel metal1 27186 12750 27186 12750 0 mem_left_ipin_0.DFFR_1_.Q
rlabel metal1 21482 10608 21482 10608 0 mem_left_ipin_0.DFFR_2_.Q
rlabel metal1 26910 8398 26910 8398 0 mem_left_ipin_0.DFFR_3_.Q
rlabel metal1 30452 8398 30452 8398 0 mem_left_ipin_0.DFFR_4_.Q
rlabel metal1 29486 8330 29486 8330 0 mem_left_ipin_0.DFFR_5_.Q
rlabel metal1 24702 16558 24702 16558 0 mem_left_ipin_1.DFFR_0_.Q
rlabel metal2 25898 15198 25898 15198 0 mem_left_ipin_1.DFFR_1_.Q
rlabel metal1 27416 16558 27416 16558 0 mem_left_ipin_1.DFFR_2_.Q
rlabel metal1 28612 12886 28612 12886 0 mem_left_ipin_1.DFFR_3_.Q
rlabel metal1 27462 13906 27462 13906 0 mem_left_ipin_1.DFFR_4_.Q
rlabel metal1 29808 5338 29808 5338 0 mem_left_ipin_1.DFFR_5_.Q
rlabel metal1 28060 2482 28060 2482 0 mem_left_ipin_2.DFFR_0_.Q
rlabel metal1 26404 14994 26404 14994 0 mem_left_ipin_2.DFFR_1_.Q
rlabel metal1 24978 13158 24978 13158 0 mem_left_ipin_2.DFFR_2_.Q
rlabel metal2 31878 3077 31878 3077 0 mem_left_ipin_2.DFFR_3_.Q
rlabel metal2 32338 4284 32338 4284 0 mem_left_ipin_2.DFFR_4_.Q
rlabel metal1 29072 8534 29072 8534 0 mem_left_ipin_2.DFFR_5_.Q
rlabel metal1 21114 4046 21114 4046 0 mem_right_ipin_0.DFFR_0_.Q
rlabel metal1 21206 5236 21206 5236 0 mem_right_ipin_0.DFFR_1_.Q
rlabel metal1 22586 8466 22586 8466 0 mem_right_ipin_0.DFFR_2_.Q
rlabel metal2 24058 6188 24058 6188 0 mem_right_ipin_0.DFFR_3_.Q
rlabel metal1 21482 7412 21482 7412 0 mem_right_ipin_0.DFFR_4_.Q
rlabel metal1 21482 6358 21482 6358 0 mem_right_ipin_0.DFFR_5_.Q
rlabel metal1 22724 2482 22724 2482 0 mem_right_ipin_1.DFFR_0_.Q
rlabel metal1 23644 2278 23644 2278 0 mem_right_ipin_1.DFFR_1_.Q
rlabel metal1 26772 2482 26772 2482 0 mem_right_ipin_1.DFFR_2_.Q
rlabel metal1 28520 14994 28520 14994 0 mem_right_ipin_1.DFFR_3_.Q
rlabel metal1 32062 3604 32062 3604 0 mem_right_ipin_1.DFFR_4_.Q
rlabel metal1 34868 3638 34868 3638 0 mem_right_ipin_1.DFFR_5_.Q
rlabel metal1 23552 19346 23552 19346 0 mem_right_ipin_2.DFFR_0_.Q
rlabel metal1 25484 18734 25484 18734 0 mem_right_ipin_2.DFFR_1_.Q
rlabel metal1 24334 17170 24334 17170 0 mem_right_ipin_2.DFFR_2_.Q
rlabel metal2 36662 3145 36662 3145 0 mem_right_ipin_2.DFFR_3_.Q
rlabel metal2 21482 15844 21482 15844 0 mem_right_ipin_2.DFFR_4_.Q
rlabel metal1 22908 13362 22908 13362 0 mux_left_ipin_0.INVTX1_0_.out
rlabel metal1 25300 31110 25300 31110 0 mux_left_ipin_0.INVTX1_1_.out
rlabel metal2 22310 9554 22310 9554 0 mux_left_ipin_0.INVTX1_2_.out
rlabel metal2 14398 10404 14398 10404 0 mux_left_ipin_0.INVTX1_3_.out
rlabel metal2 33626 10404 33626 10404 0 mux_left_ipin_0.INVTX1_4_.out
rlabel metal1 22028 10710 22028 10710 0 mux_left_ipin_0.INVTX1_5_.out
rlabel metal1 18998 12274 18998 12274 0 mux_left_ipin_0.INVTX1_6_.out
rlabel metal1 28106 12614 28106 12614 0 mux_left_ipin_0.INVTX1_7_.out
rlabel metal1 23736 13430 23736 13430 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 26634 10302 26634 10302 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 21850 12750 21850 12750 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 2300 35666 2300 35666 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 27692 14926 27692 14926 0 mux_left_ipin_1.INVTX1_2_.out
rlabel metal1 23046 29002 23046 29002 0 mux_left_ipin_1.INVTX1_3_.out
rlabel metal1 22954 16116 22954 16116 0 mux_left_ipin_1.INVTX1_4_.out
rlabel metal1 25668 27846 25668 27846 0 mux_left_ipin_1.INVTX1_5_.out
rlabel metal2 24610 18700 24610 18700 0 mux_left_ipin_1.INVTX1_6_.out
rlabel metal1 25944 11866 25944 11866 0 mux_left_ipin_1.INVTX1_7_.out
rlabel metal1 24426 14382 24426 14382 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 26128 16014 26128 16014 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 25714 15708 25714 15708 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 26680 16082 26680 16082 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 24794 9452 24794 9452 0 mux_left_ipin_2.INVTX1_2_.out
rlabel metal1 25070 12716 25070 12716 0 mux_left_ipin_2.INVTX1_3_.out
rlabel metal2 23782 19244 23782 19244 0 mux_left_ipin_2.INVTX1_4_.out
rlabel metal1 21252 16626 21252 16626 0 mux_left_ipin_2.INVTX1_5_.out
rlabel metal1 25852 14926 25852 14926 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 24058 15504 24058 15504 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 5014 11696 5014 11696 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 16560 14280 16560 14280 0 mux_right_ipin_0.INVTX1_2_.out
rlabel metal2 10626 13056 10626 13056 0 mux_right_ipin_0.INVTX1_3_.out
rlabel metal1 23276 12682 23276 12682 0 mux_right_ipin_0.INVTX1_4_.out
rlabel metal2 22126 5780 22126 5780 0 mux_right_ipin_0.INVTX1_5_.out
rlabel metal2 21390 3332 21390 3332 0 mux_right_ipin_0.INVTX1_6_.out
rlabel metal1 20470 4250 20470 4250 0 mux_right_ipin_0.INVTX1_7_.out
rlabel metal2 24150 9248 24150 9248 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 23092 12750 23092 12750 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 20562 5066 20562 5066 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 5382 5678 5382 5678 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 23414 18734 23414 18734 0 mux_right_ipin_1.INVTX1_2_.out
rlabel metal2 26450 19822 26450 19822 0 mux_right_ipin_1.INVTX1_3_.out
rlabel metal1 20470 18802 20470 18802 0 mux_right_ipin_1.INVTX1_4_.out
rlabel metal1 21022 19346 21022 19346 0 mux_right_ipin_1.INVTX1_5_.out
rlabel metal1 23000 30566 23000 30566 0 mux_right_ipin_1.INVTX1_6_.out
rlabel metal1 22402 15674 22402 15674 0 mux_right_ipin_1.INVTX1_7_.out
rlabel metal2 23138 14994 23138 14994 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 25438 18768 25438 18768 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 23138 17442 23138 17442 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 30038 36788 30038 36788 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 25530 22814 25530 22814 0 mux_right_ipin_2.INVTX1_2_.out
rlabel metal2 22494 19346 22494 19346 0 mux_right_ipin_2.INVTX1_3_.out
rlabel metal1 22448 23698 22448 23698 0 mux_right_ipin_2.INVTX1_6_.out
rlabel metal1 22632 26282 22632 26282 0 mux_right_ipin_2.INVTX1_7_.out
rlabel metal1 24518 20366 24518 20366 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 23276 17714 23276 17714 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 23506 23698 23506 23698 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 4508 36550 4508 36550 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 38042 16966 38042 16966 0 net1
rlabel metal1 24380 36754 24380 36754 0 net10
rlabel metal1 17480 12206 17480 12206 0 net11
rlabel metal1 36892 2550 36892 2550 0 net12
rlabel metal1 37950 7922 37950 7922 0 net13
rlabel metal1 10764 2550 10764 2550 0 net14
rlabel metal1 24610 37196 24610 37196 0 net15
rlabel metal1 25714 23698 25714 23698 0 net16
rlabel metal1 18216 2822 18216 2822 0 net17
rlabel metal1 34868 37298 34868 37298 0 net18
rlabel metal1 35466 14382 35466 14382 0 net19
rlabel metal1 19504 13906 19504 13906 0 net2
rlabel metal1 21758 11730 21758 11730 0 net20
rlabel metal2 25530 31858 25530 31858 0 net21
rlabel metal1 18262 30226 18262 30226 0 net22
rlabel metal1 2530 21998 2530 21998 0 net23
rlabel metal1 21344 11118 21344 11118 0 net24
rlabel metal1 14582 7378 14582 7378 0 net25
rlabel metal1 19918 20842 19918 20842 0 net26
rlabel metal1 20424 4114 20424 4114 0 net27
rlabel metal1 12650 14994 12650 14994 0 net28
rlabel metal1 2070 36618 2070 36618 0 net29
rlabel metal2 16606 20332 16606 20332 0 net3
rlabel metal1 37812 13906 37812 13906 0 net30
rlabel metal2 20746 37026 20746 37026 0 net31
rlabel metal1 37996 18734 37996 18734 0 net32
rlabel metal1 1932 2482 1932 2482 0 net33
rlabel metal1 28336 23698 28336 23698 0 net34
rlabel metal1 2346 16762 2346 16762 0 net35
rlabel metal2 1886 10370 1886 10370 0 net36
rlabel metal1 21298 36686 21298 36686 0 net37
rlabel metal1 11224 2346 11224 2346 0 net38
rlabel metal1 22264 5202 22264 5202 0 net39
rlabel metal2 1886 21352 1886 21352 0 net4
rlabel metal1 10166 30702 10166 30702 0 net40
rlabel metal1 37766 34578 37766 34578 0 net41
rlabel metal1 7774 37230 7774 37230 0 net42
rlabel metal2 17894 37060 17894 37060 0 net43
rlabel metal2 2070 23324 2070 23324 0 net44
rlabel metal2 38042 12444 38042 12444 0 net45
rlabel metal2 14122 7684 14122 7684 0 net46
rlabel metal1 2116 30702 2116 30702 0 net47
rlabel metal1 4393 3502 4393 3502 0 net48
rlabel metal1 4393 15470 4393 15470 0 net49
rlabel metal2 36202 8262 36202 8262 0 net5
rlabel metal1 23230 28424 23230 28424 0 net50
rlabel metal2 38042 14756 38042 14756 0 net51
rlabel metal2 21390 37060 21390 37060 0 net52
rlabel metal1 37904 18938 37904 18938 0 net53
rlabel metal1 1932 36550 1932 36550 0 net54
rlabel metal1 29256 37230 29256 37230 0 net55
rlabel metal2 1794 13770 1794 13770 0 net56
rlabel metal1 1886 37196 1886 37196 0 net57
rlabel metal1 26174 36652 26174 36652 0 net58
rlabel metal1 2254 34510 2254 34510 0 net59
rlabel metal1 20470 26418 20470 26418 0 net6
rlabel metal1 25806 2992 25806 2992 0 net60
rlabel metal1 4370 17170 4370 17170 0 net61
rlabel metal1 14260 29274 14260 29274 0 net62
rlabel metal1 24288 37094 24288 37094 0 net63
rlabel metal1 36432 36550 36432 36550 0 net64
rlabel metal2 1886 27778 1886 27778 0 net65
rlabel metal2 5566 2652 5566 2652 0 net66
rlabel metal2 3174 2754 3174 2754 0 net67
rlabel metal1 38042 36686 38042 36686 0 net68
rlabel metal2 24242 36448 24242 36448 0 net69
rlabel metal2 37950 19516 37950 19516 0 net7
rlabel metal1 16422 2414 16422 2414 0 net70
rlabel metal1 37996 20570 37996 20570 0 net71
rlabel metal2 38042 4284 38042 4284 0 net72
rlabel metal2 5566 30260 5566 30260 0 net73
rlabel metal1 36961 20910 36961 20910 0 net74
rlabel metal1 7728 2414 7728 2414 0 net75
rlabel metal2 14582 2618 14582 2618 0 net76
rlabel metal1 20792 2482 20792 2482 0 net77
rlabel metal1 36892 22610 36892 22610 0 net78
rlabel metal1 21252 11526 21252 11526 0 net79
rlabel via2 21482 3043 21482 3043 0 net8
rlabel metal1 3450 5678 3450 5678 0 net80
rlabel metal1 31234 36890 31234 36890 0 net81
rlabel metal2 3450 37060 3450 37060 0 net82
rlabel metal1 4508 12410 4508 12410 0 net83
rlabel metal1 1932 35802 1932 35802 0 net84
rlabel metal2 33166 18598 33166 18598 0 net85
rlabel metal1 21758 12138 21758 12138 0 net86
rlabel metal2 26358 16286 26358 16286 0 net87
rlabel metal2 22218 5066 22218 5066 0 net88
rlabel metal2 22678 18394 22678 18394 0 net89
rlabel metal1 22356 37162 22356 37162 0 net9
rlabel metal1 23000 22066 23000 22066 0 net90
rlabel metal1 26404 9010 26404 9010 0 net91
rlabel metal1 9108 37230 9108 37230 0 pReset
rlabel metal1 22264 3502 22264 3502 0 prog_clk
rlabel metal3 1188 12988 1188 12988 0 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
rlabel metal3 1188 36108 1188 36108 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
rlabel via2 38226 19125 38226 19125 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
