magic
tech sky130A
magscale 1 2
timestamp 1672417504
<< viali >>
rect 36093 37417 36127 37451
rect 37473 37281 37507 37315
rect 1593 37213 1627 37247
rect 2513 37213 2547 37247
rect 3157 37213 3191 37247
rect 4169 37213 4203 37247
rect 5457 37213 5491 37247
rect 7389 37213 7423 37247
rect 9321 37213 9355 37247
rect 10609 37213 10643 37247
rect 11897 37213 11931 37247
rect 13001 37213 13035 37247
rect 15117 37213 15151 37247
rect 17049 37213 17083 37247
rect 18153 37213 18187 37247
rect 19441 37213 19475 37247
rect 20729 37213 20763 37247
rect 22845 37213 22879 37247
rect 24593 37213 24627 37247
rect 26065 37213 26099 37247
rect 27169 37213 27203 37247
rect 29929 37213 29963 37247
rect 30573 37213 30607 37247
rect 32505 37213 32539 37247
rect 33793 37213 33827 37247
rect 35081 37213 35115 37247
rect 35909 37213 35943 37247
rect 36645 37213 36679 37247
rect 37749 37213 37783 37247
rect 1777 37077 1811 37111
rect 2329 37077 2363 37111
rect 2973 37077 3007 37111
rect 3985 37077 4019 37111
rect 5273 37077 5307 37111
rect 7205 37077 7239 37111
rect 9137 37077 9171 37111
rect 10425 37077 10459 37111
rect 11713 37077 11747 37111
rect 13185 37077 13219 37111
rect 14933 37077 14967 37111
rect 16865 37077 16899 37111
rect 18337 37077 18371 37111
rect 19625 37077 19659 37111
rect 20913 37077 20947 37111
rect 22661 37077 22695 37111
rect 24777 37077 24811 37111
rect 25881 37077 25915 37111
rect 27353 37077 27387 37111
rect 29745 37077 29779 37111
rect 30389 37077 30423 37111
rect 32321 37077 32355 37111
rect 33609 37077 33643 37111
rect 34897 37077 34931 37111
rect 36829 37077 36863 37111
rect 1777 36873 1811 36907
rect 34161 36873 34195 36907
rect 38209 36873 38243 36907
rect 1593 36737 1627 36771
rect 34345 36737 34379 36771
rect 38025 36737 38059 36771
rect 30297 36329 30331 36363
rect 38209 36329 38243 36363
rect 1777 36125 1811 36159
rect 30481 36125 30515 36159
rect 38025 36125 38059 36159
rect 1593 35989 1627 36023
rect 33425 35785 33459 35819
rect 33333 35649 33367 35683
rect 38301 35037 38335 35071
rect 38117 34901 38151 34935
rect 1777 34697 1811 34731
rect 37473 34697 37507 34731
rect 1961 34561 1995 34595
rect 15301 34561 15335 34595
rect 37657 34561 37691 34595
rect 15393 34493 15427 34527
rect 34897 34153 34931 34187
rect 1777 33949 1811 33983
rect 12817 33949 12851 33983
rect 13461 33949 13495 33983
rect 35081 33949 35115 33983
rect 1593 33813 1627 33847
rect 12633 33813 12667 33847
rect 13277 33813 13311 33847
rect 14289 33813 14323 33847
rect 1961 33609 1995 33643
rect 17233 33609 17267 33643
rect 23305 33609 23339 33643
rect 1869 33473 1903 33507
rect 2513 33473 2547 33507
rect 11713 33473 11747 33507
rect 13553 33473 13587 33507
rect 13737 33473 13771 33507
rect 17417 33473 17451 33507
rect 23489 33473 23523 33507
rect 38301 33473 38335 33507
rect 2605 33269 2639 33303
rect 11805 33269 11839 33303
rect 13921 33269 13955 33303
rect 38117 33269 38151 33303
rect 2881 33065 2915 33099
rect 23121 33065 23155 33099
rect 14749 32997 14783 33031
rect 4077 32929 4111 32963
rect 1777 32861 1811 32895
rect 3065 32861 3099 32895
rect 3985 32861 4019 32895
rect 9137 32861 9171 32895
rect 14933 32861 14967 32895
rect 15577 32861 15611 32895
rect 23305 32861 23339 32895
rect 1593 32725 1627 32759
rect 9229 32725 9263 32759
rect 15393 32725 15427 32759
rect 16037 32725 16071 32759
rect 12357 32521 12391 32555
rect 18981 32521 19015 32555
rect 19717 32521 19751 32555
rect 7205 32453 7239 32487
rect 1869 32385 1903 32419
rect 4629 32385 4663 32419
rect 6561 32385 6595 32419
rect 7665 32385 7699 32419
rect 10333 32385 10367 32419
rect 11069 32385 11103 32419
rect 11713 32385 11747 32419
rect 11897 32385 11931 32419
rect 13369 32385 13403 32419
rect 14197 32385 14231 32419
rect 14749 32385 14783 32419
rect 15669 32385 15703 32419
rect 15853 32385 15887 32419
rect 17049 32385 17083 32419
rect 19165 32385 19199 32419
rect 19625 32385 19659 32419
rect 27629 32385 27663 32419
rect 4721 32317 4755 32351
rect 5273 32317 5307 32351
rect 5457 32317 5491 32351
rect 6745 32317 6779 32351
rect 5917 32249 5951 32283
rect 10885 32249 10919 32283
rect 1961 32181 1995 32215
rect 7757 32181 7791 32215
rect 10149 32181 10183 32215
rect 13461 32181 13495 32215
rect 14013 32181 14047 32215
rect 14841 32181 14875 32215
rect 16037 32181 16071 32215
rect 16865 32181 16899 32215
rect 27721 32181 27755 32215
rect 5089 31977 5123 32011
rect 11529 31977 11563 32011
rect 13461 31977 13495 32011
rect 2053 31909 2087 31943
rect 2697 31909 2731 31943
rect 12173 31909 12207 31943
rect 14841 31909 14875 31943
rect 9781 31841 9815 31875
rect 12817 31841 12851 31875
rect 21373 31841 21407 31875
rect 25973 31841 26007 31875
rect 38301 31841 38335 31875
rect 2237 31773 2271 31807
rect 2881 31773 2915 31807
rect 5273 31773 5307 31807
rect 9689 31773 9723 31807
rect 11713 31773 11747 31807
rect 12357 31773 12391 31807
rect 13001 31773 13035 31807
rect 15025 31773 15059 31807
rect 16405 31773 16439 31807
rect 16497 31773 16531 31807
rect 17417 31773 17451 31807
rect 20729 31773 20763 31807
rect 20913 31773 20947 31807
rect 25881 31773 25915 31807
rect 38117 31773 38151 31807
rect 17233 31637 17267 31671
rect 4997 31433 5031 31467
rect 6653 31433 6687 31467
rect 19901 31433 19935 31467
rect 20729 31433 20763 31467
rect 22293 31433 22327 31467
rect 22937 31433 22971 31467
rect 9413 31365 9447 31399
rect 16957 31365 16991 31399
rect 17049 31365 17083 31399
rect 2145 31297 2179 31331
rect 5181 31297 5215 31331
rect 6561 31297 6595 31331
rect 8585 31297 8619 31331
rect 10701 31297 10735 31331
rect 12265 31297 12299 31331
rect 13645 31297 13679 31331
rect 14105 31297 14139 31331
rect 16037 31297 16071 31331
rect 19809 31297 19843 31331
rect 22477 31297 22511 31331
rect 23121 31297 23155 31331
rect 7389 31229 7423 31263
rect 7573 31229 7607 31263
rect 8677 31229 8711 31263
rect 9321 31229 9355 31263
rect 14197 31229 14231 31263
rect 14933 31229 14967 31263
rect 17601 31229 17635 31263
rect 9873 31161 9907 31195
rect 13461 31161 13495 31195
rect 1961 31093 1995 31127
rect 7757 31093 7791 31127
rect 10517 31093 10551 31127
rect 12357 31093 12391 31127
rect 16129 31093 16163 31127
rect 1961 30889 1995 30923
rect 7757 30889 7791 30923
rect 9229 30889 9263 30923
rect 13461 30889 13495 30923
rect 20821 30889 20855 30923
rect 22845 30889 22879 30923
rect 8401 30821 8435 30855
rect 15025 30821 15059 30855
rect 6561 30753 6595 30787
rect 11345 30753 11379 30787
rect 11989 30753 12023 30787
rect 15577 30753 15611 30787
rect 15761 30753 15795 30787
rect 23397 30753 23431 30787
rect 2145 30685 2179 30719
rect 2605 30685 2639 30719
rect 3249 30685 3283 30719
rect 3985 30685 4019 30719
rect 7941 30685 7975 30719
rect 8585 30685 8619 30719
rect 9413 30685 9447 30719
rect 9873 30685 9907 30719
rect 10609 30685 10643 30719
rect 13369 30685 13403 30719
rect 17141 30685 17175 30719
rect 19717 30685 19751 30719
rect 20361 30685 20395 30719
rect 21005 30685 21039 30719
rect 22753 30685 22787 30719
rect 23581 30685 23615 30719
rect 28273 30685 28307 30719
rect 6653 30617 6687 30651
rect 7205 30617 7239 30651
rect 9965 30617 9999 30651
rect 11437 30617 11471 30651
rect 14473 30617 14507 30651
rect 14565 30617 14599 30651
rect 2697 30549 2731 30583
rect 3341 30549 3375 30583
rect 4169 30549 4203 30583
rect 10701 30549 10735 30583
rect 16221 30549 16255 30583
rect 16957 30549 16991 30583
rect 19533 30549 19567 30583
rect 20177 30549 20211 30583
rect 24041 30549 24075 30583
rect 28365 30549 28399 30583
rect 3985 30277 4019 30311
rect 7021 30277 7055 30311
rect 10885 30277 10919 30311
rect 17049 30277 17083 30311
rect 17601 30277 17635 30311
rect 31585 30277 31619 30311
rect 1777 30209 1811 30243
rect 2697 30209 2731 30243
rect 2789 30209 2823 30243
rect 3525 30209 3559 30243
rect 6009 30209 6043 30243
rect 9229 30209 9263 30243
rect 10793 30209 10827 30243
rect 12449 30209 12483 30243
rect 13185 30209 13219 30243
rect 13829 30209 13863 30243
rect 18061 30209 18095 30243
rect 22017 30209 22051 30243
rect 31493 30209 31527 30243
rect 33333 30209 33367 30243
rect 33425 30209 33459 30243
rect 34345 30209 34379 30243
rect 38025 30209 38059 30243
rect 3341 30141 3375 30175
rect 4445 30141 4479 30175
rect 6929 30141 6963 30175
rect 16957 30141 16991 30175
rect 7481 30073 7515 30107
rect 34161 30073 34195 30107
rect 1593 30005 1627 30039
rect 5825 30005 5859 30039
rect 9321 30005 9355 30039
rect 12265 30005 12299 30039
rect 13277 30005 13311 30039
rect 13921 30005 13955 30039
rect 18153 30005 18187 30039
rect 22109 30005 22143 30039
rect 38209 30005 38243 30039
rect 6193 29801 6227 29835
rect 6929 29801 6963 29835
rect 18797 29801 18831 29835
rect 21833 29801 21867 29835
rect 23121 29801 23155 29835
rect 23857 29801 23891 29835
rect 4077 29733 4111 29767
rect 2789 29665 2823 29699
rect 3065 29665 3099 29699
rect 9321 29665 9355 29699
rect 11529 29665 11563 29699
rect 12541 29665 12575 29699
rect 19441 29665 19475 29699
rect 19625 29665 19659 29699
rect 21649 29665 21683 29699
rect 1869 29597 1903 29631
rect 3985 29597 4019 29631
rect 6377 29597 6411 29631
rect 6837 29597 6871 29631
rect 7481 29597 7515 29631
rect 9137 29597 9171 29631
rect 11345 29597 11379 29631
rect 14289 29597 14323 29631
rect 17325 29597 17359 29631
rect 18705 29597 18739 29631
rect 20821 29597 20855 29631
rect 21465 29597 21499 29631
rect 23029 29597 23063 29631
rect 23765 29597 23799 29631
rect 2881 29529 2915 29563
rect 12633 29529 12667 29563
rect 13185 29529 13219 29563
rect 1961 29461 1995 29495
rect 7573 29461 7607 29495
rect 9781 29461 9815 29495
rect 11989 29461 12023 29495
rect 14381 29461 14415 29495
rect 17141 29461 17175 29495
rect 20085 29461 20119 29495
rect 20913 29461 20947 29495
rect 5273 29257 5307 29291
rect 12357 29257 12391 29291
rect 13645 29257 13679 29291
rect 30481 29257 30515 29291
rect 10609 29189 10643 29223
rect 1777 29121 1811 29155
rect 5181 29121 5215 29155
rect 6653 29121 6687 29155
rect 7665 29121 7699 29155
rect 9873 29121 9907 29155
rect 12541 29121 12575 29155
rect 13185 29121 13219 29155
rect 15209 29121 15243 29155
rect 16221 29121 16255 29155
rect 18981 29121 19015 29155
rect 25329 29121 25363 29155
rect 30389 29121 30423 29155
rect 38025 29121 38059 29155
rect 6745 29053 6779 29087
rect 10517 29053 10551 29087
rect 10793 29053 10827 29087
rect 13001 29053 13035 29087
rect 18797 29053 18831 29087
rect 23397 29053 23431 29087
rect 24041 29053 24075 29087
rect 24225 29053 24259 29087
rect 7481 28985 7515 29019
rect 9689 28985 9723 29019
rect 19165 28985 19199 29019
rect 38209 28985 38243 29019
rect 1593 28917 1627 28951
rect 15025 28917 15059 28951
rect 16037 28917 16071 28951
rect 24685 28917 24719 28951
rect 25145 28917 25179 28951
rect 10609 28713 10643 28747
rect 16865 28713 16899 28747
rect 20085 28713 20119 28747
rect 24777 28713 24811 28747
rect 9781 28645 9815 28679
rect 9229 28577 9263 28611
rect 14657 28577 14691 28611
rect 15761 28577 15795 28611
rect 15945 28577 15979 28611
rect 19625 28577 19659 28611
rect 1961 28509 1995 28543
rect 4905 28509 4939 28543
rect 5365 28509 5399 28543
rect 10517 28509 10551 28543
rect 17049 28509 17083 28543
rect 19809 28509 19843 28543
rect 22017 28509 22051 28543
rect 24961 28509 24995 28543
rect 9321 28441 9355 28475
rect 14749 28441 14783 28475
rect 15301 28441 15335 28475
rect 1777 28373 1811 28407
rect 4721 28373 4755 28407
rect 5457 28373 5491 28407
rect 16405 28373 16439 28407
rect 21189 28373 21223 28407
rect 21833 28373 21867 28407
rect 14841 28169 14875 28203
rect 17509 28169 17543 28203
rect 19441 28169 19475 28203
rect 21465 28169 21499 28203
rect 24317 28169 24351 28203
rect 25697 28169 25731 28203
rect 3157 28101 3191 28135
rect 3709 28101 3743 28135
rect 4353 28101 4387 28135
rect 4905 28101 4939 28135
rect 13369 28101 13403 28135
rect 18245 28101 18279 28135
rect 1869 28033 1903 28067
rect 5549 28033 5583 28067
rect 15025 28033 15059 28067
rect 15669 28033 15703 28067
rect 16129 28033 16163 28067
rect 16865 28033 16899 28067
rect 17049 28033 17083 28067
rect 19349 28033 19383 28067
rect 20821 28033 20855 28067
rect 21005 28033 21039 28067
rect 22017 28033 22051 28067
rect 23029 28033 23063 28067
rect 25053 28033 25087 28067
rect 3065 27965 3099 27999
rect 4261 27965 4295 27999
rect 6561 27965 6595 27999
rect 13277 27965 13311 27999
rect 18153 27965 18187 27999
rect 18429 27965 18463 27999
rect 23673 27965 23707 27999
rect 23857 27965 23891 27999
rect 25237 27965 25271 27999
rect 13829 27897 13863 27931
rect 15485 27897 15519 27931
rect 1961 27829 1995 27863
rect 5365 27829 5399 27863
rect 16221 27829 16255 27863
rect 22109 27829 22143 27863
rect 22845 27829 22879 27863
rect 11240 27625 11274 27659
rect 21373 27625 21407 27659
rect 24685 27625 24719 27659
rect 25329 27625 25363 27659
rect 1593 27557 1627 27591
rect 12725 27557 12759 27591
rect 19809 27557 19843 27591
rect 20545 27557 20579 27591
rect 23397 27557 23431 27591
rect 4721 27489 4755 27523
rect 5825 27489 5859 27523
rect 18245 27489 18279 27523
rect 19441 27489 19475 27523
rect 1777 27421 1811 27455
rect 10977 27421 11011 27455
rect 16405 27421 16439 27455
rect 17049 27421 17083 27455
rect 17509 27421 17543 27455
rect 19625 27421 19659 27455
rect 20729 27421 20763 27455
rect 21557 27421 21591 27455
rect 23581 27421 23615 27455
rect 24593 27421 24627 27455
rect 25237 27421 25271 27455
rect 26065 27421 26099 27455
rect 26525 27421 26559 27455
rect 27445 27421 27479 27455
rect 4077 27353 4111 27387
rect 4169 27353 4203 27387
rect 5917 27353 5951 27387
rect 6469 27353 6503 27387
rect 17601 27353 17635 27387
rect 27537 27353 27571 27387
rect 16221 27285 16255 27319
rect 16865 27285 16899 27319
rect 25881 27285 25915 27319
rect 26617 27285 26651 27319
rect 4353 27081 4387 27115
rect 19349 27081 19383 27115
rect 8309 27013 8343 27047
rect 11989 27013 12023 27047
rect 12541 27013 12575 27047
rect 24777 27013 24811 27047
rect 1869 26945 1903 26979
rect 4261 26945 4295 26979
rect 16129 26945 16163 26979
rect 19533 26945 19567 26979
rect 20269 26945 20303 26979
rect 21005 26945 21039 26979
rect 27537 26945 27571 26979
rect 38301 26945 38335 26979
rect 8033 26877 8067 26911
rect 10057 26877 10091 26911
rect 11897 26877 11931 26911
rect 13001 26877 13035 26911
rect 13277 26877 13311 26911
rect 17325 26877 17359 26911
rect 24685 26877 24719 26911
rect 24961 26877 24995 26911
rect 1869 26741 1903 26775
rect 14749 26741 14783 26775
rect 16221 26741 16255 26775
rect 20085 26741 20119 26775
rect 21097 26741 21131 26775
rect 27629 26741 27663 26775
rect 38117 26741 38151 26775
rect 2513 26537 2547 26571
rect 5641 26537 5675 26571
rect 6180 26537 6214 26571
rect 26249 26537 26283 26571
rect 16497 26469 16531 26503
rect 20085 26469 20119 26503
rect 22569 26469 22603 26503
rect 24593 26469 24627 26503
rect 1869 26401 1903 26435
rect 2053 26401 2087 26435
rect 5917 26401 5951 26435
rect 9413 26401 9447 26435
rect 11897 26401 11931 26435
rect 14289 26401 14323 26435
rect 14565 26401 14599 26435
rect 17325 26401 17359 26435
rect 17601 26401 17635 26435
rect 19533 26401 19567 26435
rect 20637 26401 20671 26435
rect 20821 26401 20855 26435
rect 27905 26401 27939 26435
rect 28089 26401 28123 26435
rect 29101 26401 29135 26435
rect 3157 26333 3191 26367
rect 7941 26333 7975 26367
rect 16681 26333 16715 26367
rect 21281 26333 21315 26367
rect 21925 26333 21959 26367
rect 22109 26333 22143 26367
rect 24777 26333 24811 26367
rect 26433 26333 26467 26367
rect 29009 26333 29043 26367
rect 9689 26265 9723 26299
rect 11437 26265 11471 26299
rect 12173 26265 12207 26299
rect 17417 26265 17451 26299
rect 19625 26265 19659 26299
rect 2973 26197 3007 26231
rect 13645 26197 13679 26231
rect 16037 26197 16071 26231
rect 28549 26197 28583 26231
rect 2513 25993 2547 26027
rect 13277 25993 13311 26027
rect 21373 25993 21407 26027
rect 17785 25925 17819 25959
rect 19349 25925 19383 25959
rect 28917 25925 28951 25959
rect 2053 25857 2087 25891
rect 3341 25857 3375 25891
rect 13185 25857 13219 25891
rect 16957 25857 16991 25891
rect 20821 25857 20855 25891
rect 21281 25857 21315 25891
rect 23305 25857 23339 25891
rect 26617 25857 26651 25891
rect 27169 25857 27203 25891
rect 28825 25857 28859 25891
rect 29469 25857 29503 25891
rect 1869 25789 1903 25823
rect 3985 25789 4019 25823
rect 4261 25789 4295 25823
rect 17693 25789 17727 25823
rect 18521 25789 18555 25823
rect 19257 25789 19291 25823
rect 19533 25789 19567 25823
rect 27353 25789 27387 25823
rect 26433 25721 26467 25755
rect 3433 25653 3467 25687
rect 5733 25653 5767 25687
rect 17049 25653 17083 25687
rect 20637 25653 20671 25687
rect 23121 25653 23155 25687
rect 27629 25653 27663 25687
rect 29561 25653 29595 25687
rect 3341 25449 3375 25483
rect 19993 25449 20027 25483
rect 22385 25449 22419 25483
rect 27077 25449 27111 25483
rect 32965 25449 32999 25483
rect 38117 25449 38151 25483
rect 2053 25381 2087 25415
rect 4629 25381 4663 25415
rect 16405 25381 16439 25415
rect 4077 25313 4111 25347
rect 9137 25313 9171 25347
rect 18429 25313 18463 25347
rect 23397 25313 23431 25347
rect 28549 25313 28583 25347
rect 1961 25245 1995 25279
rect 2605 25245 2639 25279
rect 3249 25245 3283 25279
rect 8401 25245 8435 25279
rect 16313 25245 16347 25279
rect 20177 25245 20211 25279
rect 20913 25245 20947 25279
rect 22569 25245 22603 25279
rect 23581 25245 23615 25279
rect 24593 25245 24627 25279
rect 27261 25245 27295 25279
rect 27905 25245 27939 25279
rect 28733 25245 28767 25279
rect 32321 25245 32355 25279
rect 32413 25245 32447 25279
rect 33149 25245 33183 25279
rect 38301 25245 38335 25279
rect 4169 25177 4203 25211
rect 9413 25177 9447 25211
rect 2697 25109 2731 25143
rect 8493 25109 8527 25143
rect 10885 25109 10919 25143
rect 20729 25109 20763 25143
rect 24041 25109 24075 25143
rect 24685 25109 24719 25143
rect 27721 25109 27755 25143
rect 29193 25109 29227 25143
rect 19717 24905 19751 24939
rect 23949 24905 23983 24939
rect 17233 24837 17267 24871
rect 25329 24837 25363 24871
rect 30297 24837 30331 24871
rect 10885 24769 10919 24803
rect 16129 24769 16163 24803
rect 19901 24769 19935 24803
rect 21005 24769 21039 24803
rect 22661 24769 22695 24803
rect 23489 24769 23523 24803
rect 25881 24769 25915 24803
rect 28549 24769 28583 24803
rect 29009 24769 29043 24803
rect 29101 24769 29135 24803
rect 1777 24701 1811 24735
rect 2053 24701 2087 24735
rect 10977 24701 11011 24735
rect 13461 24701 13495 24735
rect 13737 24701 13771 24735
rect 16221 24701 16255 24735
rect 17141 24701 17175 24735
rect 17417 24701 17451 24735
rect 23305 24701 23339 24735
rect 25237 24701 25271 24735
rect 30205 24701 30239 24735
rect 30481 24701 30515 24735
rect 22753 24633 22787 24667
rect 3525 24565 3559 24599
rect 15209 24565 15243 24599
rect 20821 24565 20855 24599
rect 28365 24565 28399 24599
rect 1777 24361 1811 24395
rect 4077 24361 4111 24395
rect 15853 24361 15887 24395
rect 29009 24361 29043 24395
rect 6653 24293 6687 24327
rect 27629 24293 27663 24327
rect 20821 24225 20855 24259
rect 1593 24157 1627 24191
rect 3985 24157 4019 24191
rect 4905 24157 4939 24191
rect 9137 24157 9171 24191
rect 14565 24157 14599 24191
rect 15761 24157 15795 24191
rect 16405 24157 16439 24191
rect 18705 24157 18739 24191
rect 20637 24157 20671 24191
rect 23121 24157 23155 24191
rect 25421 24157 25455 24191
rect 27813 24157 27847 24191
rect 28457 24157 28491 24191
rect 28917 24157 28951 24191
rect 5181 24089 5215 24123
rect 16497 24089 16531 24123
rect 22017 24089 22051 24123
rect 22109 24089 22143 24123
rect 22661 24089 22695 24123
rect 9229 24021 9263 24055
rect 14657 24021 14691 24055
rect 18521 24021 18555 24055
rect 21281 24021 21315 24055
rect 23213 24021 23247 24055
rect 25237 24021 25271 24055
rect 28273 24021 28307 24055
rect 15025 23817 15059 23851
rect 21373 23817 21407 23851
rect 22109 23817 22143 23851
rect 28365 23817 28399 23851
rect 2237 23749 2271 23783
rect 6745 23749 6779 23783
rect 7297 23749 7331 23783
rect 25789 23749 25823 23783
rect 27353 23749 27387 23783
rect 27905 23749 27939 23783
rect 29929 23749 29963 23783
rect 30481 23749 30515 23783
rect 7757 23681 7791 23715
rect 16865 23681 16899 23715
rect 18061 23681 18095 23715
rect 19901 23681 19935 23715
rect 20361 23681 20395 23715
rect 20729 23681 20763 23715
rect 22017 23681 22051 23715
rect 25145 23681 25179 23715
rect 26341 23681 26375 23715
rect 28549 23681 28583 23715
rect 38301 23681 38335 23715
rect 1961 23613 1995 23647
rect 6653 23613 6687 23647
rect 13277 23613 13311 23647
rect 13553 23613 13587 23647
rect 18613 23613 18647 23647
rect 18797 23613 18831 23647
rect 20913 23613 20947 23647
rect 23305 23613 23339 23647
rect 25697 23613 25731 23647
rect 27261 23613 27295 23647
rect 29837 23613 29871 23647
rect 3709 23477 3743 23511
rect 7849 23477 7883 23511
rect 16957 23477 16991 23511
rect 17877 23477 17911 23511
rect 18981 23477 19015 23511
rect 19717 23477 19751 23511
rect 24961 23477 24995 23511
rect 38117 23477 38151 23511
rect 5733 23273 5767 23307
rect 18245 23273 18279 23307
rect 26617 23273 26651 23307
rect 27997 23273 28031 23307
rect 11161 23205 11195 23239
rect 19809 23205 19843 23239
rect 20545 23205 20579 23239
rect 22845 23205 22879 23239
rect 23673 23205 23707 23239
rect 4261 23137 4295 23171
rect 11529 23137 11563 23171
rect 13553 23137 13587 23171
rect 16405 23137 16439 23171
rect 16773 23137 16807 23171
rect 20361 23137 20395 23171
rect 22201 23137 22235 23171
rect 23305 23137 23339 23171
rect 23489 23137 23523 23171
rect 27353 23137 27387 23171
rect 28457 23137 28491 23171
rect 1593 23069 1627 23103
rect 3985 23069 4019 23103
rect 14749 23069 14783 23103
rect 15393 23069 15427 23103
rect 17509 23069 17543 23103
rect 18153 23069 18187 23103
rect 19533 23069 19567 23103
rect 20177 23069 20211 23103
rect 22385 23069 22419 23103
rect 25605 23069 25639 23103
rect 26801 23069 26835 23103
rect 27537 23069 27571 23103
rect 11805 23001 11839 23035
rect 16497 23001 16531 23035
rect 1777 22933 1811 22967
rect 14841 22933 14875 22967
rect 15485 22933 15519 22967
rect 17601 22933 17635 22967
rect 19349 22933 19383 22967
rect 25421 22933 25455 22967
rect 16221 22729 16255 22763
rect 19625 22729 19659 22763
rect 21373 22729 21407 22763
rect 25881 22729 25915 22763
rect 2053 22661 2087 22695
rect 15485 22661 15519 22695
rect 17509 22661 17543 22695
rect 18061 22661 18095 22695
rect 24777 22661 24811 22695
rect 24869 22661 24903 22695
rect 27353 22661 27387 22695
rect 2605 22593 2639 22627
rect 7573 22593 7607 22627
rect 8217 22593 8251 22627
rect 8861 22593 8895 22627
rect 10885 22593 10919 22627
rect 15393 22593 15427 22627
rect 16129 22593 16163 22627
rect 18705 22593 18739 22627
rect 19809 22593 19843 22627
rect 21281 22593 21315 22627
rect 26065 22593 26099 22627
rect 1961 22525 1995 22559
rect 9137 22525 9171 22559
rect 17417 22525 17451 22559
rect 18521 22525 18555 22559
rect 27261 22525 27295 22559
rect 27721 22525 27755 22559
rect 28365 22525 28399 22559
rect 8309 22457 8343 22491
rect 25329 22457 25363 22491
rect 7665 22389 7699 22423
rect 18889 22389 18923 22423
rect 1856 22185 1890 22219
rect 20085 22185 20119 22219
rect 26065 22185 26099 22219
rect 27261 22185 27295 22219
rect 24593 22117 24627 22151
rect 28917 22117 28951 22151
rect 1593 22049 1627 22083
rect 6837 22049 6871 22083
rect 8585 22049 8619 22083
rect 14289 22049 14323 22083
rect 14565 22049 14599 22083
rect 18153 22049 18187 22083
rect 21189 22049 21223 22083
rect 24041 22049 24075 22083
rect 28365 22049 28399 22083
rect 6561 21981 6595 22015
rect 9597 21981 9631 22015
rect 10517 21981 10551 22015
rect 13553 21981 13587 22015
rect 17325 21981 17359 22015
rect 17969 21981 18003 22015
rect 19441 21981 19475 22015
rect 19625 21981 19659 22015
rect 20545 21981 20579 22015
rect 20729 21981 20763 22015
rect 22293 21981 22327 22015
rect 24777 21981 24811 22015
rect 26249 21981 26283 22015
rect 27169 21981 27203 22015
rect 30113 21981 30147 22015
rect 38025 21981 38059 22015
rect 10793 21913 10827 21947
rect 12541 21913 12575 21947
rect 16313 21913 16347 21947
rect 23397 21913 23431 21947
rect 23489 21913 23523 21947
rect 28457 21913 28491 21947
rect 3341 21845 3375 21879
rect 9689 21845 9723 21879
rect 13645 21845 13679 21879
rect 17417 21845 17451 21879
rect 18613 21845 18647 21879
rect 22385 21845 22419 21879
rect 30205 21845 30239 21879
rect 38209 21845 38243 21879
rect 14565 21641 14599 21675
rect 16957 21641 16991 21675
rect 20177 21641 20211 21675
rect 24225 21641 24259 21675
rect 29561 21641 29595 21675
rect 22201 21573 22235 21607
rect 22293 21573 22327 21607
rect 1777 21505 1811 21539
rect 13829 21505 13863 21539
rect 14473 21505 14507 21539
rect 16865 21505 16899 21539
rect 20085 21505 20119 21539
rect 24409 21505 24443 21539
rect 28273 21505 28307 21539
rect 28365 21505 28399 21539
rect 29101 21505 29135 21539
rect 31217 21505 31251 21539
rect 6561 21437 6595 21471
rect 6837 21437 6871 21471
rect 8309 21437 8343 21471
rect 18245 21437 18279 21471
rect 18429 21437 18463 21471
rect 22477 21437 22511 21471
rect 28917 21437 28951 21471
rect 31309 21437 31343 21471
rect 8677 21369 8711 21403
rect 1593 21301 1627 21335
rect 13921 21301 13955 21335
rect 18889 21301 18923 21335
rect 4248 21097 4282 21131
rect 12081 21097 12115 21131
rect 22845 21097 22879 21131
rect 29745 21097 29779 21131
rect 30941 21097 30975 21131
rect 16773 21029 16807 21063
rect 28549 21029 28583 21063
rect 2789 20961 2823 20995
rect 3985 20961 4019 20995
rect 10609 20961 10643 20995
rect 17877 20961 17911 20995
rect 21281 20961 21315 20995
rect 27905 20961 27939 20995
rect 10333 20893 10367 20927
rect 14841 20893 14875 20927
rect 15669 20893 15703 20927
rect 16129 20893 16163 20927
rect 16957 20893 16991 20927
rect 19809 20893 19843 20927
rect 21465 20893 21499 20927
rect 23029 20893 23063 20927
rect 23489 20893 23523 20927
rect 27445 20893 27479 20927
rect 28089 20893 28123 20927
rect 29929 20893 29963 20927
rect 31125 20893 31159 20927
rect 2881 20825 2915 20859
rect 3433 20825 3467 20859
rect 16221 20825 16255 20859
rect 17969 20825 18003 20859
rect 18889 20825 18923 20859
rect 5733 20757 5767 20791
rect 14933 20757 14967 20791
rect 15485 20757 15519 20791
rect 19625 20757 19659 20791
rect 21925 20757 21959 20791
rect 23581 20757 23615 20791
rect 27261 20757 27295 20791
rect 1777 20553 1811 20587
rect 14657 20553 14691 20587
rect 20453 20553 20487 20587
rect 22017 20553 22051 20587
rect 27721 20553 27755 20587
rect 29285 20553 29319 20587
rect 31125 20553 31159 20587
rect 7573 20485 7607 20519
rect 16221 20485 16255 20519
rect 17049 20485 17083 20519
rect 19349 20485 19383 20519
rect 1961 20417 1995 20451
rect 7297 20417 7331 20451
rect 15485 20417 15519 20451
rect 16129 20417 16163 20451
rect 18061 20417 18095 20451
rect 20361 20417 20395 20451
rect 22201 20417 22235 20451
rect 23305 20417 23339 20451
rect 27905 20417 27939 20451
rect 29469 20417 29503 20451
rect 29929 20417 29963 20451
rect 31033 20417 31067 20451
rect 32965 20417 32999 20451
rect 9321 20349 9355 20383
rect 12909 20349 12943 20383
rect 13185 20349 13219 20383
rect 16957 20349 16991 20383
rect 17233 20349 17267 20383
rect 19257 20349 19291 20383
rect 19901 20349 19935 20383
rect 23121 20349 23155 20383
rect 30113 20349 30147 20383
rect 15577 20213 15611 20247
rect 18153 20213 18187 20247
rect 23489 20213 23523 20247
rect 30481 20213 30515 20247
rect 32781 20213 32815 20247
rect 1593 20009 1627 20043
rect 11253 20009 11287 20043
rect 15209 20009 15243 20043
rect 17785 20009 17819 20043
rect 21925 20009 21959 20043
rect 23213 20009 23247 20043
rect 30389 20009 30423 20043
rect 38117 20009 38151 20043
rect 25697 19941 25731 19975
rect 9505 19873 9539 19907
rect 9781 19873 9815 19907
rect 24593 19873 24627 19907
rect 28273 19873 28307 19907
rect 28917 19873 28951 19907
rect 1777 19805 1811 19839
rect 4445 19805 4479 19839
rect 7665 19805 7699 19839
rect 15117 19805 15151 19839
rect 17693 19805 17727 19839
rect 22109 19805 22143 19839
rect 22753 19805 22787 19839
rect 23397 19805 23431 19839
rect 24777 19805 24811 19839
rect 25881 19805 25915 19839
rect 26525 19805 26559 19839
rect 30297 19805 30331 19839
rect 38301 19805 38335 19839
rect 4721 19737 4755 19771
rect 6469 19737 6503 19771
rect 28365 19737 28399 19771
rect 7757 19669 7791 19703
rect 11713 19669 11747 19703
rect 22569 19669 22603 19703
rect 25237 19669 25271 19703
rect 26341 19669 26375 19703
rect 3985 19465 4019 19499
rect 21281 19465 21315 19499
rect 25329 19465 25363 19499
rect 11805 19397 11839 19431
rect 11897 19397 11931 19431
rect 15209 19397 15243 19431
rect 19349 19397 19383 19431
rect 27353 19397 27387 19431
rect 22569 19329 22603 19363
rect 25237 19329 25271 19363
rect 28365 19329 28399 19363
rect 29009 19329 29043 19363
rect 2237 19261 2271 19295
rect 2513 19261 2547 19295
rect 12265 19261 12299 19295
rect 13185 19261 13219 19295
rect 13461 19261 13495 19295
rect 16865 19261 16899 19295
rect 19257 19261 19291 19295
rect 19533 19261 19567 19295
rect 20637 19261 20671 19295
rect 20821 19261 20855 19295
rect 27261 19261 27295 19295
rect 28549 19261 28583 19295
rect 22385 19193 22419 19227
rect 27813 19193 27847 19227
rect 8309 18921 8343 18955
rect 19717 18921 19751 18955
rect 26801 18921 26835 18955
rect 27813 18921 27847 18955
rect 28457 18921 28491 18955
rect 30389 18921 30423 18955
rect 6101 18853 6135 18887
rect 15025 18853 15059 18887
rect 15669 18853 15703 18887
rect 26065 18853 26099 18887
rect 4353 18785 4387 18819
rect 6561 18785 6595 18819
rect 16405 18785 16439 18819
rect 20637 18785 20671 18819
rect 33517 18785 33551 18819
rect 2421 18717 2455 18751
rect 10333 18717 10367 18751
rect 15209 18717 15243 18751
rect 15853 18717 15887 18751
rect 19625 18717 19659 18751
rect 25605 18717 25639 18751
rect 26249 18717 26283 18751
rect 26709 18717 26743 18751
rect 27721 18717 27755 18751
rect 28365 18717 28399 18751
rect 29745 18717 29779 18751
rect 29929 18717 29963 18751
rect 33425 18717 33459 18751
rect 38301 18717 38335 18751
rect 4629 18649 4663 18683
rect 6837 18649 6871 18683
rect 10609 18649 10643 18683
rect 12357 18649 12391 18683
rect 16497 18649 16531 18683
rect 17049 18649 17083 18683
rect 17601 18649 17635 18683
rect 17693 18649 17727 18683
rect 18245 18649 18279 18683
rect 2513 18581 2547 18615
rect 22661 18581 22695 18615
rect 25421 18581 25455 18615
rect 38117 18581 38151 18615
rect 29653 18377 29687 18411
rect 24317 18309 24351 18343
rect 25513 18309 25547 18343
rect 1777 18241 1811 18275
rect 16313 18241 16347 18275
rect 17417 18241 17451 18275
rect 19809 18241 19843 18275
rect 20913 18241 20947 18275
rect 22477 18241 22511 18275
rect 30481 18241 30515 18275
rect 2329 18173 2363 18207
rect 2605 18173 2639 18207
rect 12909 18173 12943 18207
rect 13185 18173 13219 18207
rect 19993 18173 20027 18207
rect 21005 18173 21039 18207
rect 22661 18173 22695 18207
rect 24225 18173 24259 18207
rect 25421 18173 25455 18207
rect 25697 18173 25731 18207
rect 30941 18173 30975 18207
rect 14657 18105 14691 18139
rect 16129 18105 16163 18139
rect 24777 18105 24811 18139
rect 1593 18037 1627 18071
rect 4077 18037 4111 18071
rect 17233 18037 17267 18071
rect 20453 18037 20487 18071
rect 22845 18037 22879 18071
rect 30297 18037 30331 18071
rect 4616 17833 4650 17867
rect 14933 17833 14967 17867
rect 17693 17833 17727 17867
rect 22109 17833 22143 17867
rect 25145 17833 25179 17867
rect 29745 17833 29779 17867
rect 20913 17765 20947 17799
rect 26801 17765 26835 17799
rect 28089 17765 28123 17799
rect 4353 17697 4387 17731
rect 17233 17697 17267 17731
rect 18245 17697 18279 17731
rect 20361 17697 20395 17731
rect 22661 17697 22695 17731
rect 22845 17697 22879 17731
rect 27721 17697 27755 17731
rect 30389 17697 30423 17731
rect 9137 17629 9171 17663
rect 14841 17629 14875 17663
rect 15761 17629 15795 17663
rect 16405 17629 16439 17663
rect 17049 17629 17083 17663
rect 22017 17629 22051 17663
rect 25053 17629 25087 17663
rect 26157 17629 26191 17663
rect 26341 17629 26375 17663
rect 27905 17629 27939 17663
rect 29193 17629 29227 17663
rect 29929 17629 29963 17663
rect 30573 17629 30607 17663
rect 6377 17561 6411 17595
rect 9413 17561 9447 17595
rect 16497 17561 16531 17595
rect 18337 17561 18371 17595
rect 18889 17561 18923 17595
rect 20453 17561 20487 17595
rect 10885 17493 10919 17527
rect 15853 17493 15887 17527
rect 23305 17493 23339 17527
rect 29009 17493 29043 17527
rect 31033 17493 31067 17527
rect 9137 17289 9171 17323
rect 18245 17289 18279 17323
rect 21189 17289 21223 17323
rect 27261 17289 27295 17323
rect 29837 17289 29871 17323
rect 32965 17289 32999 17323
rect 7665 17221 7699 17255
rect 13553 17221 13587 17255
rect 18981 17221 19015 17255
rect 25973 17221 26007 17255
rect 26065 17221 26099 17255
rect 16129 17153 16163 17187
rect 16221 17153 16255 17187
rect 17049 17153 17083 17187
rect 18153 17153 18187 17187
rect 19993 17153 20027 17187
rect 20637 17153 20671 17187
rect 21097 17153 21131 17187
rect 22569 17153 22603 17187
rect 27169 17153 27203 17187
rect 30021 17153 30055 17187
rect 30481 17153 30515 17187
rect 30573 17153 30607 17187
rect 32505 17153 32539 17187
rect 38301 17153 38335 17187
rect 7389 17085 7423 17119
rect 13277 17085 13311 17119
rect 16865 17085 16899 17119
rect 18889 17085 18923 17119
rect 20177 17085 20211 17119
rect 22753 17085 22787 17119
rect 32321 17085 32355 17119
rect 19441 17017 19475 17051
rect 26525 17017 26559 17051
rect 15025 16949 15059 16983
rect 17509 16949 17543 16983
rect 22937 16949 22971 16983
rect 38117 16949 38151 16983
rect 6180 16745 6214 16779
rect 18429 16745 18463 16779
rect 21005 16745 21039 16779
rect 32413 16745 32447 16779
rect 16589 16677 16623 16711
rect 5917 16609 5951 16643
rect 10609 16609 10643 16643
rect 16037 16609 16071 16643
rect 30481 16609 30515 16643
rect 1777 16541 1811 16575
rect 10333 16541 10367 16575
rect 12817 16541 12851 16575
rect 15301 16541 15335 16575
rect 18337 16541 18371 16575
rect 21189 16541 21223 16575
rect 25145 16541 25179 16575
rect 26065 16541 26099 16575
rect 26525 16541 26559 16575
rect 27353 16541 27387 16575
rect 30665 16541 30699 16575
rect 32413 16541 32447 16575
rect 33517 16541 33551 16575
rect 12909 16473 12943 16507
rect 16129 16473 16163 16507
rect 1593 16405 1627 16439
rect 7665 16405 7699 16439
rect 12081 16405 12115 16439
rect 15393 16405 15427 16439
rect 24961 16405 24995 16439
rect 25881 16405 25915 16439
rect 26617 16405 26651 16439
rect 27169 16405 27203 16439
rect 31125 16405 31159 16439
rect 33609 16405 33643 16439
rect 19993 16201 20027 16235
rect 21005 16201 21039 16235
rect 23213 16201 23247 16235
rect 24409 16201 24443 16235
rect 25513 16201 25547 16235
rect 1869 16133 1903 16167
rect 13185 16133 13219 16167
rect 17509 16133 17543 16167
rect 18705 16133 18739 16167
rect 1593 16065 1627 16099
rect 8953 16065 8987 16099
rect 19257 16065 19291 16099
rect 20177 16065 20211 16099
rect 21189 16065 21223 16099
rect 25697 16065 25731 16099
rect 3617 15997 3651 16031
rect 9229 15997 9263 16031
rect 12909 15997 12943 16031
rect 14657 15997 14691 16031
rect 17417 15997 17451 16031
rect 18613 15997 18647 16031
rect 22569 15997 22603 16031
rect 22753 15997 22787 16031
rect 23765 15997 23799 16031
rect 23949 15997 23983 16031
rect 24869 15997 24903 16031
rect 28457 15997 28491 16031
rect 28641 15997 28675 16031
rect 29561 15997 29595 16031
rect 29745 15997 29779 16031
rect 17969 15929 18003 15963
rect 29101 15929 29135 15963
rect 29929 15929 29963 15963
rect 10701 15861 10735 15895
rect 14381 15657 14415 15691
rect 16405 15657 16439 15691
rect 17233 15657 17267 15691
rect 22753 15657 22787 15691
rect 23949 15657 23983 15691
rect 25237 15657 25271 15691
rect 27813 15657 27847 15691
rect 29837 15657 29871 15691
rect 30389 15657 30423 15691
rect 4077 15589 4111 15623
rect 15761 15589 15795 15623
rect 17877 15589 17911 15623
rect 21557 15589 21591 15623
rect 27077 15589 27111 15623
rect 32321 15589 32355 15623
rect 10977 15521 11011 15555
rect 18705 15521 18739 15555
rect 19809 15521 19843 15555
rect 20913 15521 20947 15555
rect 24593 15521 24627 15555
rect 26433 15521 26467 15555
rect 28457 15521 28491 15555
rect 3985 15453 4019 15487
rect 14289 15453 14323 15487
rect 15945 15453 15979 15487
rect 16589 15453 16623 15487
rect 17417 15453 17451 15487
rect 18061 15453 18095 15487
rect 21097 15453 21131 15487
rect 22661 15453 22695 15487
rect 23857 15453 23891 15487
rect 24777 15453 24811 15487
rect 26617 15453 26651 15487
rect 27997 15453 28031 15487
rect 29745 15453 29779 15487
rect 30573 15453 30607 15487
rect 31033 15453 31067 15487
rect 31677 15453 31711 15487
rect 32505 15453 32539 15487
rect 38025 15453 38059 15487
rect 11253 15385 11287 15419
rect 13001 15385 13035 15419
rect 19901 15385 19935 15419
rect 20453 15385 20487 15419
rect 31125 15385 31159 15419
rect 31769 15317 31803 15351
rect 38209 15317 38243 15351
rect 4445 15113 4479 15147
rect 17601 15113 17635 15147
rect 19901 15113 19935 15147
rect 21005 15113 21039 15147
rect 25421 15113 25455 15147
rect 25881 15113 25915 15147
rect 27261 15113 27295 15147
rect 28365 15113 28399 15147
rect 29009 15113 29043 15147
rect 5089 15045 5123 15079
rect 1869 14977 1903 15011
rect 3893 14977 3927 15011
rect 4353 14977 4387 15011
rect 4997 14977 5031 15011
rect 20085 14977 20119 15011
rect 20913 14977 20947 15011
rect 22201 14977 22235 15011
rect 26065 14977 26099 15011
rect 27169 14977 27203 15011
rect 28549 14977 28583 15011
rect 29193 14977 29227 15011
rect 2145 14909 2179 14943
rect 7481 14909 7515 14943
rect 7757 14909 7791 14943
rect 9505 14909 9539 14943
rect 13737 14909 13771 14943
rect 14013 14909 14047 14943
rect 15761 14909 15795 14943
rect 16957 14909 16991 14943
rect 17141 14909 17175 14943
rect 24777 14909 24811 14943
rect 24961 14909 24995 14943
rect 22017 14773 22051 14807
rect 3341 14569 3375 14603
rect 6653 14569 6687 14603
rect 11161 14569 11195 14603
rect 15485 14569 15519 14603
rect 21373 14569 21407 14603
rect 26341 14569 26375 14603
rect 28641 14569 28675 14603
rect 4169 14501 4203 14535
rect 11713 14501 11747 14535
rect 22017 14501 22051 14535
rect 25605 14501 25639 14535
rect 4905 14433 4939 14467
rect 9413 14433 9447 14467
rect 14841 14433 14875 14467
rect 16589 14433 16623 14467
rect 17233 14433 17267 14467
rect 19809 14433 19843 14467
rect 27997 14433 28031 14467
rect 3249 14365 3283 14399
rect 4077 14365 4111 14399
rect 11621 14365 11655 14399
rect 14749 14365 14783 14399
rect 15393 14365 15427 14399
rect 16313 14365 16347 14399
rect 18245 14365 18279 14399
rect 20453 14365 20487 14399
rect 21557 14365 21591 14399
rect 22201 14365 22235 14399
rect 22845 14365 22879 14399
rect 25789 14365 25823 14399
rect 26249 14365 26283 14399
rect 27537 14365 27571 14399
rect 28181 14365 28215 14399
rect 5181 14297 5215 14331
rect 9689 14297 9723 14331
rect 19901 14297 19935 14331
rect 18061 14229 18095 14263
rect 18705 14229 18739 14263
rect 22661 14229 22695 14263
rect 27353 14229 27387 14263
rect 22845 14025 22879 14059
rect 24501 14025 24535 14059
rect 26065 14025 26099 14059
rect 28273 14025 28307 14059
rect 38117 14025 38151 14059
rect 17233 13957 17267 13991
rect 18889 13957 18923 13991
rect 18981 13957 19015 13991
rect 23489 13957 23523 13991
rect 24041 13957 24075 13991
rect 2605 13889 2639 13923
rect 15853 13889 15887 13923
rect 24685 13889 24719 13923
rect 26249 13889 26283 13923
rect 27353 13889 27387 13923
rect 28457 13889 28491 13923
rect 38301 13889 38335 13923
rect 4353 13821 4387 13855
rect 16129 13821 16163 13855
rect 17141 13821 17175 13855
rect 17601 13821 17635 13855
rect 19349 13821 19383 13855
rect 19993 13821 20027 13855
rect 22201 13821 22235 13855
rect 22385 13821 22419 13855
rect 23397 13821 23431 13855
rect 2868 13685 2902 13719
rect 27169 13685 27203 13719
rect 11529 13481 11563 13515
rect 13001 13481 13035 13515
rect 15853 13481 15887 13515
rect 17969 13481 18003 13515
rect 24777 13481 24811 13515
rect 29929 13481 29963 13515
rect 30849 13413 30883 13447
rect 9781 13345 9815 13379
rect 10057 13345 10091 13379
rect 19441 13345 19475 13379
rect 23397 13345 23431 13379
rect 26893 13345 26927 13379
rect 30481 13345 30515 13379
rect 1593 13277 1627 13311
rect 12909 13277 12943 13311
rect 15025 13277 15059 13311
rect 15761 13277 15795 13311
rect 18153 13277 18187 13311
rect 19625 13277 19659 13311
rect 21741 13277 21775 13311
rect 24961 13277 24995 13311
rect 26709 13277 26743 13311
rect 28365 13277 28399 13311
rect 29009 13277 29043 13311
rect 29837 13277 29871 13311
rect 30665 13277 30699 13311
rect 1777 13141 1811 13175
rect 15117 13141 15151 13175
rect 20085 13141 20119 13175
rect 21557 13141 21591 13175
rect 27353 13141 27387 13175
rect 28181 13141 28215 13175
rect 28825 13141 28859 13175
rect 18705 12937 18739 12971
rect 26433 12937 26467 12971
rect 29101 12937 29135 12971
rect 2789 12869 2823 12903
rect 13369 12869 13403 12903
rect 16037 12869 16071 12903
rect 17417 12869 17451 12903
rect 20913 12869 20947 12903
rect 22109 12869 22143 12903
rect 22201 12869 22235 12903
rect 23305 12869 23339 12903
rect 2513 12801 2547 12835
rect 9229 12801 9263 12835
rect 15761 12801 15795 12835
rect 18889 12801 18923 12835
rect 23213 12801 23247 12835
rect 24409 12801 24443 12835
rect 25237 12801 25271 12835
rect 25881 12801 25915 12835
rect 26341 12801 26375 12835
rect 27169 12801 27203 12835
rect 27813 12801 27847 12835
rect 27905 12801 27939 12835
rect 28641 12801 28675 12835
rect 4261 12733 4295 12767
rect 6929 12733 6963 12767
rect 7205 12733 7239 12767
rect 13093 12733 13127 12767
rect 15117 12733 15151 12767
rect 17325 12733 17359 12767
rect 17601 12733 17635 12767
rect 20821 12733 20855 12767
rect 21189 12733 21223 12767
rect 22385 12733 22419 12767
rect 28457 12733 28491 12767
rect 25053 12665 25087 12699
rect 25697 12665 25731 12699
rect 8677 12597 8711 12631
rect 9321 12597 9355 12631
rect 24501 12597 24535 12631
rect 27261 12597 27295 12631
rect 3249 12393 3283 12427
rect 16589 12393 16623 12427
rect 18245 12393 18279 12427
rect 20821 12393 20855 12427
rect 22017 12393 22051 12427
rect 6377 12257 6411 12291
rect 12725 12257 12759 12291
rect 17325 12257 17359 12291
rect 20361 12257 20395 12291
rect 21465 12257 21499 12291
rect 3157 12189 3191 12223
rect 6101 12189 6135 12223
rect 11713 12189 11747 12223
rect 12633 12189 12667 12223
rect 13553 12189 13587 12223
rect 14289 12189 14323 12223
rect 16497 12189 16531 12223
rect 18429 12189 18463 12223
rect 20177 12189 20211 12223
rect 21373 12189 21407 12223
rect 22201 12189 22235 12223
rect 23489 12189 23523 12223
rect 25881 12189 25915 12223
rect 32137 12189 32171 12223
rect 14565 12121 14599 12155
rect 7849 12053 7883 12087
rect 11529 12053 11563 12087
rect 13645 12053 13679 12087
rect 16037 12053 16071 12087
rect 22661 12053 22695 12087
rect 23305 12053 23339 12087
rect 25697 12053 25731 12087
rect 32229 12053 32263 12087
rect 5733 11849 5767 11883
rect 14749 11849 14783 11883
rect 16221 11849 16255 11883
rect 27813 11849 27847 11883
rect 38117 11849 38151 11883
rect 8401 11781 8435 11815
rect 15393 11781 15427 11815
rect 17785 11781 17819 11815
rect 17877 11781 17911 11815
rect 18981 11781 19015 11815
rect 19073 11781 19107 11815
rect 25605 11781 25639 11815
rect 3985 11713 4019 11747
rect 8125 11713 8159 11747
rect 13553 11713 13587 11747
rect 14657 11713 14691 11747
rect 15301 11713 15335 11747
rect 16129 11713 16163 11747
rect 19625 11713 19659 11747
rect 23213 11713 23247 11747
rect 27353 11713 27387 11747
rect 32505 11713 32539 11747
rect 38301 11713 38335 11747
rect 4261 11645 4295 11679
rect 13277 11645 13311 11679
rect 13921 11645 13955 11679
rect 17049 11645 17083 11679
rect 18061 11645 18095 11679
rect 23397 11645 23431 11679
rect 25513 11645 25547 11679
rect 25789 11645 25823 11679
rect 27169 11645 27203 11679
rect 23581 11577 23615 11611
rect 9873 11509 9907 11543
rect 11805 11509 11839 11543
rect 32321 11509 32355 11543
rect 15761 11305 15795 11339
rect 18613 11305 18647 11339
rect 23397 11305 23431 11339
rect 25237 11305 25271 11339
rect 25973 11305 26007 11339
rect 27813 11305 27847 11339
rect 6745 11237 6779 11271
rect 15117 11237 15151 11271
rect 1869 11169 1903 11203
rect 4997 11169 5031 11203
rect 10517 11169 10551 11203
rect 16589 11169 16623 11203
rect 17509 11169 17543 11203
rect 20545 11169 20579 11203
rect 25053 11169 25087 11203
rect 1593 11101 1627 11135
rect 10241 11101 10275 11135
rect 15025 11101 15059 11135
rect 15669 11101 15703 11135
rect 16313 11101 16347 11135
rect 18797 11101 18831 11135
rect 19625 11101 19659 11135
rect 21649 11101 21683 11135
rect 22753 11101 22787 11135
rect 23581 11101 23615 11135
rect 24869 11101 24903 11135
rect 26157 11101 26191 11135
rect 27721 11101 27755 11135
rect 31309 11101 31343 11135
rect 5273 11033 5307 11067
rect 17601 11033 17635 11067
rect 18153 11033 18187 11067
rect 20637 11033 20671 11067
rect 21189 11033 21223 11067
rect 21741 11033 21775 11067
rect 11989 10965 12023 10999
rect 19441 10965 19475 10999
rect 22845 10965 22879 10999
rect 31401 10965 31435 10999
rect 8769 10761 8803 10795
rect 16129 10761 16163 10795
rect 18337 10761 18371 10795
rect 38117 10761 38151 10795
rect 16865 10693 16899 10727
rect 19349 10693 19383 10727
rect 19901 10693 19935 10727
rect 1593 10625 1627 10659
rect 7021 10625 7055 10659
rect 13829 10625 13863 10659
rect 16313 10625 16347 10659
rect 18245 10625 18279 10659
rect 23121 10625 23155 10659
rect 24225 10625 24259 10659
rect 24685 10625 24719 10659
rect 25513 10625 25547 10659
rect 27169 10625 27203 10659
rect 30849 10625 30883 10659
rect 38301 10625 38335 10659
rect 7297 10557 7331 10591
rect 14105 10557 14139 10591
rect 17601 10557 17635 10591
rect 19257 10557 19291 10591
rect 22937 10557 22971 10591
rect 27261 10489 27295 10523
rect 1777 10421 1811 10455
rect 15577 10421 15611 10455
rect 23581 10421 23615 10455
rect 24041 10421 24075 10455
rect 24777 10421 24811 10455
rect 25329 10421 25363 10455
rect 30941 10421 30975 10455
rect 4077 10217 4111 10251
rect 17785 10217 17819 10251
rect 18613 10217 18647 10251
rect 23121 10217 23155 10251
rect 3341 10149 3375 10183
rect 1593 10081 1627 10115
rect 7481 10081 7515 10115
rect 17141 10081 17175 10115
rect 20085 10081 20119 10115
rect 24869 10081 24903 10115
rect 26525 10081 26559 10115
rect 3985 10013 4019 10047
rect 5457 10013 5491 10047
rect 9873 10013 9907 10047
rect 17969 10013 18003 10047
rect 18797 10013 18831 10047
rect 20269 10013 20303 10047
rect 21741 10013 21775 10047
rect 21925 10013 21959 10047
rect 23305 10013 23339 10047
rect 24685 10013 24719 10047
rect 31401 10013 31435 10047
rect 33149 10013 33183 10047
rect 1869 9945 1903 9979
rect 5733 9945 5767 9979
rect 10149 9945 10183 9979
rect 16405 9945 16439 9979
rect 25881 9945 25915 9979
rect 25973 9945 26007 9979
rect 11621 9877 11655 9911
rect 20729 9877 20763 9911
rect 22385 9877 22419 9911
rect 25329 9877 25363 9911
rect 31217 9877 31251 9911
rect 32965 9877 32999 9911
rect 24685 9673 24719 9707
rect 27169 9673 27203 9707
rect 11161 9605 11195 9639
rect 17325 9605 17359 9639
rect 19717 9605 19751 9639
rect 29101 9605 29135 9639
rect 1593 9537 1627 9571
rect 3893 9537 3927 9571
rect 6837 9537 6871 9571
rect 11713 9537 11747 9571
rect 14197 9537 14231 9571
rect 18337 9537 18371 9571
rect 19625 9537 19659 9571
rect 22017 9537 22051 9571
rect 24041 9537 24075 9571
rect 25329 9537 25363 9571
rect 27353 9537 27387 9571
rect 27997 9537 28031 9571
rect 29009 9537 29043 9571
rect 1869 9469 1903 9503
rect 4169 9469 4203 9503
rect 7113 9469 7147 9503
rect 9137 9469 9171 9503
rect 9413 9469 9447 9503
rect 11989 9469 12023 9503
rect 13737 9469 13771 9503
rect 14473 9469 14507 9503
rect 17233 9469 17267 9503
rect 17509 9469 17543 9503
rect 18981 9469 19015 9503
rect 20637 9469 20671 9503
rect 20821 9469 20855 9503
rect 22753 9469 22787 9503
rect 24225 9469 24259 9503
rect 18429 9401 18463 9435
rect 25145 9401 25179 9435
rect 27813 9401 27847 9435
rect 3341 9333 3375 9367
rect 5641 9333 5675 9367
rect 8585 9333 8619 9367
rect 15945 9333 15979 9367
rect 21005 9333 21039 9367
rect 22109 9333 22143 9367
rect 4537 9129 4571 9163
rect 5457 9129 5491 9163
rect 6745 9129 6779 9163
rect 17141 9129 17175 9163
rect 26249 9129 26283 9163
rect 15301 9061 15335 9095
rect 18429 9061 18463 9095
rect 22569 9061 22603 9095
rect 7849 8993 7883 9027
rect 15945 8993 15979 9027
rect 17877 8993 17911 9027
rect 19625 8993 19659 9027
rect 19809 8993 19843 9027
rect 23213 8993 23247 9027
rect 23489 8993 23523 9027
rect 4721 8925 4755 8959
rect 5365 8925 5399 8959
rect 6009 8925 6043 8959
rect 6653 8925 6687 8959
rect 7757 8925 7791 8959
rect 15209 8925 15243 8959
rect 15853 8925 15887 8959
rect 16497 8925 16531 8959
rect 17325 8925 17359 8959
rect 20729 8925 20763 8959
rect 20821 8925 20855 8959
rect 25421 8925 25455 8959
rect 26157 8925 26191 8959
rect 27537 8925 27571 8959
rect 38025 8925 38059 8959
rect 6101 8857 6135 8891
rect 16589 8857 16623 8891
rect 17946 8857 17980 8891
rect 22017 8857 22051 8891
rect 22109 8857 22143 8891
rect 23305 8857 23339 8891
rect 20269 8789 20303 8823
rect 25237 8789 25271 8823
rect 27629 8789 27663 8823
rect 38209 8789 38243 8823
rect 6561 8585 6595 8619
rect 16957 8585 16991 8619
rect 19441 8585 19475 8619
rect 23581 8585 23615 8619
rect 8401 8517 8435 8551
rect 18153 8517 18187 8551
rect 1593 8449 1627 8483
rect 5825 8449 5859 8483
rect 5917 8449 5951 8483
rect 6745 8449 6779 8483
rect 8309 8449 8343 8483
rect 13277 8449 13311 8483
rect 15485 8449 15519 8483
rect 16129 8449 16163 8483
rect 16865 8449 16899 8483
rect 18797 8449 18831 8483
rect 19625 8449 19659 8483
rect 23029 8449 23063 8483
rect 23765 8449 23799 8483
rect 26433 8449 26467 8483
rect 13553 8381 13587 8415
rect 15025 8381 15059 8415
rect 17509 8381 17543 8415
rect 17693 8381 17727 8415
rect 25145 8381 25179 8415
rect 25329 8381 25363 8415
rect 1777 8313 1811 8347
rect 15577 8313 15611 8347
rect 16221 8313 16255 8347
rect 18613 8313 18647 8347
rect 22845 8313 22879 8347
rect 25513 8313 25547 8347
rect 26249 8313 26283 8347
rect 5365 8041 5399 8075
rect 9689 8041 9723 8075
rect 13185 8041 13219 8075
rect 17509 8041 17543 8075
rect 23949 8041 23983 8075
rect 26709 8041 26743 8075
rect 25145 7905 25179 7939
rect 5273 7837 5307 7871
rect 9597 7837 9631 7871
rect 10241 7837 10275 7871
rect 10885 7837 10919 7871
rect 12541 7837 12575 7871
rect 13093 7837 13127 7871
rect 16957 7837 16991 7871
rect 17693 7837 17727 7871
rect 18337 7837 18371 7871
rect 23857 7837 23891 7871
rect 26617 7837 26651 7871
rect 28733 7837 28767 7871
rect 14473 7769 14507 7803
rect 14565 7769 14599 7803
rect 15117 7769 15151 7803
rect 15577 7769 15611 7803
rect 16313 7769 16347 7803
rect 16405 7769 16439 7803
rect 10333 7701 10367 7735
rect 10977 7701 11011 7735
rect 12357 7701 12391 7735
rect 18153 7701 18187 7735
rect 28825 7701 28859 7735
rect 13001 7497 13035 7531
rect 14473 7497 14507 7531
rect 16957 7497 16991 7531
rect 22017 7497 22051 7531
rect 11897 7429 11931 7463
rect 19257 7429 19291 7463
rect 4813 7361 4847 7395
rect 6009 7361 6043 7395
rect 12909 7361 12943 7395
rect 15485 7361 15519 7395
rect 15945 7361 15979 7395
rect 16865 7361 16899 7395
rect 17509 7361 17543 7395
rect 22201 7361 22235 7395
rect 22845 7361 22879 7395
rect 23397 7361 23431 7395
rect 23489 7361 23523 7395
rect 24225 7361 24259 7395
rect 38025 7361 38059 7395
rect 9229 7293 9263 7327
rect 11805 7293 11839 7327
rect 12265 7293 12299 7327
rect 19165 7293 19199 7327
rect 24041 7293 24075 7327
rect 15301 7225 15335 7259
rect 19717 7225 19751 7259
rect 22661 7225 22695 7259
rect 4905 7157 4939 7191
rect 5825 7157 5859 7191
rect 16037 7157 16071 7191
rect 17601 7157 17635 7191
rect 24409 7157 24443 7191
rect 38209 7157 38243 7191
rect 6009 6953 6043 6987
rect 15485 6953 15519 6987
rect 9229 6817 9263 6851
rect 9873 6817 9907 6851
rect 19533 6817 19567 6851
rect 25145 6817 25179 6851
rect 2881 6749 2915 6783
rect 4721 6749 4755 6783
rect 6009 6749 6043 6783
rect 6745 6749 6779 6783
rect 7389 6749 7423 6783
rect 11713 6749 11747 6783
rect 11897 6749 11931 6783
rect 15669 6749 15703 6783
rect 16313 6749 16347 6783
rect 22201 6749 22235 6783
rect 22661 6749 22695 6783
rect 22845 6749 22879 6783
rect 23949 6749 23983 6783
rect 25053 6749 25087 6783
rect 9321 6681 9355 6715
rect 17785 6681 17819 6715
rect 17877 6681 17911 6715
rect 18429 6681 18463 6715
rect 19625 6681 19659 6715
rect 20177 6681 20211 6715
rect 2697 6613 2731 6647
rect 4813 6613 4847 6647
rect 6561 6613 6595 6647
rect 7205 6613 7239 6647
rect 12357 6613 12391 6647
rect 16129 6613 16163 6647
rect 22017 6613 22051 6647
rect 23305 6613 23339 6647
rect 23765 6613 23799 6647
rect 6745 6409 6779 6443
rect 14013 6409 14047 6443
rect 16865 6409 16899 6443
rect 19717 6409 19751 6443
rect 20361 6409 20395 6443
rect 23397 6409 23431 6443
rect 25789 6409 25823 6443
rect 8585 6341 8619 6375
rect 9965 6341 9999 6375
rect 15025 6341 15059 6375
rect 15761 6341 15795 6375
rect 1593 6273 1627 6307
rect 2329 6273 2363 6307
rect 4997 6273 5031 6307
rect 5641 6273 5675 6307
rect 6745 6273 6779 6307
rect 7573 6273 7607 6307
rect 9689 6273 9723 6307
rect 12265 6273 12299 6307
rect 13001 6273 13035 6307
rect 13921 6273 13955 6307
rect 14933 6273 14967 6307
rect 17049 6273 17083 6307
rect 17601 6273 17635 6307
rect 18613 6273 18647 6307
rect 19901 6273 19935 6307
rect 20545 6273 20579 6307
rect 23581 6273 23615 6307
rect 25697 6273 25731 6307
rect 8493 6205 8527 6239
rect 9137 6205 9171 6239
rect 15669 6205 15703 6239
rect 17693 6205 17727 6239
rect 1777 6137 1811 6171
rect 5457 6137 5491 6171
rect 16221 6137 16255 6171
rect 2421 6069 2455 6103
rect 4813 6069 4847 6103
rect 7389 6069 7423 6103
rect 12081 6069 12115 6103
rect 13093 6069 13127 6103
rect 18705 6069 18739 6103
rect 6377 5865 6411 5899
rect 7849 5865 7883 5899
rect 12265 5865 12299 5899
rect 14657 5865 14691 5899
rect 21373 5865 21407 5899
rect 29837 5865 29871 5899
rect 12909 5797 12943 5831
rect 13553 5797 13587 5831
rect 4905 5729 4939 5763
rect 14289 5729 14323 5763
rect 14473 5729 14507 5763
rect 37749 5729 37783 5763
rect 4353 5661 4387 5695
rect 4813 5661 4847 5695
rect 6285 5661 6319 5695
rect 7113 5661 7147 5695
rect 7757 5661 7791 5695
rect 12449 5661 12483 5695
rect 13093 5661 13127 5695
rect 13737 5661 13771 5695
rect 15853 5661 15887 5695
rect 16497 5661 16531 5695
rect 18889 5661 18923 5695
rect 21281 5661 21315 5695
rect 29745 5661 29779 5695
rect 37473 5661 37507 5695
rect 7205 5593 7239 5627
rect 16589 5593 16623 5627
rect 4169 5525 4203 5559
rect 15945 5525 15979 5559
rect 18705 5525 18739 5559
rect 7389 5253 7423 5287
rect 10425 5253 10459 5287
rect 1593 5185 1627 5219
rect 6561 5185 6595 5219
rect 10149 5185 10183 5219
rect 11713 5185 11747 5219
rect 14013 5185 14047 5219
rect 15301 5185 15335 5219
rect 31677 5185 31711 5219
rect 32505 5185 32539 5219
rect 7297 5117 7331 5151
rect 7941 5117 7975 5151
rect 15393 5117 15427 5151
rect 31493 5049 31527 5083
rect 1777 4981 1811 5015
rect 6653 4981 6687 5015
rect 11805 4981 11839 5015
rect 13829 4981 13863 5015
rect 32321 4981 32355 5015
rect 12081 4573 12115 4607
rect 17693 4573 17727 4607
rect 27721 4573 27755 4607
rect 11161 4437 11195 4471
rect 11897 4437 11931 4471
rect 17785 4437 17819 4471
rect 27813 4437 27847 4471
rect 12357 4233 12391 4267
rect 11713 4097 11747 4131
rect 11897 4097 11931 4131
rect 17049 4097 17083 4131
rect 16865 3961 16899 3995
rect 1593 3689 1627 3723
rect 1777 3485 1811 3519
rect 6653 3485 6687 3519
rect 11161 3485 11195 3519
rect 18613 3485 18647 3519
rect 38025 3485 38059 3519
rect 6469 3349 6503 3383
rect 11253 3349 11287 3383
rect 18429 3349 18463 3383
rect 38209 3349 38243 3383
rect 6653 3145 6687 3179
rect 13369 3145 13403 3179
rect 16865 3145 16899 3179
rect 17601 3145 17635 3179
rect 36737 3145 36771 3179
rect 18337 3077 18371 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 6561 3009 6595 3043
rect 9689 3009 9723 3043
rect 11069 3009 11103 3043
rect 13277 3009 13311 3043
rect 17049 3009 17083 3043
rect 17509 3009 17543 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 18245 2941 18279 2975
rect 2329 2873 2363 2907
rect 10885 2873 10919 2907
rect 18797 2873 18831 2907
rect 1777 2805 1811 2839
rect 9505 2805 9539 2839
rect 38209 2805 38243 2839
rect 2697 2601 2731 2635
rect 10425 2601 10459 2635
rect 15577 2601 15611 2635
rect 22017 2601 22051 2635
rect 24593 2601 24627 2635
rect 27169 2601 27203 2635
rect 27813 2601 27847 2635
rect 29745 2601 29779 2635
rect 32321 2601 32355 2635
rect 35541 2601 35575 2635
rect 36737 2601 36771 2635
rect 12357 2533 12391 2567
rect 31033 2533 31067 2567
rect 1593 2397 1627 2431
rect 2881 2397 2915 2431
rect 4629 2397 4663 2431
rect 6561 2397 6595 2431
rect 7849 2397 7883 2431
rect 9137 2397 9171 2431
rect 10609 2397 10643 2431
rect 12541 2397 12575 2431
rect 14289 2397 14323 2431
rect 15761 2397 15795 2431
rect 16865 2397 16899 2431
rect 18613 2397 18647 2431
rect 20085 2397 20119 2431
rect 22201 2397 22235 2431
rect 23305 2397 23339 2431
rect 24777 2397 24811 2431
rect 27353 2397 27387 2431
rect 27997 2397 28031 2431
rect 29929 2397 29963 2431
rect 31217 2397 31251 2431
rect 32505 2397 32539 2431
rect 35081 2397 35115 2431
rect 35725 2397 35759 2431
rect 36921 2397 36955 2431
rect 37473 2397 37507 2431
rect 1777 2261 1811 2295
rect 4813 2261 4847 2295
rect 6745 2261 6779 2295
rect 8033 2261 8067 2295
rect 9321 2261 9355 2295
rect 14473 2261 14507 2295
rect 17049 2261 17083 2295
rect 18797 2261 18831 2295
rect 20269 2261 20303 2295
rect 23489 2261 23523 2295
rect 34897 2261 34931 2295
rect 37657 2261 37691 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 36081 37451 36139 37457
rect 36081 37417 36093 37451
rect 36127 37448 36139 37451
rect 39298 37448 39304 37460
rect 36127 37420 39304 37448
rect 36127 37417 36139 37420
rect 36081 37411 36139 37417
rect 39298 37408 39304 37420
rect 39356 37408 39362 37460
rect 37458 37312 37464 37324
rect 37419 37284 37464 37312
rect 37458 37272 37464 37284
rect 37516 37272 37522 37324
rect 1578 37244 1584 37256
rect 1539 37216 1584 37244
rect 1578 37204 1584 37216
rect 1636 37204 1642 37256
rect 1946 37204 1952 37256
rect 2004 37244 2010 37256
rect 2501 37247 2559 37253
rect 2501 37244 2513 37247
rect 2004 37216 2513 37244
rect 2004 37204 2010 37216
rect 2501 37213 2513 37216
rect 2547 37213 2559 37247
rect 3142 37244 3148 37256
rect 3103 37216 3148 37244
rect 2501 37207 2559 37213
rect 3142 37204 3148 37216
rect 3200 37204 3206 37256
rect 4154 37244 4160 37256
rect 4115 37216 4160 37244
rect 4154 37204 4160 37216
rect 4212 37204 4218 37256
rect 5166 37204 5172 37256
rect 5224 37244 5230 37256
rect 5445 37247 5503 37253
rect 5445 37244 5457 37247
rect 5224 37216 5457 37244
rect 5224 37204 5230 37216
rect 5445 37213 5457 37216
rect 5491 37213 5503 37247
rect 5445 37207 5503 37213
rect 7098 37204 7104 37256
rect 7156 37244 7162 37256
rect 7377 37247 7435 37253
rect 7377 37244 7389 37247
rect 7156 37216 7389 37244
rect 7156 37204 7162 37216
rect 7377 37213 7389 37216
rect 7423 37213 7435 37247
rect 7377 37207 7435 37213
rect 8386 37204 8392 37256
rect 8444 37244 8450 37256
rect 9309 37247 9367 37253
rect 9309 37244 9321 37247
rect 8444 37216 9321 37244
rect 8444 37204 8450 37216
rect 9309 37213 9321 37216
rect 9355 37213 9367 37247
rect 9309 37207 9367 37213
rect 10318 37204 10324 37256
rect 10376 37244 10382 37256
rect 10597 37247 10655 37253
rect 10597 37244 10609 37247
rect 10376 37216 10609 37244
rect 10376 37204 10382 37216
rect 10597 37213 10609 37216
rect 10643 37213 10655 37247
rect 10597 37207 10655 37213
rect 11606 37204 11612 37256
rect 11664 37244 11670 37256
rect 11885 37247 11943 37253
rect 11885 37244 11897 37247
rect 11664 37216 11897 37244
rect 11664 37204 11670 37216
rect 11885 37213 11897 37216
rect 11931 37213 11943 37247
rect 11885 37207 11943 37213
rect 11974 37204 11980 37256
rect 12032 37244 12038 37256
rect 12989 37247 13047 37253
rect 12989 37244 13001 37247
rect 12032 37216 13001 37244
rect 12032 37204 12038 37216
rect 12989 37213 13001 37216
rect 13035 37213 13047 37247
rect 12989 37207 13047 37213
rect 14826 37204 14832 37256
rect 14884 37244 14890 37256
rect 15105 37247 15163 37253
rect 15105 37244 15117 37247
rect 14884 37216 15117 37244
rect 14884 37204 14890 37216
rect 15105 37213 15117 37216
rect 15151 37213 15163 37247
rect 15105 37207 15163 37213
rect 16114 37204 16120 37256
rect 16172 37244 16178 37256
rect 17037 37247 17095 37253
rect 17037 37244 17049 37247
rect 16172 37216 17049 37244
rect 16172 37204 16178 37216
rect 17037 37213 17049 37216
rect 17083 37213 17095 37247
rect 17037 37207 17095 37213
rect 17218 37204 17224 37256
rect 17276 37244 17282 37256
rect 18141 37247 18199 37253
rect 18141 37244 18153 37247
rect 17276 37216 18153 37244
rect 17276 37204 17282 37216
rect 18141 37213 18153 37216
rect 18187 37213 18199 37247
rect 18141 37207 18199 37213
rect 18966 37204 18972 37256
rect 19024 37244 19030 37256
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 19024 37216 19441 37244
rect 19024 37204 19030 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 19429 37207 19487 37213
rect 20717 37247 20775 37253
rect 20717 37213 20729 37247
rect 20763 37244 20775 37247
rect 20806 37244 20812 37256
rect 20763 37216 20812 37244
rect 20763 37213 20775 37216
rect 20717 37207 20775 37213
rect 20806 37204 20812 37216
rect 20864 37204 20870 37256
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 22612 37216 22845 37244
rect 22612 37204 22618 37216
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 22833 37207 22891 37213
rect 23290 37204 23296 37256
rect 23348 37244 23354 37256
rect 24581 37247 24639 37253
rect 24581 37244 24593 37247
rect 23348 37216 24593 37244
rect 23348 37204 23354 37216
rect 24581 37213 24593 37216
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 26053 37247 26111 37253
rect 26053 37244 26065 37247
rect 25832 37216 26065 37244
rect 25832 37204 25838 37216
rect 26053 37213 26065 37216
rect 26099 37213 26111 37247
rect 27154 37244 27160 37256
rect 27115 37216 27160 37244
rect 26053 37207 26111 37213
rect 27154 37204 27160 37216
rect 27212 37204 27218 37256
rect 28994 37204 29000 37256
rect 29052 37244 29058 37256
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29052 37216 29929 37244
rect 29052 37204 29058 37216
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 29917 37207 29975 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30561 37247 30619 37253
rect 30561 37244 30573 37247
rect 30432 37216 30573 37244
rect 30432 37204 30438 37216
rect 30561 37213 30573 37216
rect 30607 37213 30619 37247
rect 30561 37207 30619 37213
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 31812 37216 32505 37244
rect 31812 37204 31818 37216
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33560 37216 33793 37244
rect 33560 37204 33566 37216
rect 33781 37213 33793 37216
rect 33827 37213 33839 37247
rect 33781 37207 33839 37213
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34848 37216 35081 37244
rect 34848 37204 34854 37216
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 35434 37204 35440 37256
rect 35492 37244 35498 37256
rect 35897 37247 35955 37253
rect 35897 37244 35909 37247
rect 35492 37216 35909 37244
rect 35492 37204 35498 37216
rect 35897 37213 35909 37216
rect 35943 37213 35955 37247
rect 36630 37244 36636 37256
rect 36591 37216 36636 37244
rect 35897 37207 35955 37213
rect 36630 37204 36636 37216
rect 36688 37204 36694 37256
rect 37734 37244 37740 37256
rect 37695 37216 37740 37244
rect 37734 37204 37740 37216
rect 37792 37204 37798 37256
rect 2774 37176 2780 37188
rect 1780 37148 2780 37176
rect 1780 37117 1808 37148
rect 2774 37136 2780 37148
rect 2832 37136 2838 37188
rect 6822 37176 6828 37188
rect 3988 37148 6828 37176
rect 1765 37111 1823 37117
rect 1765 37077 1777 37111
rect 1811 37077 1823 37111
rect 2314 37108 2320 37120
rect 2275 37080 2320 37108
rect 1765 37071 1823 37077
rect 2314 37068 2320 37080
rect 2372 37068 2378 37120
rect 2961 37111 3019 37117
rect 2961 37077 2973 37111
rect 3007 37108 3019 37111
rect 3878 37108 3884 37120
rect 3007 37080 3884 37108
rect 3007 37077 3019 37080
rect 2961 37071 3019 37077
rect 3878 37068 3884 37080
rect 3936 37068 3942 37120
rect 3988 37117 4016 37148
rect 6822 37136 6828 37148
rect 6880 37136 6886 37188
rect 23750 37136 23756 37188
rect 23808 37176 23814 37188
rect 23808 37148 25912 37176
rect 23808 37136 23814 37148
rect 3973 37111 4031 37117
rect 3973 37077 3985 37111
rect 4019 37077 4031 37111
rect 3973 37071 4031 37077
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 5261 37111 5319 37117
rect 5261 37108 5273 37111
rect 4672 37080 5273 37108
rect 4672 37068 4678 37080
rect 5261 37077 5273 37080
rect 5307 37077 5319 37111
rect 7190 37108 7196 37120
rect 7151 37080 7196 37108
rect 5261 37071 5319 37077
rect 7190 37068 7196 37080
rect 7248 37068 7254 37120
rect 9122 37108 9128 37120
rect 9083 37080 9128 37108
rect 9122 37068 9128 37080
rect 9180 37068 9186 37120
rect 10410 37108 10416 37120
rect 10371 37080 10416 37108
rect 10410 37068 10416 37080
rect 10468 37068 10474 37120
rect 11698 37108 11704 37120
rect 11659 37080 11704 37108
rect 11698 37068 11704 37080
rect 11756 37068 11762 37120
rect 12894 37068 12900 37120
rect 12952 37108 12958 37120
rect 13173 37111 13231 37117
rect 13173 37108 13185 37111
rect 12952 37080 13185 37108
rect 12952 37068 12958 37080
rect 13173 37077 13185 37080
rect 13219 37077 13231 37111
rect 13173 37071 13231 37077
rect 14734 37068 14740 37120
rect 14792 37108 14798 37120
rect 14921 37111 14979 37117
rect 14921 37108 14933 37111
rect 14792 37080 14933 37108
rect 14792 37068 14798 37080
rect 14921 37077 14933 37080
rect 14967 37077 14979 37111
rect 14921 37071 14979 37077
rect 16574 37068 16580 37120
rect 16632 37108 16638 37120
rect 16853 37111 16911 37117
rect 16853 37108 16865 37111
rect 16632 37080 16865 37108
rect 16632 37068 16638 37080
rect 16853 37077 16865 37080
rect 16899 37077 16911 37111
rect 16853 37071 16911 37077
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18325 37111 18383 37117
rect 18325 37108 18337 37111
rect 18104 37080 18337 37108
rect 18104 37068 18110 37080
rect 18325 37077 18337 37080
rect 18371 37077 18383 37111
rect 18325 37071 18383 37077
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 19613 37111 19671 37117
rect 19613 37108 19625 37111
rect 19392 37080 19625 37108
rect 19392 37068 19398 37080
rect 19613 37077 19625 37080
rect 19659 37077 19671 37111
rect 19613 37071 19671 37077
rect 20714 37068 20720 37120
rect 20772 37108 20778 37120
rect 20901 37111 20959 37117
rect 20901 37108 20913 37111
rect 20772 37080 20913 37108
rect 20772 37068 20778 37080
rect 20901 37077 20913 37080
rect 20947 37077 20959 37111
rect 20901 37071 20959 37077
rect 20990 37068 20996 37120
rect 21048 37108 21054 37120
rect 22649 37111 22707 37117
rect 22649 37108 22661 37111
rect 21048 37080 22661 37108
rect 21048 37068 21054 37080
rect 22649 37077 22661 37080
rect 22695 37077 22707 37111
rect 22649 37071 22707 37077
rect 23842 37068 23848 37120
rect 23900 37108 23906 37120
rect 25884 37117 25912 37148
rect 27430 37136 27436 37188
rect 27488 37176 27494 37188
rect 27488 37148 32352 37176
rect 27488 37136 27494 37148
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 23900 37080 24777 37108
rect 23900 37068 23906 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25869 37111 25927 37117
rect 25869 37077 25881 37111
rect 25915 37077 25927 37111
rect 25869 37071 25927 37077
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27120 37080 27353 37108
rect 27120 37068 27126 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 29730 37108 29736 37120
rect 29691 37080 29736 37108
rect 27341 37071 27399 37077
rect 29730 37068 29736 37080
rect 29788 37068 29794 37120
rect 30374 37108 30380 37120
rect 30335 37080 30380 37108
rect 30374 37068 30380 37080
rect 30432 37068 30438 37120
rect 32324 37117 32352 37148
rect 32309 37111 32367 37117
rect 32309 37077 32321 37111
rect 32355 37077 32367 37111
rect 32309 37071 32367 37077
rect 32398 37068 32404 37120
rect 32456 37108 32462 37120
rect 33597 37111 33655 37117
rect 33597 37108 33609 37111
rect 32456 37080 33609 37108
rect 32456 37068 32462 37080
rect 33597 37077 33609 37080
rect 33643 37077 33655 37111
rect 33597 37071 33655 37077
rect 34606 37068 34612 37120
rect 34664 37108 34670 37120
rect 34885 37111 34943 37117
rect 34885 37108 34897 37111
rect 34664 37080 34897 37108
rect 34664 37068 34670 37080
rect 34885 37077 34897 37080
rect 34931 37077 34943 37111
rect 34885 37071 34943 37077
rect 36722 37068 36728 37120
rect 36780 37108 36786 37120
rect 36817 37111 36875 37117
rect 36817 37108 36829 37111
rect 36780 37080 36829 37108
rect 36780 37068 36786 37080
rect 36817 37077 36829 37080
rect 36863 37077 36875 37111
rect 36817 37071 36875 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 658 36864 664 36916
rect 716 36904 722 36916
rect 1765 36907 1823 36913
rect 1765 36904 1777 36907
rect 716 36876 1777 36904
rect 716 36864 722 36876
rect 1765 36873 1777 36876
rect 1811 36873 1823 36907
rect 1765 36867 1823 36873
rect 34149 36907 34207 36913
rect 34149 36873 34161 36907
rect 34195 36904 34207 36907
rect 34195 36876 35894 36904
rect 34195 36873 34207 36876
rect 34149 36867 34207 36873
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36768 1639 36771
rect 2866 36768 2872 36780
rect 1627 36740 2872 36768
rect 1627 36737 1639 36740
rect 1581 36731 1639 36737
rect 2866 36728 2872 36740
rect 2924 36728 2930 36780
rect 34330 36768 34336 36780
rect 34291 36740 34336 36768
rect 34330 36728 34336 36740
rect 34388 36728 34394 36780
rect 35866 36768 35894 36876
rect 38010 36864 38016 36916
rect 38068 36904 38074 36916
rect 38197 36907 38255 36913
rect 38197 36904 38209 36907
rect 38068 36876 38209 36904
rect 38068 36864 38074 36876
rect 38197 36873 38209 36876
rect 38243 36873 38255 36907
rect 38197 36867 38255 36873
rect 38013 36771 38071 36777
rect 38013 36768 38025 36771
rect 35866 36740 38025 36768
rect 38013 36737 38025 36740
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 30285 36363 30343 36369
rect 30285 36329 30297 36363
rect 30331 36360 30343 36363
rect 36630 36360 36636 36372
rect 30331 36332 36636 36360
rect 30331 36329 30343 36332
rect 30285 36323 30343 36329
rect 36630 36320 36636 36332
rect 36688 36320 36694 36372
rect 38194 36360 38200 36372
rect 38155 36332 38200 36360
rect 38194 36320 38200 36332
rect 38252 36320 38258 36372
rect 1762 36156 1768 36168
rect 1723 36128 1768 36156
rect 1762 36116 1768 36128
rect 1820 36116 1826 36168
rect 29822 36116 29828 36168
rect 29880 36156 29886 36168
rect 30469 36159 30527 36165
rect 30469 36156 30481 36159
rect 29880 36128 30481 36156
rect 29880 36116 29886 36128
rect 30469 36125 30481 36128
rect 30515 36125 30527 36159
rect 38010 36156 38016 36168
rect 37971 36128 38016 36156
rect 30469 36119 30527 36125
rect 38010 36116 38016 36128
rect 38068 36116 38074 36168
rect 1581 36023 1639 36029
rect 1581 35989 1593 36023
rect 1627 36020 1639 36023
rect 3510 36020 3516 36032
rect 1627 35992 3516 36020
rect 1627 35989 1639 35992
rect 1581 35983 1639 35989
rect 3510 35980 3516 35992
rect 3568 35980 3574 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 33413 35819 33471 35825
rect 33413 35785 33425 35819
rect 33459 35816 33471 35819
rect 34330 35816 34336 35828
rect 33459 35788 34336 35816
rect 33459 35785 33471 35788
rect 33413 35779 33471 35785
rect 34330 35776 34336 35788
rect 34388 35776 34394 35828
rect 33318 35680 33324 35692
rect 33279 35652 33324 35680
rect 33318 35640 33324 35652
rect 33376 35640 33382 35692
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 38286 35068 38292 35080
rect 38247 35040 38292 35068
rect 38286 35028 38292 35040
rect 38344 35028 38350 35080
rect 37274 34892 37280 34944
rect 37332 34932 37338 34944
rect 38105 34935 38163 34941
rect 38105 34932 38117 34935
rect 37332 34904 38117 34932
rect 37332 34892 37338 34904
rect 38105 34901 38117 34904
rect 38151 34901 38163 34935
rect 38105 34895 38163 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1578 34688 1584 34740
rect 1636 34728 1642 34740
rect 1765 34731 1823 34737
rect 1765 34728 1777 34731
rect 1636 34700 1777 34728
rect 1636 34688 1642 34700
rect 1765 34697 1777 34700
rect 1811 34697 1823 34731
rect 1765 34691 1823 34697
rect 37461 34731 37519 34737
rect 37461 34697 37473 34731
rect 37507 34728 37519 34731
rect 38010 34728 38016 34740
rect 37507 34700 38016 34728
rect 37507 34697 37519 34700
rect 37461 34691 37519 34697
rect 38010 34688 38016 34700
rect 38068 34688 38074 34740
rect 1946 34592 1952 34604
rect 1907 34564 1952 34592
rect 1946 34552 1952 34564
rect 2004 34552 2010 34604
rect 15286 34592 15292 34604
rect 15247 34564 15292 34592
rect 15286 34552 15292 34564
rect 15344 34552 15350 34604
rect 36446 34552 36452 34604
rect 36504 34592 36510 34604
rect 37645 34595 37703 34601
rect 37645 34592 37657 34595
rect 36504 34564 37657 34592
rect 36504 34552 36510 34564
rect 37645 34561 37657 34564
rect 37691 34561 37703 34595
rect 37645 34555 37703 34561
rect 15381 34527 15439 34533
rect 15381 34493 15393 34527
rect 15427 34524 15439 34527
rect 17402 34524 17408 34536
rect 15427 34496 17408 34524
rect 15427 34493 15439 34496
rect 15381 34487 15439 34493
rect 17402 34484 17408 34496
rect 17460 34484 17466 34536
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 34885 34187 34943 34193
rect 34885 34153 34897 34187
rect 34931 34184 34943 34187
rect 35434 34184 35440 34196
rect 34931 34156 35440 34184
rect 34931 34153 34943 34156
rect 34885 34147 34943 34153
rect 35434 34144 35440 34156
rect 35492 34144 35498 34196
rect 12158 34008 12164 34060
rect 12216 34048 12222 34060
rect 12216 34020 13492 34048
rect 12216 34008 12222 34020
rect 1762 33980 1768 33992
rect 1723 33952 1768 33980
rect 1762 33940 1768 33952
rect 1820 33940 1826 33992
rect 13464 33989 13492 34020
rect 12805 33983 12863 33989
rect 12805 33949 12817 33983
rect 12851 33980 12863 33983
rect 13449 33983 13507 33989
rect 12851 33952 13308 33980
rect 12851 33949 12863 33952
rect 12805 33943 12863 33949
rect 1581 33847 1639 33853
rect 1581 33813 1593 33847
rect 1627 33844 1639 33847
rect 1670 33844 1676 33856
rect 1627 33816 1676 33844
rect 1627 33813 1639 33816
rect 1581 33807 1639 33813
rect 1670 33804 1676 33816
rect 1728 33804 1734 33856
rect 12618 33844 12624 33856
rect 12579 33816 12624 33844
rect 12618 33804 12624 33816
rect 12676 33804 12682 33856
rect 13280 33853 13308 33952
rect 13449 33949 13461 33983
rect 13495 33949 13507 33983
rect 13449 33943 13507 33949
rect 34514 33940 34520 33992
rect 34572 33980 34578 33992
rect 35069 33983 35127 33989
rect 35069 33980 35081 33983
rect 34572 33952 35081 33980
rect 34572 33940 34578 33952
rect 35069 33949 35081 33952
rect 35115 33949 35127 33983
rect 35069 33943 35127 33949
rect 13265 33847 13323 33853
rect 13265 33813 13277 33847
rect 13311 33813 13323 33847
rect 13265 33807 13323 33813
rect 13538 33804 13544 33856
rect 13596 33844 13602 33856
rect 14277 33847 14335 33853
rect 14277 33844 14289 33847
rect 13596 33816 14289 33844
rect 13596 33804 13602 33816
rect 14277 33813 14289 33816
rect 14323 33813 14335 33847
rect 14277 33807 14335 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1946 33640 1952 33652
rect 1907 33612 1952 33640
rect 1946 33600 1952 33612
rect 2004 33600 2010 33652
rect 17218 33640 17224 33652
rect 17179 33612 17224 33640
rect 17218 33600 17224 33612
rect 17276 33600 17282 33652
rect 23290 33640 23296 33652
rect 23251 33612 23296 33640
rect 23290 33600 23296 33612
rect 23348 33600 23354 33652
rect 12618 33532 12624 33584
rect 12676 33572 12682 33584
rect 12676 33544 13768 33572
rect 12676 33532 12682 33544
rect 1857 33507 1915 33513
rect 1857 33473 1869 33507
rect 1903 33473 1915 33507
rect 1857 33467 1915 33473
rect 1872 33436 1900 33467
rect 2130 33464 2136 33516
rect 2188 33504 2194 33516
rect 2501 33507 2559 33513
rect 2501 33504 2513 33507
rect 2188 33476 2513 33504
rect 2188 33464 2194 33476
rect 2501 33473 2513 33476
rect 2547 33473 2559 33507
rect 2501 33467 2559 33473
rect 11701 33507 11759 33513
rect 11701 33473 11713 33507
rect 11747 33504 11759 33507
rect 12158 33504 12164 33516
rect 11747 33476 12164 33504
rect 11747 33473 11759 33476
rect 11701 33467 11759 33473
rect 12158 33464 12164 33476
rect 12216 33464 12222 33516
rect 13538 33504 13544 33516
rect 13499 33476 13544 33504
rect 13538 33464 13544 33476
rect 13596 33464 13602 33516
rect 13740 33513 13768 33544
rect 13725 33507 13783 33513
rect 13725 33473 13737 33507
rect 13771 33473 13783 33507
rect 17402 33504 17408 33516
rect 17363 33476 17408 33504
rect 13725 33467 13783 33473
rect 17402 33464 17408 33476
rect 17460 33464 17466 33516
rect 22830 33464 22836 33516
rect 22888 33504 22894 33516
rect 23477 33507 23535 33513
rect 23477 33504 23489 33507
rect 22888 33476 23489 33504
rect 22888 33464 22894 33476
rect 23477 33473 23489 33476
rect 23523 33473 23535 33507
rect 38286 33504 38292 33516
rect 38247 33476 38292 33504
rect 23477 33467 23535 33473
rect 38286 33464 38292 33476
rect 38344 33464 38350 33516
rect 3050 33436 3056 33448
rect 1872 33408 3056 33436
rect 3050 33396 3056 33408
rect 3108 33396 3114 33448
rect 2222 33260 2228 33312
rect 2280 33300 2286 33312
rect 2593 33303 2651 33309
rect 2593 33300 2605 33303
rect 2280 33272 2605 33300
rect 2280 33260 2286 33272
rect 2593 33269 2605 33272
rect 2639 33269 2651 33303
rect 11790 33300 11796 33312
rect 11751 33272 11796 33300
rect 2593 33263 2651 33269
rect 11790 33260 11796 33272
rect 11848 33260 11854 33312
rect 13906 33300 13912 33312
rect 13867 33272 13912 33300
rect 13906 33260 13912 33272
rect 13964 33300 13970 33312
rect 15286 33300 15292 33312
rect 13964 33272 15292 33300
rect 13964 33260 13970 33272
rect 15286 33260 15292 33272
rect 15344 33260 15350 33312
rect 29454 33260 29460 33312
rect 29512 33300 29518 33312
rect 38105 33303 38163 33309
rect 38105 33300 38117 33303
rect 29512 33272 38117 33300
rect 29512 33260 29518 33272
rect 38105 33269 38117 33272
rect 38151 33269 38163 33303
rect 38105 33263 38163 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 2866 33096 2872 33108
rect 2827 33068 2872 33096
rect 2866 33056 2872 33068
rect 2924 33056 2930 33108
rect 23109 33099 23167 33105
rect 23109 33065 23121 33099
rect 23155 33096 23167 33099
rect 27154 33096 27160 33108
rect 23155 33068 27160 33096
rect 23155 33065 23167 33068
rect 23109 33059 23167 33065
rect 27154 33056 27160 33068
rect 27212 33056 27218 33108
rect 14737 33031 14795 33037
rect 14737 32997 14749 33031
rect 14783 32997 14795 33031
rect 14737 32991 14795 32997
rect 4065 32963 4123 32969
rect 4065 32960 4077 32963
rect 3068 32932 4077 32960
rect 1762 32892 1768 32904
rect 1723 32864 1768 32892
rect 1762 32852 1768 32864
rect 1820 32852 1826 32904
rect 3068 32901 3096 32932
rect 4065 32929 4077 32932
rect 4111 32929 4123 32963
rect 14752 32960 14780 32991
rect 14752 32932 15608 32960
rect 4065 32923 4123 32929
rect 3053 32895 3111 32901
rect 3053 32861 3065 32895
rect 3099 32861 3111 32895
rect 3053 32855 3111 32861
rect 3973 32895 4031 32901
rect 3973 32861 3985 32895
rect 4019 32892 4031 32895
rect 6178 32892 6184 32904
rect 4019 32864 6184 32892
rect 4019 32861 4031 32864
rect 3973 32855 4031 32861
rect 6178 32852 6184 32864
rect 6236 32852 6242 32904
rect 9122 32892 9128 32904
rect 9083 32864 9128 32892
rect 9122 32852 9128 32864
rect 9180 32852 9186 32904
rect 13354 32852 13360 32904
rect 13412 32892 13418 32904
rect 15580 32901 15608 32932
rect 14921 32895 14979 32901
rect 14921 32892 14933 32895
rect 13412 32864 14933 32892
rect 13412 32852 13418 32864
rect 14921 32861 14933 32864
rect 14967 32861 14979 32895
rect 14921 32855 14979 32861
rect 15565 32895 15623 32901
rect 15565 32861 15577 32895
rect 15611 32861 15623 32895
rect 23290 32892 23296 32904
rect 23251 32864 23296 32892
rect 15565 32855 15623 32861
rect 23290 32852 23296 32864
rect 23348 32852 23354 32904
rect 1581 32759 1639 32765
rect 1581 32725 1593 32759
rect 1627 32756 1639 32759
rect 1854 32756 1860 32768
rect 1627 32728 1860 32756
rect 1627 32725 1639 32728
rect 1581 32719 1639 32725
rect 1854 32716 1860 32728
rect 1912 32716 1918 32768
rect 6546 32716 6552 32768
rect 6604 32756 6610 32768
rect 9217 32759 9275 32765
rect 9217 32756 9229 32759
rect 6604 32728 9229 32756
rect 6604 32716 6610 32728
rect 9217 32725 9229 32728
rect 9263 32756 9275 32759
rect 11238 32756 11244 32768
rect 9263 32728 11244 32756
rect 9263 32725 9275 32728
rect 9217 32719 9275 32725
rect 11238 32716 11244 32728
rect 11296 32716 11302 32768
rect 15378 32756 15384 32768
rect 15339 32728 15384 32756
rect 15378 32716 15384 32728
rect 15436 32716 15442 32768
rect 15654 32716 15660 32768
rect 15712 32756 15718 32768
rect 16025 32759 16083 32765
rect 16025 32756 16037 32759
rect 15712 32728 16037 32756
rect 15712 32716 15718 32728
rect 16025 32725 16037 32728
rect 16071 32725 16083 32759
rect 16025 32719 16083 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 12345 32555 12403 32561
rect 12345 32521 12357 32555
rect 12391 32552 12403 32555
rect 13906 32552 13912 32564
rect 12391 32524 13912 32552
rect 12391 32521 12403 32524
rect 12345 32515 12403 32521
rect 13906 32512 13912 32524
rect 13964 32512 13970 32564
rect 18966 32552 18972 32564
rect 18927 32524 18972 32552
rect 18966 32512 18972 32524
rect 19024 32512 19030 32564
rect 19705 32555 19763 32561
rect 19705 32521 19717 32555
rect 19751 32552 19763 32555
rect 23290 32552 23296 32564
rect 19751 32524 23296 32552
rect 19751 32521 19763 32524
rect 19705 32515 19763 32521
rect 23290 32512 23296 32524
rect 23348 32512 23354 32564
rect 7193 32487 7251 32493
rect 7193 32453 7205 32487
rect 7239 32484 7251 32487
rect 7239 32456 11744 32484
rect 7239 32453 7251 32456
rect 7193 32447 7251 32453
rect 1486 32376 1492 32428
rect 1544 32416 1550 32428
rect 1857 32419 1915 32425
rect 1857 32416 1869 32419
rect 1544 32388 1869 32416
rect 1544 32376 1550 32388
rect 1857 32385 1869 32388
rect 1903 32385 1915 32419
rect 4614 32416 4620 32428
rect 4575 32388 4620 32416
rect 1857 32379 1915 32385
rect 4614 32376 4620 32388
rect 4672 32376 4678 32428
rect 6546 32416 6552 32428
rect 6507 32388 6552 32416
rect 6546 32376 6552 32388
rect 6604 32376 6610 32428
rect 6822 32376 6828 32428
rect 6880 32416 6886 32428
rect 7653 32419 7711 32425
rect 7653 32416 7665 32419
rect 6880 32388 7665 32416
rect 6880 32376 6886 32388
rect 7653 32385 7665 32388
rect 7699 32385 7711 32419
rect 7653 32379 7711 32385
rect 4709 32351 4767 32357
rect 4709 32317 4721 32351
rect 4755 32348 4767 32351
rect 5261 32351 5319 32357
rect 5261 32348 5273 32351
rect 4755 32320 5273 32348
rect 4755 32317 4767 32320
rect 4709 32311 4767 32317
rect 5261 32317 5273 32320
rect 5307 32317 5319 32351
rect 5442 32348 5448 32360
rect 5403 32320 5448 32348
rect 5261 32311 5319 32317
rect 5442 32308 5448 32320
rect 5500 32308 5506 32360
rect 6730 32348 6736 32360
rect 6691 32320 6736 32348
rect 6730 32308 6736 32320
rect 6788 32308 6794 32360
rect 5905 32283 5963 32289
rect 5905 32249 5917 32283
rect 5951 32280 5963 32283
rect 7760 32280 7788 32456
rect 10321 32419 10379 32425
rect 10321 32385 10333 32419
rect 10367 32416 10379 32419
rect 11057 32419 11115 32425
rect 10367 32388 10916 32416
rect 10367 32385 10379 32388
rect 10321 32379 10379 32385
rect 10888 32289 10916 32388
rect 11057 32385 11069 32419
rect 11103 32416 11115 32419
rect 11146 32416 11152 32428
rect 11103 32388 11152 32416
rect 11103 32385 11115 32388
rect 11057 32379 11115 32385
rect 11146 32376 11152 32388
rect 11204 32376 11210 32428
rect 11716 32425 11744 32456
rect 15378 32444 15384 32496
rect 15436 32484 15442 32496
rect 15436 32456 15884 32484
rect 15436 32444 15442 32456
rect 11701 32419 11759 32425
rect 11701 32385 11713 32419
rect 11747 32385 11759 32419
rect 11701 32379 11759 32385
rect 11790 32376 11796 32428
rect 11848 32416 11854 32428
rect 11885 32419 11943 32425
rect 11885 32416 11897 32419
rect 11848 32388 11897 32416
rect 11848 32376 11854 32388
rect 11885 32385 11897 32388
rect 11931 32385 11943 32419
rect 11885 32379 11943 32385
rect 13357 32419 13415 32425
rect 13357 32385 13369 32419
rect 13403 32416 13415 32419
rect 13446 32416 13452 32428
rect 13403 32388 13452 32416
rect 13403 32385 13415 32388
rect 13357 32379 13415 32385
rect 13446 32376 13452 32388
rect 13504 32376 13510 32428
rect 14182 32416 14188 32428
rect 14143 32388 14188 32416
rect 14182 32376 14188 32388
rect 14240 32376 14246 32428
rect 14734 32416 14740 32428
rect 14695 32388 14740 32416
rect 14734 32376 14740 32388
rect 14792 32376 14798 32428
rect 15654 32416 15660 32428
rect 15615 32388 15660 32416
rect 15654 32376 15660 32388
rect 15712 32376 15718 32428
rect 15856 32425 15884 32456
rect 15841 32419 15899 32425
rect 15841 32385 15853 32419
rect 15887 32385 15899 32419
rect 15841 32379 15899 32385
rect 16390 32376 16396 32428
rect 16448 32416 16454 32428
rect 17037 32419 17095 32425
rect 17037 32416 17049 32419
rect 16448 32388 17049 32416
rect 16448 32376 16454 32388
rect 17037 32385 17049 32388
rect 17083 32385 17095 32419
rect 17037 32379 17095 32385
rect 19153 32419 19211 32425
rect 19153 32385 19165 32419
rect 19199 32416 19211 32419
rect 19426 32416 19432 32428
rect 19199 32388 19432 32416
rect 19199 32385 19211 32388
rect 19153 32379 19211 32385
rect 19426 32376 19432 32388
rect 19484 32376 19490 32428
rect 19613 32419 19671 32425
rect 19613 32385 19625 32419
rect 19659 32385 19671 32419
rect 19613 32379 19671 32385
rect 27617 32419 27675 32425
rect 27617 32385 27629 32419
rect 27663 32416 27675 32419
rect 34606 32416 34612 32428
rect 27663 32388 34612 32416
rect 27663 32385 27675 32388
rect 27617 32379 27675 32385
rect 19334 32308 19340 32360
rect 19392 32348 19398 32360
rect 19628 32348 19656 32379
rect 34606 32376 34612 32388
rect 34664 32376 34670 32428
rect 19392 32320 19656 32348
rect 19392 32308 19398 32320
rect 5951 32252 7788 32280
rect 10873 32283 10931 32289
rect 5951 32249 5963 32252
rect 5905 32243 5963 32249
rect 10873 32249 10885 32283
rect 10919 32249 10931 32283
rect 10873 32243 10931 32249
rect 1946 32212 1952 32224
rect 1907 32184 1952 32212
rect 1946 32172 1952 32184
rect 2004 32172 2010 32224
rect 7742 32212 7748 32224
rect 7703 32184 7748 32212
rect 7742 32172 7748 32184
rect 7800 32172 7806 32224
rect 10134 32212 10140 32224
rect 10095 32184 10140 32212
rect 10134 32172 10140 32184
rect 10192 32172 10198 32224
rect 11882 32172 11888 32224
rect 11940 32212 11946 32224
rect 13449 32215 13507 32221
rect 13449 32212 13461 32215
rect 11940 32184 13461 32212
rect 11940 32172 11946 32184
rect 13449 32181 13461 32184
rect 13495 32181 13507 32215
rect 13998 32212 14004 32224
rect 13959 32184 14004 32212
rect 13449 32175 13507 32181
rect 13998 32172 14004 32184
rect 14056 32172 14062 32224
rect 14090 32172 14096 32224
rect 14148 32212 14154 32224
rect 14829 32215 14887 32221
rect 14829 32212 14841 32215
rect 14148 32184 14841 32212
rect 14148 32172 14154 32184
rect 14829 32181 14841 32184
rect 14875 32181 14887 32215
rect 16022 32212 16028 32224
rect 15983 32184 16028 32212
rect 14829 32175 14887 32181
rect 16022 32172 16028 32184
rect 16080 32172 16086 32224
rect 16853 32215 16911 32221
rect 16853 32181 16865 32215
rect 16899 32212 16911 32215
rect 17402 32212 17408 32224
rect 16899 32184 17408 32212
rect 16899 32181 16911 32184
rect 16853 32175 16911 32181
rect 17402 32172 17408 32184
rect 17460 32172 17466 32224
rect 25038 32172 25044 32224
rect 25096 32212 25102 32224
rect 27709 32215 27767 32221
rect 27709 32212 27721 32215
rect 25096 32184 27721 32212
rect 25096 32172 25102 32184
rect 27709 32181 27721 32184
rect 27755 32181 27767 32215
rect 27709 32175 27767 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 5077 32011 5135 32017
rect 5077 31977 5089 32011
rect 5123 32008 5135 32011
rect 5442 32008 5448 32020
rect 5123 31980 5448 32008
rect 5123 31977 5135 31980
rect 5077 31971 5135 31977
rect 5442 31968 5448 31980
rect 5500 31968 5506 32020
rect 11517 32011 11575 32017
rect 11517 31977 11529 32011
rect 11563 32008 11575 32011
rect 11974 32008 11980 32020
rect 11563 31980 11980 32008
rect 11563 31977 11575 31980
rect 11517 31971 11575 31977
rect 11974 31968 11980 31980
rect 12032 31968 12038 32020
rect 13449 32011 13507 32017
rect 13449 31977 13461 32011
rect 13495 32008 13507 32011
rect 16022 32008 16028 32020
rect 13495 31980 16028 32008
rect 13495 31977 13507 31980
rect 13449 31971 13507 31977
rect 16022 31968 16028 31980
rect 16080 32008 16086 32020
rect 16942 32008 16948 32020
rect 16080 31980 16948 32008
rect 16080 31968 16086 31980
rect 16942 31968 16948 31980
rect 17000 31968 17006 32020
rect 2041 31943 2099 31949
rect 2041 31909 2053 31943
rect 2087 31909 2099 31943
rect 2041 31903 2099 31909
rect 2685 31943 2743 31949
rect 2685 31909 2697 31943
rect 2731 31940 2743 31943
rect 2866 31940 2872 31952
rect 2731 31912 2872 31940
rect 2731 31909 2743 31912
rect 2685 31903 2743 31909
rect 2056 31872 2084 31903
rect 2866 31900 2872 31912
rect 2924 31900 2930 31952
rect 7374 31900 7380 31952
rect 7432 31940 7438 31952
rect 7742 31940 7748 31952
rect 7432 31912 7748 31940
rect 7432 31900 7438 31912
rect 7742 31900 7748 31912
rect 7800 31940 7806 31952
rect 12161 31943 12219 31949
rect 7800 31912 9904 31940
rect 7800 31900 7806 31912
rect 2056 31844 2912 31872
rect 2225 31807 2283 31813
rect 2225 31773 2237 31807
rect 2271 31804 2283 31807
rect 2774 31804 2780 31816
rect 2271 31776 2780 31804
rect 2271 31773 2283 31776
rect 2225 31767 2283 31773
rect 2774 31764 2780 31776
rect 2832 31764 2838 31816
rect 2884 31813 2912 31844
rect 9214 31832 9220 31884
rect 9272 31872 9278 31884
rect 9769 31875 9827 31881
rect 9769 31872 9781 31875
rect 9272 31844 9781 31872
rect 9272 31832 9278 31844
rect 9769 31841 9781 31844
rect 9815 31841 9827 31875
rect 9876 31872 9904 31912
rect 12161 31909 12173 31943
rect 12207 31940 12219 31943
rect 13630 31940 13636 31952
rect 12207 31912 13636 31940
rect 12207 31909 12219 31912
rect 12161 31903 12219 31909
rect 13630 31900 13636 31912
rect 13688 31900 13694 31952
rect 14829 31943 14887 31949
rect 14829 31909 14841 31943
rect 14875 31940 14887 31943
rect 15746 31940 15752 31952
rect 14875 31912 15752 31940
rect 14875 31909 14887 31912
rect 14829 31903 14887 31909
rect 15746 31900 15752 31912
rect 15804 31900 15810 31952
rect 17586 31900 17592 31952
rect 17644 31940 17650 31952
rect 17644 31912 25912 31940
rect 17644 31900 17650 31912
rect 12805 31875 12863 31881
rect 12805 31872 12817 31875
rect 9876 31844 12817 31872
rect 9769 31835 9827 31841
rect 12805 31841 12817 31844
rect 12851 31841 12863 31875
rect 21358 31872 21364 31884
rect 21319 31844 21364 31872
rect 12805 31835 12863 31841
rect 21358 31832 21364 31844
rect 21416 31832 21422 31884
rect 2869 31807 2927 31813
rect 2869 31773 2881 31807
rect 2915 31773 2927 31807
rect 5258 31804 5264 31816
rect 5219 31776 5264 31804
rect 2869 31767 2927 31773
rect 5258 31764 5264 31776
rect 5316 31764 5322 31816
rect 9677 31807 9735 31813
rect 9677 31773 9689 31807
rect 9723 31804 9735 31807
rect 10410 31804 10416 31816
rect 9723 31776 10416 31804
rect 9723 31773 9735 31776
rect 9677 31767 9735 31773
rect 10410 31764 10416 31776
rect 10468 31764 10474 31816
rect 10870 31764 10876 31816
rect 10928 31804 10934 31816
rect 11701 31807 11759 31813
rect 11701 31804 11713 31807
rect 10928 31776 11713 31804
rect 10928 31764 10934 31776
rect 11701 31773 11713 31776
rect 11747 31773 11759 31807
rect 11701 31767 11759 31773
rect 12345 31807 12403 31813
rect 12345 31773 12357 31807
rect 12391 31773 12403 31807
rect 12986 31804 12992 31816
rect 12947 31776 12992 31804
rect 12345 31767 12403 31773
rect 10594 31696 10600 31748
rect 10652 31736 10658 31748
rect 12360 31736 12388 31767
rect 12986 31764 12992 31776
rect 13044 31764 13050 31816
rect 13998 31764 14004 31816
rect 14056 31804 14062 31816
rect 15013 31807 15071 31813
rect 15013 31804 15025 31807
rect 14056 31776 15025 31804
rect 14056 31764 14062 31776
rect 15013 31773 15025 31776
rect 15059 31773 15071 31807
rect 16390 31804 16396 31816
rect 16351 31776 16396 31804
rect 15013 31767 15071 31773
rect 16390 31764 16396 31776
rect 16448 31764 16454 31816
rect 16485 31807 16543 31813
rect 16485 31773 16497 31807
rect 16531 31804 16543 31807
rect 16758 31804 16764 31816
rect 16531 31776 16764 31804
rect 16531 31773 16543 31776
rect 16485 31767 16543 31773
rect 16758 31764 16764 31776
rect 16816 31764 16822 31816
rect 17402 31804 17408 31816
rect 17363 31776 17408 31804
rect 17402 31764 17408 31776
rect 17460 31764 17466 31816
rect 20714 31804 20720 31816
rect 20675 31776 20720 31804
rect 20714 31764 20720 31776
rect 20772 31764 20778 31816
rect 20901 31807 20959 31813
rect 20901 31773 20913 31807
rect 20947 31804 20959 31807
rect 22922 31804 22928 31816
rect 20947 31776 22928 31804
rect 20947 31773 20959 31776
rect 20901 31767 20959 31773
rect 22922 31764 22928 31776
rect 22980 31764 22986 31816
rect 25884 31813 25912 31912
rect 25961 31875 26019 31881
rect 25961 31841 25973 31875
rect 26007 31872 26019 31875
rect 29822 31872 29828 31884
rect 26007 31844 29828 31872
rect 26007 31841 26019 31844
rect 25961 31835 26019 31841
rect 29822 31832 29828 31844
rect 29880 31832 29886 31884
rect 37366 31832 37372 31884
rect 37424 31872 37430 31884
rect 38289 31875 38347 31881
rect 38289 31872 38301 31875
rect 37424 31844 38301 31872
rect 37424 31832 37430 31844
rect 38289 31841 38301 31844
rect 38335 31841 38347 31875
rect 38289 31835 38347 31841
rect 25869 31807 25927 31813
rect 25869 31773 25881 31807
rect 25915 31773 25927 31807
rect 38102 31804 38108 31816
rect 38063 31776 38108 31804
rect 25869 31767 25927 31773
rect 38102 31764 38108 31776
rect 38160 31764 38166 31816
rect 10652 31708 12388 31736
rect 10652 31696 10658 31708
rect 3694 31628 3700 31680
rect 3752 31668 3758 31680
rect 11146 31668 11152 31680
rect 3752 31640 11152 31668
rect 3752 31628 3758 31640
rect 11146 31628 11152 31640
rect 11204 31628 11210 31680
rect 17218 31668 17224 31680
rect 17179 31640 17224 31668
rect 17218 31628 17224 31640
rect 17276 31628 17282 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 4985 31467 5043 31473
rect 4985 31433 4997 31467
rect 5031 31464 5043 31467
rect 5258 31464 5264 31476
rect 5031 31436 5264 31464
rect 5031 31433 5043 31436
rect 4985 31427 5043 31433
rect 5258 31424 5264 31436
rect 5316 31424 5322 31476
rect 6641 31467 6699 31473
rect 6641 31433 6653 31467
rect 6687 31464 6699 31467
rect 6730 31464 6736 31476
rect 6687 31436 6736 31464
rect 6687 31433 6699 31436
rect 6641 31427 6699 31433
rect 6730 31424 6736 31436
rect 6788 31424 6794 31476
rect 13446 31464 13452 31476
rect 12406 31436 13452 31464
rect 9401 31399 9459 31405
rect 9401 31365 9413 31399
rect 9447 31396 9459 31399
rect 10134 31396 10140 31408
rect 9447 31368 10140 31396
rect 9447 31365 9459 31368
rect 9401 31359 9459 31365
rect 10134 31356 10140 31368
rect 10192 31356 10198 31408
rect 1946 31288 1952 31340
rect 2004 31328 2010 31340
rect 2133 31331 2191 31337
rect 2133 31328 2145 31331
rect 2004 31300 2145 31328
rect 2004 31288 2010 31300
rect 2133 31297 2145 31300
rect 2179 31297 2191 31331
rect 5166 31328 5172 31340
rect 5127 31300 5172 31328
rect 2133 31291 2191 31297
rect 5166 31288 5172 31300
rect 5224 31328 5230 31340
rect 6549 31331 6607 31337
rect 6549 31328 6561 31331
rect 5224 31300 6561 31328
rect 5224 31288 5230 31300
rect 6549 31297 6561 31300
rect 6595 31297 6607 31331
rect 6549 31291 6607 31297
rect 7190 31288 7196 31340
rect 7248 31328 7254 31340
rect 8573 31331 8631 31337
rect 8573 31328 8585 31331
rect 7248 31300 8585 31328
rect 7248 31288 7254 31300
rect 8573 31297 8585 31300
rect 8619 31297 8631 31331
rect 10686 31328 10692 31340
rect 10647 31300 10692 31328
rect 8573 31291 8631 31297
rect 10686 31288 10692 31300
rect 10744 31288 10750 31340
rect 12253 31331 12311 31337
rect 12253 31297 12265 31331
rect 12299 31328 12311 31331
rect 12406 31328 12434 31436
rect 13446 31424 13452 31436
rect 13504 31464 13510 31476
rect 16390 31464 16396 31476
rect 13504 31436 16396 31464
rect 13504 31424 13510 31436
rect 16390 31424 16396 31436
rect 16448 31424 16454 31476
rect 19426 31424 19432 31476
rect 19484 31464 19490 31476
rect 19889 31467 19947 31473
rect 19889 31464 19901 31467
rect 19484 31436 19901 31464
rect 19484 31424 19490 31436
rect 19889 31433 19901 31436
rect 19935 31433 19947 31467
rect 20714 31464 20720 31476
rect 20675 31436 20720 31464
rect 19889 31427 19947 31433
rect 20714 31424 20720 31436
rect 20772 31424 20778 31476
rect 22281 31467 22339 31473
rect 22281 31433 22293 31467
rect 22327 31433 22339 31467
rect 22922 31464 22928 31476
rect 22883 31436 22928 31464
rect 22281 31427 22339 31433
rect 16574 31396 16580 31408
rect 14108 31368 16580 31396
rect 13630 31328 13636 31340
rect 12299 31300 12434 31328
rect 13591 31300 13636 31328
rect 12299 31297 12311 31300
rect 12253 31291 12311 31297
rect 13630 31288 13636 31300
rect 13688 31288 13694 31340
rect 14108 31337 14136 31368
rect 16574 31356 16580 31368
rect 16632 31356 16638 31408
rect 16942 31396 16948 31408
rect 16903 31368 16948 31396
rect 16942 31356 16948 31368
rect 17000 31356 17006 31408
rect 17037 31399 17095 31405
rect 17037 31365 17049 31399
rect 17083 31396 17095 31399
rect 17218 31396 17224 31408
rect 17083 31368 17224 31396
rect 17083 31365 17095 31368
rect 17037 31359 17095 31365
rect 17218 31356 17224 31368
rect 17276 31356 17282 31408
rect 22296 31396 22324 31427
rect 22922 31424 22928 31436
rect 22980 31424 22986 31476
rect 22296 31368 23152 31396
rect 14093 31331 14151 31337
rect 14093 31297 14105 31331
rect 14139 31297 14151 31331
rect 14093 31291 14151 31297
rect 16025 31331 16083 31337
rect 16025 31297 16037 31331
rect 16071 31328 16083 31331
rect 16390 31328 16396 31340
rect 16071 31300 16396 31328
rect 16071 31297 16083 31300
rect 16025 31291 16083 31297
rect 16390 31288 16396 31300
rect 16448 31288 16454 31340
rect 19797 31331 19855 31337
rect 19797 31297 19809 31331
rect 19843 31328 19855 31331
rect 21358 31328 21364 31340
rect 19843 31300 21364 31328
rect 19843 31297 19855 31300
rect 19797 31291 19855 31297
rect 21358 31288 21364 31300
rect 21416 31288 21422 31340
rect 22462 31328 22468 31340
rect 22423 31300 22468 31328
rect 22462 31288 22468 31300
rect 22520 31288 22526 31340
rect 23124 31337 23152 31368
rect 23109 31331 23167 31337
rect 23109 31297 23121 31331
rect 23155 31297 23167 31331
rect 23109 31291 23167 31297
rect 7374 31260 7380 31272
rect 7335 31232 7380 31260
rect 7374 31220 7380 31232
rect 7432 31220 7438 31272
rect 7561 31263 7619 31269
rect 7561 31229 7573 31263
rect 7607 31260 7619 31263
rect 7742 31260 7748 31272
rect 7607 31232 7748 31260
rect 7607 31229 7619 31232
rect 7561 31223 7619 31229
rect 7742 31220 7748 31232
rect 7800 31220 7806 31272
rect 8665 31263 8723 31269
rect 8665 31229 8677 31263
rect 8711 31260 8723 31263
rect 9309 31263 9367 31269
rect 9309 31260 9321 31263
rect 8711 31232 9321 31260
rect 8711 31229 8723 31232
rect 8665 31223 8723 31229
rect 9309 31229 9321 31232
rect 9355 31260 9367 31263
rect 9355 31232 10180 31260
rect 9355 31229 9367 31232
rect 9309 31223 9367 31229
rect 9582 31152 9588 31204
rect 9640 31192 9646 31204
rect 9861 31195 9919 31201
rect 9861 31192 9873 31195
rect 9640 31164 9873 31192
rect 9640 31152 9646 31164
rect 9861 31161 9873 31164
rect 9907 31161 9919 31195
rect 10152 31192 10180 31232
rect 11054 31220 11060 31272
rect 11112 31260 11118 31272
rect 14185 31263 14243 31269
rect 14185 31260 14197 31263
rect 11112 31232 14197 31260
rect 11112 31220 11118 31232
rect 14185 31229 14197 31232
rect 14231 31229 14243 31263
rect 14185 31223 14243 31229
rect 14921 31263 14979 31269
rect 14921 31229 14933 31263
rect 14967 31260 14979 31263
rect 15562 31260 15568 31272
rect 14967 31232 15568 31260
rect 14967 31229 14979 31232
rect 14921 31223 14979 31229
rect 15562 31220 15568 31232
rect 15620 31220 15626 31272
rect 17586 31260 17592 31272
rect 17547 31232 17592 31260
rect 17586 31220 17592 31232
rect 17644 31220 17650 31272
rect 13449 31195 13507 31201
rect 10152 31164 13400 31192
rect 9861 31155 9919 31161
rect 1949 31127 2007 31133
rect 1949 31093 1961 31127
rect 1995 31124 2007 31127
rect 2498 31124 2504 31136
rect 1995 31096 2504 31124
rect 1995 31093 2007 31096
rect 1949 31087 2007 31093
rect 2498 31084 2504 31096
rect 2556 31084 2562 31136
rect 5442 31084 5448 31136
rect 5500 31124 5506 31136
rect 7745 31127 7803 31133
rect 7745 31124 7757 31127
rect 5500 31096 7757 31124
rect 5500 31084 5506 31096
rect 7745 31093 7757 31096
rect 7791 31124 7803 31127
rect 10410 31124 10416 31136
rect 7791 31096 10416 31124
rect 7791 31093 7803 31096
rect 7745 31087 7803 31093
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 10505 31127 10563 31133
rect 10505 31093 10517 31127
rect 10551 31124 10563 31127
rect 12066 31124 12072 31136
rect 10551 31096 12072 31124
rect 10551 31093 10563 31096
rect 10505 31087 10563 31093
rect 12066 31084 12072 31096
rect 12124 31084 12130 31136
rect 12345 31127 12403 31133
rect 12345 31093 12357 31127
rect 12391 31124 12403 31127
rect 13078 31124 13084 31136
rect 12391 31096 13084 31124
rect 12391 31093 12403 31096
rect 12345 31087 12403 31093
rect 13078 31084 13084 31096
rect 13136 31084 13142 31136
rect 13372 31124 13400 31164
rect 13449 31161 13461 31195
rect 13495 31192 13507 31195
rect 14550 31192 14556 31204
rect 13495 31164 14556 31192
rect 13495 31161 13507 31164
rect 13449 31155 13507 31161
rect 14550 31152 14556 31164
rect 14608 31152 14614 31204
rect 13722 31124 13728 31136
rect 13372 31096 13728 31124
rect 13722 31084 13728 31096
rect 13780 31084 13786 31136
rect 13814 31084 13820 31136
rect 13872 31124 13878 31136
rect 16117 31127 16175 31133
rect 16117 31124 16129 31127
rect 13872 31096 16129 31124
rect 13872 31084 13878 31096
rect 16117 31093 16129 31096
rect 16163 31093 16175 31127
rect 16117 31087 16175 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1946 30920 1952 30932
rect 1907 30892 1952 30920
rect 1946 30880 1952 30892
rect 2004 30880 2010 30932
rect 7742 30920 7748 30932
rect 7703 30892 7748 30920
rect 7742 30880 7748 30892
rect 7800 30880 7806 30932
rect 9217 30923 9275 30929
rect 9217 30889 9229 30923
rect 9263 30920 9275 30923
rect 10686 30920 10692 30932
rect 9263 30892 10692 30920
rect 9263 30889 9275 30892
rect 9217 30883 9275 30889
rect 10686 30880 10692 30892
rect 10744 30880 10750 30932
rect 12986 30880 12992 30932
rect 13044 30920 13050 30932
rect 13449 30923 13507 30929
rect 13449 30920 13461 30923
rect 13044 30892 13461 30920
rect 13044 30880 13050 30892
rect 13449 30889 13461 30892
rect 13495 30889 13507 30923
rect 13449 30883 13507 30889
rect 13722 30880 13728 30932
rect 13780 30920 13786 30932
rect 15654 30920 15660 30932
rect 13780 30892 15660 30920
rect 13780 30880 13786 30892
rect 15654 30880 15660 30892
rect 15712 30880 15718 30932
rect 20806 30920 20812 30932
rect 20767 30892 20812 30920
rect 20806 30880 20812 30892
rect 20864 30880 20870 30932
rect 22830 30920 22836 30932
rect 22791 30892 22836 30920
rect 22830 30880 22836 30892
rect 22888 30880 22894 30932
rect 8389 30855 8447 30861
rect 8389 30821 8401 30855
rect 8435 30821 8447 30855
rect 8389 30815 8447 30821
rect 5718 30784 5724 30796
rect 3252 30756 5724 30784
rect 2133 30719 2191 30725
rect 2133 30685 2145 30719
rect 2179 30716 2191 30719
rect 2593 30719 2651 30725
rect 2593 30716 2605 30719
rect 2179 30688 2605 30716
rect 2179 30685 2191 30688
rect 2133 30679 2191 30685
rect 2593 30685 2605 30688
rect 2639 30685 2651 30719
rect 2593 30679 2651 30685
rect 2608 30648 2636 30679
rect 2774 30676 2780 30728
rect 2832 30716 2838 30728
rect 3252 30725 3280 30756
rect 5718 30744 5724 30756
rect 5776 30744 5782 30796
rect 6549 30787 6607 30793
rect 6549 30753 6561 30787
rect 6595 30784 6607 30787
rect 7374 30784 7380 30796
rect 6595 30756 7380 30784
rect 6595 30753 6607 30756
rect 6549 30747 6607 30753
rect 7374 30744 7380 30756
rect 7432 30744 7438 30796
rect 3237 30719 3295 30725
rect 3237 30716 3249 30719
rect 2832 30688 3249 30716
rect 2832 30676 2838 30688
rect 3237 30685 3249 30688
rect 3283 30685 3295 30719
rect 3237 30679 3295 30685
rect 3878 30676 3884 30728
rect 3936 30716 3942 30728
rect 3973 30719 4031 30725
rect 3973 30716 3985 30719
rect 3936 30688 3985 30716
rect 3936 30676 3942 30688
rect 3973 30685 3985 30688
rect 4019 30685 4031 30719
rect 3973 30679 4031 30685
rect 7929 30719 7987 30725
rect 7929 30685 7941 30719
rect 7975 30716 7987 30719
rect 8404 30716 8432 30815
rect 11146 30812 11152 30864
rect 11204 30852 11210 30864
rect 13354 30852 13360 30864
rect 11204 30824 13360 30852
rect 11204 30812 11210 30824
rect 13354 30812 13360 30824
rect 13412 30812 13418 30864
rect 15013 30855 15071 30861
rect 15013 30821 15025 30855
rect 15059 30852 15071 30855
rect 19334 30852 19340 30864
rect 15059 30824 19340 30852
rect 15059 30821 15071 30824
rect 15013 30815 15071 30821
rect 10410 30744 10416 30796
rect 10468 30784 10474 30796
rect 11333 30787 11391 30793
rect 11333 30784 11345 30787
rect 10468 30756 11345 30784
rect 10468 30744 10474 30756
rect 11333 30753 11345 30756
rect 11379 30753 11391 30787
rect 11333 30747 11391 30753
rect 11977 30787 12035 30793
rect 11977 30753 11989 30787
rect 12023 30784 12035 30787
rect 15028 30784 15056 30815
rect 19334 30812 19340 30824
rect 19392 30812 19398 30864
rect 15562 30784 15568 30796
rect 12023 30756 15056 30784
rect 15523 30756 15568 30784
rect 12023 30753 12035 30756
rect 11977 30747 12035 30753
rect 15562 30744 15568 30756
rect 15620 30744 15626 30796
rect 15746 30784 15752 30796
rect 15707 30756 15752 30784
rect 15746 30744 15752 30756
rect 15804 30744 15810 30796
rect 23385 30787 23443 30793
rect 23385 30753 23397 30787
rect 23431 30784 23443 30787
rect 23842 30784 23848 30796
rect 23431 30756 23848 30784
rect 23431 30753 23443 30756
rect 23385 30747 23443 30753
rect 23842 30744 23848 30756
rect 23900 30744 23906 30796
rect 8570 30716 8576 30728
rect 7975 30688 8432 30716
rect 8531 30688 8576 30716
rect 7975 30685 7987 30688
rect 7929 30679 7987 30685
rect 8570 30676 8576 30688
rect 8628 30676 8634 30728
rect 9398 30716 9404 30728
rect 9359 30688 9404 30716
rect 9398 30676 9404 30688
rect 9456 30716 9462 30728
rect 9861 30719 9919 30725
rect 9861 30716 9873 30719
rect 9456 30688 9873 30716
rect 9456 30676 9462 30688
rect 9861 30685 9873 30688
rect 9907 30685 9919 30719
rect 9861 30679 9919 30685
rect 10134 30676 10140 30728
rect 10192 30716 10198 30728
rect 10594 30716 10600 30728
rect 10192 30688 10600 30716
rect 10192 30676 10198 30688
rect 10594 30676 10600 30688
rect 10652 30676 10658 30728
rect 13354 30716 13360 30728
rect 13315 30688 13360 30716
rect 13354 30676 13360 30688
rect 13412 30676 13418 30728
rect 16574 30676 16580 30728
rect 16632 30716 16638 30728
rect 17129 30719 17187 30725
rect 17129 30716 17141 30719
rect 16632 30688 17141 30716
rect 16632 30676 16638 30688
rect 17129 30685 17141 30688
rect 17175 30716 17187 30719
rect 17862 30716 17868 30728
rect 17175 30688 17868 30716
rect 17175 30685 17187 30688
rect 17129 30679 17187 30685
rect 17862 30676 17868 30688
rect 17920 30676 17926 30728
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30716 19763 30719
rect 19978 30716 19984 30728
rect 19751 30688 19984 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 19978 30676 19984 30688
rect 20036 30676 20042 30728
rect 20349 30719 20407 30725
rect 20349 30685 20361 30719
rect 20395 30685 20407 30719
rect 20349 30679 20407 30685
rect 4614 30648 4620 30660
rect 2608 30620 4620 30648
rect 4614 30608 4620 30620
rect 4672 30608 4678 30660
rect 6638 30608 6644 30660
rect 6696 30648 6702 30660
rect 7193 30651 7251 30657
rect 6696 30620 6741 30648
rect 6696 30608 6702 30620
rect 7193 30617 7205 30651
rect 7239 30648 7251 30651
rect 7466 30648 7472 30660
rect 7239 30620 7472 30648
rect 7239 30617 7251 30620
rect 7193 30611 7251 30617
rect 7466 30608 7472 30620
rect 7524 30608 7530 30660
rect 9953 30651 10011 30657
rect 9953 30617 9965 30651
rect 9999 30648 10011 30651
rect 11146 30648 11152 30660
rect 9999 30620 11152 30648
rect 9999 30617 10011 30620
rect 9953 30611 10011 30617
rect 11146 30608 11152 30620
rect 11204 30608 11210 30660
rect 11425 30651 11483 30657
rect 11425 30617 11437 30651
rect 11471 30617 11483 30651
rect 14458 30648 14464 30660
rect 14419 30620 14464 30648
rect 11425 30611 11483 30617
rect 2406 30540 2412 30592
rect 2464 30580 2470 30592
rect 2685 30583 2743 30589
rect 2685 30580 2697 30583
rect 2464 30552 2697 30580
rect 2464 30540 2470 30552
rect 2685 30549 2697 30552
rect 2731 30549 2743 30583
rect 2685 30543 2743 30549
rect 3142 30540 3148 30592
rect 3200 30580 3206 30592
rect 3329 30583 3387 30589
rect 3329 30580 3341 30583
rect 3200 30552 3341 30580
rect 3200 30540 3206 30552
rect 3329 30549 3341 30552
rect 3375 30549 3387 30583
rect 4154 30580 4160 30592
rect 4115 30552 4160 30580
rect 3329 30543 3387 30549
rect 4154 30540 4160 30552
rect 4212 30540 4218 30592
rect 10689 30583 10747 30589
rect 10689 30549 10701 30583
rect 10735 30580 10747 30583
rect 11440 30580 11468 30611
rect 14458 30608 14464 30620
rect 14516 30608 14522 30660
rect 14550 30608 14556 30660
rect 14608 30648 14614 30660
rect 20364 30648 20392 30679
rect 20438 30676 20444 30728
rect 20496 30716 20502 30728
rect 20993 30719 21051 30725
rect 20993 30716 21005 30719
rect 20496 30688 21005 30716
rect 20496 30676 20502 30688
rect 20993 30685 21005 30688
rect 21039 30685 21051 30719
rect 22738 30716 22744 30728
rect 22699 30688 22744 30716
rect 20993 30679 21051 30685
rect 22738 30676 22744 30688
rect 22796 30676 22802 30728
rect 23566 30716 23572 30728
rect 23527 30688 23572 30716
rect 23566 30676 23572 30688
rect 23624 30676 23630 30728
rect 28261 30719 28319 30725
rect 28261 30685 28273 30719
rect 28307 30716 28319 30719
rect 32398 30716 32404 30728
rect 28307 30688 32404 30716
rect 28307 30685 28319 30688
rect 28261 30679 28319 30685
rect 32398 30676 32404 30688
rect 32456 30676 32462 30728
rect 14608 30620 14653 30648
rect 19536 30620 20392 30648
rect 14608 30608 14614 30620
rect 10735 30552 11468 30580
rect 14476 30580 14504 30608
rect 16209 30583 16267 30589
rect 16209 30580 16221 30583
rect 14476 30552 16221 30580
rect 10735 30549 10747 30552
rect 10689 30543 10747 30549
rect 16209 30549 16221 30552
rect 16255 30549 16267 30583
rect 16209 30543 16267 30549
rect 16945 30583 17003 30589
rect 16945 30549 16957 30583
rect 16991 30580 17003 30583
rect 17310 30580 17316 30592
rect 16991 30552 17316 30580
rect 16991 30549 17003 30552
rect 16945 30543 17003 30549
rect 17310 30540 17316 30552
rect 17368 30540 17374 30592
rect 19536 30589 19564 30620
rect 19521 30583 19579 30589
rect 19521 30549 19533 30583
rect 19567 30549 19579 30583
rect 20162 30580 20168 30592
rect 20123 30552 20168 30580
rect 19521 30543 19579 30549
rect 20162 30540 20168 30552
rect 20220 30540 20226 30592
rect 24026 30580 24032 30592
rect 23987 30552 24032 30580
rect 24026 30540 24032 30552
rect 24084 30540 24090 30592
rect 27890 30540 27896 30592
rect 27948 30580 27954 30592
rect 28353 30583 28411 30589
rect 28353 30580 28365 30583
rect 27948 30552 28365 30580
rect 27948 30540 27954 30552
rect 28353 30549 28365 30552
rect 28399 30549 28411 30583
rect 28353 30543 28411 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 9582 30336 9588 30388
rect 9640 30376 9646 30388
rect 9640 30348 11008 30376
rect 9640 30336 9646 30348
rect 3973 30311 4031 30317
rect 3973 30277 3985 30311
rect 4019 30308 4031 30311
rect 5442 30308 5448 30320
rect 4019 30280 5448 30308
rect 4019 30277 4031 30280
rect 3973 30271 4031 30277
rect 5442 30268 5448 30280
rect 5500 30268 5506 30320
rect 6914 30268 6920 30320
rect 6972 30308 6978 30320
rect 7009 30311 7067 30317
rect 7009 30308 7021 30311
rect 6972 30280 7021 30308
rect 6972 30268 6978 30280
rect 7009 30277 7021 30280
rect 7055 30277 7067 30311
rect 7009 30271 7067 30277
rect 8570 30268 8576 30320
rect 8628 30308 8634 30320
rect 9490 30308 9496 30320
rect 8628 30280 9496 30308
rect 8628 30268 8634 30280
rect 9490 30268 9496 30280
rect 9548 30268 9554 30320
rect 10870 30308 10876 30320
rect 10831 30280 10876 30308
rect 10870 30268 10876 30280
rect 10928 30268 10934 30320
rect 10980 30308 11008 30348
rect 10980 30280 14688 30308
rect 1762 30240 1768 30252
rect 1723 30212 1768 30240
rect 1762 30200 1768 30212
rect 1820 30200 1826 30252
rect 2590 30200 2596 30252
rect 2648 30240 2654 30252
rect 2685 30243 2743 30249
rect 2685 30240 2697 30243
rect 2648 30212 2697 30240
rect 2648 30200 2654 30212
rect 2685 30209 2697 30212
rect 2731 30209 2743 30243
rect 2685 30203 2743 30209
rect 2777 30243 2835 30249
rect 2777 30209 2789 30243
rect 2823 30240 2835 30243
rect 3513 30243 3571 30249
rect 3513 30240 3525 30243
rect 2823 30212 3525 30240
rect 2823 30209 2835 30212
rect 2777 30203 2835 30209
rect 3513 30209 3525 30212
rect 3559 30209 3571 30243
rect 5994 30240 6000 30252
rect 5955 30212 6000 30240
rect 3513 30203 3571 30209
rect 5994 30200 6000 30212
rect 6052 30200 6058 30252
rect 9217 30243 9275 30249
rect 9217 30209 9229 30243
rect 9263 30209 9275 30243
rect 9217 30203 9275 30209
rect 3329 30175 3387 30181
rect 3329 30141 3341 30175
rect 3375 30172 3387 30175
rect 4154 30172 4160 30184
rect 3375 30144 4160 30172
rect 3375 30141 3387 30144
rect 3329 30135 3387 30141
rect 4154 30132 4160 30144
rect 4212 30132 4218 30184
rect 4433 30175 4491 30181
rect 4433 30141 4445 30175
rect 4479 30141 4491 30175
rect 4433 30135 4491 30141
rect 6917 30175 6975 30181
rect 6917 30141 6929 30175
rect 6963 30172 6975 30175
rect 9232 30172 9260 30203
rect 10686 30200 10692 30252
rect 10744 30240 10750 30252
rect 10781 30243 10839 30249
rect 10781 30240 10793 30243
rect 10744 30212 10793 30240
rect 10744 30200 10750 30212
rect 10781 30209 10793 30212
rect 10827 30209 10839 30243
rect 10781 30203 10839 30209
rect 12342 30200 12348 30252
rect 12400 30240 12406 30252
rect 12437 30243 12495 30249
rect 12437 30240 12449 30243
rect 12400 30212 12449 30240
rect 12400 30200 12406 30212
rect 12437 30209 12449 30212
rect 12483 30209 12495 30243
rect 12437 30203 12495 30209
rect 13173 30243 13231 30249
rect 13173 30209 13185 30243
rect 13219 30209 13231 30243
rect 13173 30203 13231 30209
rect 13817 30243 13875 30249
rect 13817 30209 13829 30243
rect 13863 30240 13875 30243
rect 14090 30240 14096 30252
rect 13863 30212 14096 30240
rect 13863 30209 13875 30212
rect 13817 30203 13875 30209
rect 11330 30172 11336 30184
rect 6963 30144 9168 30172
rect 9232 30144 11336 30172
rect 6963 30141 6975 30144
rect 6917 30135 6975 30141
rect 2774 30064 2780 30116
rect 2832 30104 2838 30116
rect 4448 30104 4476 30135
rect 7466 30104 7472 30116
rect 2832 30076 4476 30104
rect 7427 30076 7472 30104
rect 2832 30064 2838 30076
rect 7466 30064 7472 30076
rect 7524 30064 7530 30116
rect 9140 30104 9168 30144
rect 11330 30132 11336 30144
rect 11388 30132 11394 30184
rect 13188 30172 13216 30203
rect 14090 30200 14096 30212
rect 14148 30200 14154 30252
rect 14182 30172 14188 30184
rect 11440 30144 14188 30172
rect 11054 30104 11060 30116
rect 9140 30076 11060 30104
rect 11054 30064 11060 30076
rect 11112 30064 11118 30116
rect 1578 30036 1584 30048
rect 1539 30008 1584 30036
rect 1578 29996 1584 30008
rect 1636 29996 1642 30048
rect 5813 30039 5871 30045
rect 5813 30005 5825 30039
rect 5859 30036 5871 30039
rect 6362 30036 6368 30048
rect 5859 30008 6368 30036
rect 5859 30005 5871 30008
rect 5813 29999 5871 30005
rect 6362 29996 6368 30008
rect 6420 29996 6426 30048
rect 9306 30036 9312 30048
rect 9267 30008 9312 30036
rect 9306 29996 9312 30008
rect 9364 29996 9370 30048
rect 9490 29996 9496 30048
rect 9548 30036 9554 30048
rect 11440 30036 11468 30144
rect 14182 30132 14188 30144
rect 14240 30132 14246 30184
rect 14660 30172 14688 30280
rect 16758 30268 16764 30320
rect 16816 30308 16822 30320
rect 17037 30311 17095 30317
rect 17037 30308 17049 30311
rect 16816 30280 17049 30308
rect 16816 30268 16822 30280
rect 17037 30277 17049 30280
rect 17083 30277 17095 30311
rect 17586 30308 17592 30320
rect 17547 30280 17592 30308
rect 17037 30271 17095 30277
rect 17586 30268 17592 30280
rect 17644 30268 17650 30320
rect 31573 30311 31631 30317
rect 31573 30277 31585 30311
rect 31619 30308 31631 30311
rect 34514 30308 34520 30320
rect 31619 30280 34520 30308
rect 31619 30277 31631 30280
rect 31573 30271 31631 30277
rect 34514 30268 34520 30280
rect 34572 30268 34578 30320
rect 17862 30200 17868 30252
rect 17920 30240 17926 30252
rect 18049 30243 18107 30249
rect 18049 30240 18061 30243
rect 17920 30212 18061 30240
rect 17920 30200 17926 30212
rect 18049 30209 18061 30212
rect 18095 30209 18107 30243
rect 18049 30203 18107 30209
rect 21910 30200 21916 30252
rect 21968 30240 21974 30252
rect 22005 30243 22063 30249
rect 22005 30240 22017 30243
rect 21968 30212 22017 30240
rect 21968 30200 21974 30212
rect 22005 30209 22017 30212
rect 22051 30240 22063 30243
rect 22462 30240 22468 30252
rect 22051 30212 22468 30240
rect 22051 30209 22063 30212
rect 22005 30203 22063 30209
rect 22462 30200 22468 30212
rect 22520 30200 22526 30252
rect 30466 30200 30472 30252
rect 30524 30240 30530 30252
rect 31481 30243 31539 30249
rect 31481 30240 31493 30243
rect 30524 30212 31493 30240
rect 30524 30200 30530 30212
rect 31481 30209 31493 30212
rect 31527 30209 31539 30243
rect 31481 30203 31539 30209
rect 31754 30200 31760 30252
rect 31812 30240 31818 30252
rect 33321 30243 33379 30249
rect 33321 30240 33333 30243
rect 31812 30212 33333 30240
rect 31812 30200 31818 30212
rect 33321 30209 33333 30212
rect 33367 30209 33379 30243
rect 33321 30203 33379 30209
rect 33413 30243 33471 30249
rect 33413 30209 33425 30243
rect 33459 30240 33471 30243
rect 34333 30243 34391 30249
rect 34333 30240 34345 30243
rect 33459 30212 34345 30240
rect 33459 30209 33471 30212
rect 33413 30203 33471 30209
rect 34333 30209 34345 30212
rect 34379 30209 34391 30243
rect 38013 30243 38071 30249
rect 38013 30240 38025 30243
rect 34333 30203 34391 30209
rect 35866 30212 38025 30240
rect 16945 30175 17003 30181
rect 16945 30172 16957 30175
rect 14660 30144 16957 30172
rect 16945 30141 16957 30144
rect 16991 30141 17003 30175
rect 16945 30135 17003 30141
rect 11698 30064 11704 30116
rect 11756 30104 11762 30116
rect 14274 30104 14280 30116
rect 11756 30076 14280 30104
rect 11756 30064 11762 30076
rect 14274 30064 14280 30076
rect 14332 30064 14338 30116
rect 34149 30107 34207 30113
rect 34149 30073 34161 30107
rect 34195 30104 34207 30107
rect 35866 30104 35894 30212
rect 38013 30209 38025 30212
rect 38059 30209 38071 30243
rect 38013 30203 38071 30209
rect 34195 30076 35894 30104
rect 34195 30073 34207 30076
rect 34149 30067 34207 30073
rect 9548 30008 11468 30036
rect 9548 29996 9554 30008
rect 11514 29996 11520 30048
rect 11572 30036 11578 30048
rect 12253 30039 12311 30045
rect 12253 30036 12265 30039
rect 11572 30008 12265 30036
rect 11572 29996 11578 30008
rect 12253 30005 12265 30008
rect 12299 30005 12311 30039
rect 12253 29999 12311 30005
rect 13170 29996 13176 30048
rect 13228 30036 13234 30048
rect 13265 30039 13323 30045
rect 13265 30036 13277 30039
rect 13228 30008 13277 30036
rect 13228 29996 13234 30008
rect 13265 30005 13277 30008
rect 13311 30005 13323 30039
rect 13906 30036 13912 30048
rect 13867 30008 13912 30036
rect 13265 29999 13323 30005
rect 13906 29996 13912 30008
rect 13964 29996 13970 30048
rect 18141 30039 18199 30045
rect 18141 30005 18153 30039
rect 18187 30036 18199 30039
rect 18966 30036 18972 30048
rect 18187 30008 18972 30036
rect 18187 30005 18199 30008
rect 18141 29999 18199 30005
rect 18966 29996 18972 30008
rect 19024 29996 19030 30048
rect 21634 29996 21640 30048
rect 21692 30036 21698 30048
rect 22097 30039 22155 30045
rect 22097 30036 22109 30039
rect 21692 30008 22109 30036
rect 21692 29996 21698 30008
rect 22097 30005 22109 30008
rect 22143 30005 22155 30039
rect 38194 30036 38200 30048
rect 38155 30008 38200 30036
rect 22097 29999 22155 30005
rect 38194 29996 38200 30008
rect 38252 29996 38258 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 6181 29835 6239 29841
rect 6181 29801 6193 29835
rect 6227 29832 6239 29835
rect 6638 29832 6644 29844
rect 6227 29804 6644 29832
rect 6227 29801 6239 29804
rect 6181 29795 6239 29801
rect 6638 29792 6644 29804
rect 6696 29792 6702 29844
rect 6914 29832 6920 29844
rect 6875 29804 6920 29832
rect 6914 29792 6920 29804
rect 6972 29792 6978 29844
rect 9122 29792 9128 29844
rect 9180 29832 9186 29844
rect 18785 29835 18843 29841
rect 9180 29804 17540 29832
rect 9180 29792 9186 29804
rect 4065 29767 4123 29773
rect 4065 29733 4077 29767
rect 4111 29764 4123 29767
rect 4111 29736 12434 29764
rect 4111 29733 4123 29736
rect 4065 29727 4123 29733
rect 2774 29656 2780 29708
rect 2832 29696 2838 29708
rect 3050 29696 3056 29708
rect 2832 29668 2877 29696
rect 3011 29668 3056 29696
rect 2832 29656 2838 29668
rect 3050 29656 3056 29668
rect 3108 29656 3114 29708
rect 5994 29656 6000 29708
rect 6052 29696 6058 29708
rect 9306 29696 9312 29708
rect 6052 29668 6868 29696
rect 9267 29668 9312 29696
rect 6052 29656 6058 29668
rect 1854 29628 1860 29640
rect 1815 29600 1860 29628
rect 1854 29588 1860 29600
rect 1912 29588 1918 29640
rect 3970 29628 3976 29640
rect 3931 29600 3976 29628
rect 3970 29588 3976 29600
rect 4028 29588 4034 29640
rect 6362 29628 6368 29640
rect 6323 29600 6368 29628
rect 6362 29588 6368 29600
rect 6420 29588 6426 29640
rect 6840 29637 6868 29668
rect 9306 29656 9312 29668
rect 9364 29656 9370 29708
rect 11514 29696 11520 29708
rect 11475 29668 11520 29696
rect 11514 29656 11520 29668
rect 11572 29656 11578 29708
rect 12406 29696 12434 29736
rect 12529 29699 12587 29705
rect 12529 29696 12541 29699
rect 12406 29668 12541 29696
rect 12529 29665 12541 29668
rect 12575 29696 12587 29699
rect 12986 29696 12992 29708
rect 12575 29668 12992 29696
rect 12575 29665 12587 29668
rect 12529 29659 12587 29665
rect 12986 29656 12992 29668
rect 13044 29656 13050 29708
rect 17512 29696 17540 29804
rect 18785 29801 18797 29835
rect 18831 29832 18843 29835
rect 20438 29832 20444 29844
rect 18831 29804 20444 29832
rect 18831 29801 18843 29804
rect 18785 29795 18843 29801
rect 20438 29792 20444 29804
rect 20496 29792 20502 29844
rect 21358 29792 21364 29844
rect 21416 29832 21422 29844
rect 21821 29835 21879 29841
rect 21821 29832 21833 29835
rect 21416 29804 21833 29832
rect 21416 29792 21422 29804
rect 21821 29801 21833 29804
rect 21867 29801 21879 29835
rect 21821 29795 21879 29801
rect 23109 29835 23167 29841
rect 23109 29801 23121 29835
rect 23155 29832 23167 29835
rect 23566 29832 23572 29844
rect 23155 29804 23572 29832
rect 23155 29801 23167 29804
rect 23109 29795 23167 29801
rect 23566 29792 23572 29804
rect 23624 29792 23630 29844
rect 23842 29832 23848 29844
rect 23803 29804 23848 29832
rect 23842 29792 23848 29804
rect 23900 29792 23906 29844
rect 19429 29699 19487 29705
rect 19429 29696 19441 29699
rect 17512 29668 19441 29696
rect 19429 29665 19441 29668
rect 19475 29665 19487 29699
rect 19429 29659 19487 29665
rect 19613 29699 19671 29705
rect 19613 29665 19625 29699
rect 19659 29696 19671 29699
rect 20162 29696 20168 29708
rect 19659 29668 20168 29696
rect 19659 29665 19671 29668
rect 19613 29659 19671 29665
rect 6825 29631 6883 29637
rect 6825 29597 6837 29631
rect 6871 29597 6883 29631
rect 6825 29591 6883 29597
rect 7469 29631 7527 29637
rect 7469 29597 7481 29631
rect 7515 29628 7527 29631
rect 7742 29628 7748 29640
rect 7515 29600 7748 29628
rect 7515 29597 7527 29600
rect 7469 29591 7527 29597
rect 7742 29588 7748 29600
rect 7800 29588 7806 29640
rect 9122 29628 9128 29640
rect 9083 29600 9128 29628
rect 9122 29588 9128 29600
rect 9180 29588 9186 29640
rect 11238 29588 11244 29640
rect 11296 29628 11302 29640
rect 11333 29631 11391 29637
rect 11333 29628 11345 29631
rect 11296 29600 11345 29628
rect 11296 29588 11302 29600
rect 11333 29597 11345 29600
rect 11379 29597 11391 29631
rect 14274 29628 14280 29640
rect 14235 29600 14280 29628
rect 11333 29591 11391 29597
rect 2866 29520 2872 29572
rect 2924 29560 2930 29572
rect 11348 29560 11376 29591
rect 14274 29588 14280 29600
rect 14332 29588 14338 29640
rect 17310 29628 17316 29640
rect 17271 29600 17316 29628
rect 17310 29588 17316 29600
rect 17368 29588 17374 29640
rect 18693 29631 18751 29637
rect 18693 29597 18705 29631
rect 18739 29628 18751 29631
rect 19150 29628 19156 29640
rect 18739 29600 19156 29628
rect 18739 29597 18751 29600
rect 18693 29591 18751 29597
rect 19150 29588 19156 29600
rect 19208 29588 19214 29640
rect 19444 29628 19472 29659
rect 20162 29656 20168 29668
rect 20220 29656 20226 29708
rect 21634 29696 21640 29708
rect 21595 29668 21640 29696
rect 21634 29656 21640 29668
rect 21692 29656 21698 29708
rect 20622 29628 20628 29640
rect 19444 29600 20628 29628
rect 20622 29588 20628 29600
rect 20680 29588 20686 29640
rect 20809 29631 20867 29637
rect 20809 29597 20821 29631
rect 20855 29628 20867 29631
rect 20990 29628 20996 29640
rect 20855 29600 20996 29628
rect 20855 29597 20867 29600
rect 20809 29591 20867 29597
rect 20990 29588 20996 29600
rect 21048 29588 21054 29640
rect 21453 29631 21511 29637
rect 21453 29597 21465 29631
rect 21499 29597 21511 29631
rect 23014 29628 23020 29640
rect 22975 29600 23020 29628
rect 21453 29591 21511 29597
rect 11514 29560 11520 29572
rect 2924 29532 2969 29560
rect 11348 29532 11520 29560
rect 2924 29520 2930 29532
rect 11514 29520 11520 29532
rect 11572 29520 11578 29572
rect 12621 29563 12679 29569
rect 12621 29529 12633 29563
rect 12667 29529 12679 29563
rect 12621 29523 12679 29529
rect 1949 29495 2007 29501
rect 1949 29461 1961 29495
rect 1995 29492 2007 29495
rect 2130 29492 2136 29504
rect 1995 29464 2136 29492
rect 1995 29461 2007 29464
rect 1949 29455 2007 29461
rect 2130 29452 2136 29464
rect 2188 29452 2194 29504
rect 7558 29492 7564 29504
rect 7519 29464 7564 29492
rect 7558 29452 7564 29464
rect 7616 29452 7622 29504
rect 9769 29495 9827 29501
rect 9769 29461 9781 29495
rect 9815 29492 9827 29495
rect 10502 29492 10508 29504
rect 9815 29464 10508 29492
rect 9815 29461 9827 29464
rect 9769 29455 9827 29461
rect 10502 29452 10508 29464
rect 10560 29492 10566 29504
rect 11977 29495 12035 29501
rect 11977 29492 11989 29495
rect 10560 29464 11989 29492
rect 10560 29452 10566 29464
rect 11977 29461 11989 29464
rect 12023 29461 12035 29495
rect 11977 29455 12035 29461
rect 12066 29452 12072 29504
rect 12124 29492 12130 29504
rect 12636 29492 12664 29523
rect 12802 29520 12808 29572
rect 12860 29560 12866 29572
rect 13173 29563 13231 29569
rect 13173 29560 13185 29563
rect 12860 29532 13185 29560
rect 12860 29520 12866 29532
rect 13173 29529 13185 29532
rect 13219 29529 13231 29563
rect 21468 29560 21496 29591
rect 23014 29588 23020 29600
rect 23072 29588 23078 29640
rect 23750 29628 23756 29640
rect 23711 29600 23756 29628
rect 23750 29588 23756 29600
rect 23808 29588 23814 29640
rect 24026 29560 24032 29572
rect 21468 29532 24032 29560
rect 13173 29523 13231 29529
rect 24026 29520 24032 29532
rect 24084 29520 24090 29572
rect 14366 29492 14372 29504
rect 12124 29464 12664 29492
rect 14327 29464 14372 29492
rect 12124 29452 12130 29464
rect 14366 29452 14372 29464
rect 14424 29452 14430 29504
rect 17126 29492 17132 29504
rect 17087 29464 17132 29492
rect 17126 29452 17132 29464
rect 17184 29452 17190 29504
rect 20070 29492 20076 29504
rect 20031 29464 20076 29492
rect 20070 29452 20076 29464
rect 20128 29452 20134 29504
rect 20901 29495 20959 29501
rect 20901 29461 20913 29495
rect 20947 29492 20959 29495
rect 22186 29492 22192 29504
rect 20947 29464 22192 29492
rect 20947 29461 20959 29464
rect 20901 29455 20959 29461
rect 22186 29452 22192 29464
rect 22244 29452 22250 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 5261 29291 5319 29297
rect 5261 29257 5273 29291
rect 5307 29288 5319 29291
rect 9122 29288 9128 29300
rect 5307 29260 9128 29288
rect 5307 29257 5319 29260
rect 5261 29251 5319 29257
rect 9122 29248 9128 29260
rect 9180 29248 9186 29300
rect 12342 29288 12348 29300
rect 12303 29260 12348 29288
rect 12342 29248 12348 29260
rect 12400 29248 12406 29300
rect 12526 29248 12532 29300
rect 12584 29288 12590 29300
rect 12802 29288 12808 29300
rect 12584 29260 12808 29288
rect 12584 29248 12590 29260
rect 12802 29248 12808 29260
rect 12860 29248 12866 29300
rect 13633 29291 13691 29297
rect 13633 29257 13645 29291
rect 13679 29288 13691 29291
rect 14458 29288 14464 29300
rect 13679 29260 14464 29288
rect 13679 29257 13691 29260
rect 13633 29251 13691 29257
rect 14458 29248 14464 29260
rect 14516 29248 14522 29300
rect 30469 29291 30527 29297
rect 30469 29257 30481 29291
rect 30515 29288 30527 29291
rect 36446 29288 36452 29300
rect 30515 29260 36452 29288
rect 30515 29257 30527 29260
rect 30469 29251 30527 29257
rect 36446 29248 36452 29260
rect 36504 29248 36510 29300
rect 8570 29220 8576 29232
rect 5460 29192 8576 29220
rect 1762 29152 1768 29164
rect 1723 29124 1768 29152
rect 1762 29112 1768 29124
rect 1820 29112 1826 29164
rect 2314 29112 2320 29164
rect 2372 29152 2378 29164
rect 5169 29155 5227 29161
rect 5169 29152 5181 29155
rect 2372 29124 5181 29152
rect 2372 29112 2378 29124
rect 5169 29121 5181 29124
rect 5215 29121 5227 29155
rect 5169 29115 5227 29121
rect 2590 29044 2596 29096
rect 2648 29084 2654 29096
rect 5460 29084 5488 29192
rect 8570 29180 8576 29192
rect 8628 29180 8634 29232
rect 10594 29220 10600 29232
rect 10555 29192 10600 29220
rect 10594 29180 10600 29192
rect 10652 29180 10658 29232
rect 5534 29112 5540 29164
rect 5592 29152 5598 29164
rect 6641 29155 6699 29161
rect 6641 29152 6653 29155
rect 5592 29124 6653 29152
rect 5592 29112 5598 29124
rect 6641 29121 6653 29124
rect 6687 29121 6699 29155
rect 6641 29115 6699 29121
rect 7653 29155 7711 29161
rect 7653 29121 7665 29155
rect 7699 29152 7711 29155
rect 9858 29152 9864 29164
rect 7699 29124 9720 29152
rect 9819 29124 9864 29152
rect 7699 29121 7711 29124
rect 7653 29115 7711 29121
rect 2648 29056 5488 29084
rect 6733 29087 6791 29093
rect 2648 29044 2654 29056
rect 6733 29053 6745 29087
rect 6779 29084 6791 29087
rect 8202 29084 8208 29096
rect 6779 29056 8208 29084
rect 6779 29053 6791 29056
rect 6733 29047 6791 29053
rect 8202 29044 8208 29056
rect 8260 29044 8266 29096
rect 6822 28976 6828 29028
rect 6880 29016 6886 29028
rect 9692 29025 9720 29124
rect 9858 29112 9864 29124
rect 9916 29112 9922 29164
rect 11330 29112 11336 29164
rect 11388 29152 11394 29164
rect 12434 29152 12440 29164
rect 11388 29124 12440 29152
rect 11388 29112 11394 29124
rect 12434 29112 12440 29124
rect 12492 29152 12498 29164
rect 12529 29155 12587 29161
rect 12529 29152 12541 29155
rect 12492 29124 12541 29152
rect 12492 29112 12498 29124
rect 12529 29121 12541 29124
rect 12575 29121 12587 29155
rect 13170 29152 13176 29164
rect 13131 29124 13176 29152
rect 12529 29115 12587 29121
rect 13170 29112 13176 29124
rect 13228 29112 13234 29164
rect 14090 29112 14096 29164
rect 14148 29152 14154 29164
rect 15197 29155 15255 29161
rect 15197 29152 15209 29155
rect 14148 29124 15209 29152
rect 14148 29112 14154 29124
rect 15197 29121 15209 29124
rect 15243 29121 15255 29155
rect 15197 29115 15255 29121
rect 16209 29155 16267 29161
rect 16209 29121 16221 29155
rect 16255 29152 16267 29155
rect 16850 29152 16856 29164
rect 16255 29124 16856 29152
rect 16255 29121 16267 29124
rect 16209 29115 16267 29121
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 18966 29152 18972 29164
rect 18927 29124 18972 29152
rect 18966 29112 18972 29124
rect 19024 29112 19030 29164
rect 25314 29152 25320 29164
rect 25275 29124 25320 29152
rect 25314 29112 25320 29124
rect 25372 29112 25378 29164
rect 27982 29112 27988 29164
rect 28040 29152 28046 29164
rect 30377 29155 30435 29161
rect 30377 29152 30389 29155
rect 28040 29124 30389 29152
rect 28040 29112 28046 29124
rect 30377 29121 30389 29124
rect 30423 29121 30435 29155
rect 30377 29115 30435 29121
rect 36630 29112 36636 29164
rect 36688 29152 36694 29164
rect 38013 29155 38071 29161
rect 38013 29152 38025 29155
rect 36688 29124 38025 29152
rect 36688 29112 36694 29124
rect 38013 29121 38025 29124
rect 38059 29121 38071 29155
rect 38013 29115 38071 29121
rect 10502 29084 10508 29096
rect 10463 29056 10508 29084
rect 10502 29044 10508 29056
rect 10560 29044 10566 29096
rect 10686 29044 10692 29096
rect 10744 29084 10750 29096
rect 10781 29087 10839 29093
rect 10781 29084 10793 29087
rect 10744 29056 10793 29084
rect 10744 29044 10750 29056
rect 10781 29053 10793 29056
rect 10827 29053 10839 29087
rect 12986 29084 12992 29096
rect 12947 29056 12992 29084
rect 10781 29047 10839 29053
rect 12986 29044 12992 29056
rect 13044 29044 13050 29096
rect 18785 29087 18843 29093
rect 18785 29053 18797 29087
rect 18831 29084 18843 29087
rect 20070 29084 20076 29096
rect 18831 29056 20076 29084
rect 18831 29053 18843 29056
rect 18785 29047 18843 29053
rect 20070 29044 20076 29056
rect 20128 29044 20134 29096
rect 23385 29087 23443 29093
rect 23385 29053 23397 29087
rect 23431 29084 23443 29087
rect 24029 29087 24087 29093
rect 24029 29084 24041 29087
rect 23431 29056 24041 29084
rect 23431 29053 23443 29056
rect 23385 29047 23443 29053
rect 24029 29053 24041 29056
rect 24075 29053 24087 29087
rect 24210 29084 24216 29096
rect 24171 29056 24216 29084
rect 24029 29047 24087 29053
rect 24210 29044 24216 29056
rect 24268 29044 24274 29096
rect 7469 29019 7527 29025
rect 7469 29016 7481 29019
rect 6880 28988 7481 29016
rect 6880 28976 6886 28988
rect 7469 28985 7481 28988
rect 7515 28985 7527 29019
rect 7469 28979 7527 28985
rect 9677 29019 9735 29025
rect 9677 28985 9689 29019
rect 9723 28985 9735 29019
rect 19150 29016 19156 29028
rect 19111 28988 19156 29016
rect 9677 28979 9735 28985
rect 19150 28976 19156 28988
rect 19208 28976 19214 29028
rect 38194 29016 38200 29028
rect 38155 28988 38200 29016
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 1581 28951 1639 28957
rect 1581 28917 1593 28951
rect 1627 28948 1639 28951
rect 1946 28948 1952 28960
rect 1627 28920 1952 28948
rect 1627 28917 1639 28920
rect 1581 28911 1639 28917
rect 1946 28908 1952 28920
rect 2004 28908 2010 28960
rect 15010 28948 15016 28960
rect 14971 28920 15016 28948
rect 15010 28908 15016 28920
rect 15068 28908 15074 28960
rect 16022 28948 16028 28960
rect 15983 28920 16028 28948
rect 16022 28908 16028 28920
rect 16080 28908 16086 28960
rect 24670 28948 24676 28960
rect 24631 28920 24676 28948
rect 24670 28908 24676 28920
rect 24728 28908 24734 28960
rect 24946 28908 24952 28960
rect 25004 28948 25010 28960
rect 25133 28951 25191 28957
rect 25133 28948 25145 28951
rect 25004 28920 25145 28948
rect 25004 28908 25010 28920
rect 25133 28917 25145 28920
rect 25179 28917 25191 28951
rect 25133 28911 25191 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 10594 28744 10600 28756
rect 10555 28716 10600 28744
rect 10594 28704 10600 28716
rect 10652 28704 10658 28756
rect 16850 28744 16856 28756
rect 16811 28716 16856 28744
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 20070 28744 20076 28756
rect 20031 28716 20076 28744
rect 20070 28704 20076 28716
rect 20128 28704 20134 28756
rect 24210 28704 24216 28756
rect 24268 28744 24274 28756
rect 24765 28747 24823 28753
rect 24765 28744 24777 28747
rect 24268 28716 24777 28744
rect 24268 28704 24274 28716
rect 24765 28713 24777 28716
rect 24811 28713 24823 28747
rect 24765 28707 24823 28713
rect 9769 28679 9827 28685
rect 9769 28645 9781 28679
rect 9815 28676 9827 28679
rect 17586 28676 17592 28688
rect 9815 28648 17592 28676
rect 9815 28645 9827 28648
rect 9769 28639 9827 28645
rect 17586 28636 17592 28648
rect 17644 28636 17650 28688
rect 3510 28568 3516 28620
rect 3568 28608 3574 28620
rect 9214 28608 9220 28620
rect 3568 28580 5396 28608
rect 9175 28580 9220 28608
rect 3568 28568 3574 28580
rect 1946 28540 1952 28552
rect 1907 28512 1952 28540
rect 1946 28500 1952 28512
rect 2004 28500 2010 28552
rect 4893 28543 4951 28549
rect 4893 28509 4905 28543
rect 4939 28540 4951 28543
rect 5074 28540 5080 28552
rect 4939 28512 5080 28540
rect 4939 28509 4951 28512
rect 4893 28503 4951 28509
rect 5074 28500 5080 28512
rect 5132 28500 5138 28552
rect 5368 28549 5396 28580
rect 9214 28568 9220 28580
rect 9272 28568 9278 28620
rect 12986 28568 12992 28620
rect 13044 28608 13050 28620
rect 14645 28611 14703 28617
rect 14645 28608 14657 28611
rect 13044 28580 14657 28608
rect 13044 28568 13050 28580
rect 14645 28577 14657 28580
rect 14691 28577 14703 28611
rect 14645 28571 14703 28577
rect 15654 28568 15660 28620
rect 15712 28608 15718 28620
rect 15749 28611 15807 28617
rect 15749 28608 15761 28611
rect 15712 28580 15761 28608
rect 15712 28568 15718 28580
rect 15749 28577 15761 28580
rect 15795 28577 15807 28611
rect 15749 28571 15807 28577
rect 15933 28611 15991 28617
rect 15933 28577 15945 28611
rect 15979 28608 15991 28611
rect 16022 28608 16028 28620
rect 15979 28580 16028 28608
rect 15979 28577 15991 28580
rect 15933 28571 15991 28577
rect 16022 28568 16028 28580
rect 16080 28568 16086 28620
rect 19613 28611 19671 28617
rect 19613 28577 19625 28611
rect 19659 28608 19671 28611
rect 24578 28608 24584 28620
rect 19659 28580 24584 28608
rect 19659 28577 19671 28580
rect 19613 28571 19671 28577
rect 24578 28568 24584 28580
rect 24636 28568 24642 28620
rect 5353 28543 5411 28549
rect 5353 28509 5365 28543
rect 5399 28509 5411 28543
rect 5353 28503 5411 28509
rect 9858 28500 9864 28552
rect 9916 28540 9922 28552
rect 10505 28543 10563 28549
rect 10505 28540 10517 28543
rect 9916 28512 10517 28540
rect 9916 28500 9922 28512
rect 10505 28509 10517 28512
rect 10551 28540 10563 28543
rect 10870 28540 10876 28552
rect 10551 28512 10876 28540
rect 10551 28509 10563 28512
rect 10505 28503 10563 28509
rect 10870 28500 10876 28512
rect 10928 28500 10934 28552
rect 14458 28540 14464 28552
rect 12406 28512 14464 28540
rect 8202 28432 8208 28484
rect 8260 28472 8266 28484
rect 9309 28475 9367 28481
rect 9309 28472 9321 28475
rect 8260 28444 9321 28472
rect 8260 28432 8266 28444
rect 9309 28441 9321 28444
rect 9355 28441 9367 28475
rect 9309 28435 9367 28441
rect 1765 28407 1823 28413
rect 1765 28373 1777 28407
rect 1811 28404 1823 28407
rect 1946 28404 1952 28416
rect 1811 28376 1952 28404
rect 1811 28373 1823 28376
rect 1765 28367 1823 28373
rect 1946 28364 1952 28376
rect 2004 28364 2010 28416
rect 4709 28407 4767 28413
rect 4709 28373 4721 28407
rect 4755 28404 4767 28407
rect 5350 28404 5356 28416
rect 4755 28376 5356 28404
rect 4755 28373 4767 28376
rect 4709 28367 4767 28373
rect 5350 28364 5356 28376
rect 5408 28364 5414 28416
rect 5442 28364 5448 28416
rect 5500 28404 5506 28416
rect 5500 28376 5545 28404
rect 5500 28364 5506 28376
rect 5626 28364 5632 28416
rect 5684 28404 5690 28416
rect 12406 28404 12434 28512
rect 14458 28500 14464 28512
rect 14516 28500 14522 28552
rect 15838 28500 15844 28552
rect 15896 28540 15902 28552
rect 17037 28543 17095 28549
rect 17037 28540 17049 28543
rect 15896 28512 17049 28540
rect 15896 28500 15902 28512
rect 17037 28509 17049 28512
rect 17083 28509 17095 28543
rect 17037 28503 17095 28509
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28509 19855 28543
rect 22002 28540 22008 28552
rect 21963 28512 22008 28540
rect 19797 28503 19855 28509
rect 14737 28475 14795 28481
rect 14737 28441 14749 28475
rect 14783 28472 14795 28475
rect 14826 28472 14832 28484
rect 14783 28444 14832 28472
rect 14783 28441 14795 28444
rect 14737 28435 14795 28441
rect 14826 28432 14832 28444
rect 14884 28432 14890 28484
rect 15289 28475 15347 28481
rect 15289 28441 15301 28475
rect 15335 28441 15347 28475
rect 15289 28435 15347 28441
rect 5684 28376 12434 28404
rect 15304 28404 15332 28435
rect 19426 28432 19432 28484
rect 19484 28472 19490 28484
rect 19812 28472 19840 28503
rect 22002 28500 22008 28512
rect 22060 28500 22066 28552
rect 24946 28540 24952 28552
rect 24907 28512 24952 28540
rect 24946 28500 24952 28512
rect 25004 28500 25010 28552
rect 19484 28444 19840 28472
rect 19484 28432 19490 28444
rect 15746 28404 15752 28416
rect 15304 28376 15752 28404
rect 5684 28364 5690 28376
rect 15746 28364 15752 28376
rect 15804 28364 15810 28416
rect 16393 28407 16451 28413
rect 16393 28373 16405 28407
rect 16439 28404 16451 28407
rect 19334 28404 19340 28416
rect 16439 28376 19340 28404
rect 16439 28373 16451 28376
rect 16393 28367 16451 28373
rect 19334 28364 19340 28376
rect 19392 28364 19398 28416
rect 20806 28364 20812 28416
rect 20864 28404 20870 28416
rect 21177 28407 21235 28413
rect 21177 28404 21189 28407
rect 20864 28376 21189 28404
rect 20864 28364 20870 28376
rect 21177 28373 21189 28376
rect 21223 28373 21235 28407
rect 21818 28404 21824 28416
rect 21779 28376 21824 28404
rect 21177 28367 21235 28373
rect 21818 28364 21824 28376
rect 21876 28364 21882 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 3050 28160 3056 28212
rect 3108 28200 3114 28212
rect 3108 28172 3740 28200
rect 3108 28160 3114 28172
rect 3142 28132 3148 28144
rect 3103 28104 3148 28132
rect 3142 28092 3148 28104
rect 3200 28092 3206 28144
rect 3712 28141 3740 28172
rect 5442 28160 5448 28212
rect 5500 28200 5506 28212
rect 14826 28200 14832 28212
rect 5500 28172 14412 28200
rect 14787 28172 14832 28200
rect 5500 28160 5506 28172
rect 3697 28135 3755 28141
rect 3697 28101 3709 28135
rect 3743 28101 3755 28135
rect 3697 28095 3755 28101
rect 3786 28092 3792 28144
rect 3844 28132 3850 28144
rect 4341 28135 4399 28141
rect 4341 28132 4353 28135
rect 3844 28104 4353 28132
rect 3844 28092 3850 28104
rect 4341 28101 4353 28104
rect 4387 28101 4399 28135
rect 4341 28095 4399 28101
rect 4893 28135 4951 28141
rect 4893 28101 4905 28135
rect 4939 28132 4951 28135
rect 9582 28132 9588 28144
rect 4939 28104 9588 28132
rect 4939 28101 4951 28104
rect 4893 28095 4951 28101
rect 9582 28092 9588 28104
rect 9640 28092 9646 28144
rect 13357 28135 13415 28141
rect 13357 28101 13369 28135
rect 13403 28132 13415 28135
rect 13906 28132 13912 28144
rect 13403 28104 13912 28132
rect 13403 28101 13415 28104
rect 13357 28095 13415 28101
rect 13906 28092 13912 28104
rect 13964 28092 13970 28144
rect 1578 28024 1584 28076
rect 1636 28064 1642 28076
rect 1857 28067 1915 28073
rect 1857 28064 1869 28067
rect 1636 28036 1869 28064
rect 1636 28024 1642 28036
rect 1857 28033 1869 28036
rect 1903 28033 1915 28067
rect 1857 28027 1915 28033
rect 5350 28024 5356 28076
rect 5408 28064 5414 28076
rect 5537 28067 5595 28073
rect 5537 28064 5549 28067
rect 5408 28036 5549 28064
rect 5408 28024 5414 28036
rect 5537 28033 5549 28036
rect 5583 28033 5595 28067
rect 14384 28064 14412 28172
rect 14826 28160 14832 28172
rect 14884 28160 14890 28212
rect 17497 28203 17555 28209
rect 17497 28169 17509 28203
rect 17543 28200 17555 28203
rect 19150 28200 19156 28212
rect 17543 28172 19156 28200
rect 17543 28169 17555 28172
rect 17497 28163 17555 28169
rect 19150 28160 19156 28172
rect 19208 28160 19214 28212
rect 19426 28200 19432 28212
rect 19387 28172 19432 28200
rect 19426 28160 19432 28172
rect 19484 28160 19490 28212
rect 21453 28203 21511 28209
rect 21453 28169 21465 28203
rect 21499 28200 21511 28203
rect 22738 28200 22744 28212
rect 21499 28172 22744 28200
rect 21499 28169 21511 28172
rect 21453 28163 21511 28169
rect 22738 28160 22744 28172
rect 22796 28160 22802 28212
rect 24026 28160 24032 28212
rect 24084 28200 24090 28212
rect 24305 28203 24363 28209
rect 24305 28200 24317 28203
rect 24084 28172 24317 28200
rect 24084 28160 24090 28172
rect 24305 28169 24317 28172
rect 24351 28169 24363 28203
rect 24305 28163 24363 28169
rect 24670 28160 24676 28212
rect 24728 28200 24734 28212
rect 25685 28203 25743 28209
rect 25685 28200 25697 28203
rect 24728 28172 25697 28200
rect 24728 28160 24734 28172
rect 25685 28169 25697 28172
rect 25731 28169 25743 28203
rect 25685 28163 25743 28169
rect 14458 28092 14464 28144
rect 14516 28132 14522 28144
rect 18233 28135 18291 28141
rect 14516 28104 16896 28132
rect 14516 28092 14522 28104
rect 15010 28064 15016 28076
rect 14384 28036 14872 28064
rect 14971 28036 15016 28064
rect 5537 28027 5595 28033
rect 3050 27996 3056 28008
rect 3011 27968 3056 27996
rect 3050 27956 3056 27968
rect 3108 27956 3114 28008
rect 3510 27956 3516 28008
rect 3568 27996 3574 28008
rect 4249 27999 4307 28005
rect 4249 27996 4261 27999
rect 3568 27968 4261 27996
rect 3568 27956 3574 27968
rect 4249 27965 4261 27968
rect 4295 27965 4307 27999
rect 4249 27959 4307 27965
rect 5810 27956 5816 28008
rect 5868 27996 5874 28008
rect 6549 27999 6607 28005
rect 6549 27996 6561 27999
rect 5868 27968 6561 27996
rect 5868 27956 5874 27968
rect 6549 27965 6561 27968
rect 6595 27965 6607 27999
rect 6549 27959 6607 27965
rect 13265 27999 13323 28005
rect 13265 27965 13277 27999
rect 13311 27996 13323 27999
rect 14366 27996 14372 28008
rect 13311 27968 14372 27996
rect 13311 27965 13323 27968
rect 13265 27959 13323 27965
rect 14366 27956 14372 27968
rect 14424 27956 14430 28008
rect 14844 27996 14872 28036
rect 15010 28024 15016 28036
rect 15068 28024 15074 28076
rect 15562 28024 15568 28076
rect 15620 28064 15626 28076
rect 15657 28067 15715 28073
rect 15657 28064 15669 28067
rect 15620 28036 15669 28064
rect 15620 28024 15626 28036
rect 15657 28033 15669 28036
rect 15703 28033 15715 28067
rect 15657 28027 15715 28033
rect 15838 28024 15844 28076
rect 15896 28064 15902 28076
rect 16868 28073 16896 28104
rect 18233 28101 18245 28135
rect 18279 28132 18291 28135
rect 20530 28132 20536 28144
rect 18279 28104 20536 28132
rect 18279 28101 18291 28104
rect 18233 28095 18291 28101
rect 20530 28092 20536 28104
rect 20588 28092 20594 28144
rect 29730 28132 29736 28144
rect 22020 28104 29736 28132
rect 16117 28067 16175 28073
rect 16117 28064 16129 28067
rect 15896 28036 16129 28064
rect 15896 28024 15902 28036
rect 16117 28033 16129 28036
rect 16163 28033 16175 28067
rect 16117 28027 16175 28033
rect 16853 28067 16911 28073
rect 16853 28033 16865 28067
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 17037 28067 17095 28073
rect 17037 28033 17049 28067
rect 17083 28064 17095 28067
rect 17126 28064 17132 28076
rect 17083 28036 17132 28064
rect 17083 28033 17095 28036
rect 17037 28027 17095 28033
rect 16758 27996 16764 28008
rect 14844 27968 16764 27996
rect 16758 27956 16764 27968
rect 16816 27956 16822 28008
rect 16868 27996 16896 28027
rect 17126 28024 17132 28036
rect 17184 28024 17190 28076
rect 19337 28067 19395 28073
rect 19337 28033 19349 28067
rect 19383 28064 19395 28067
rect 19426 28064 19432 28076
rect 19383 28036 19432 28064
rect 19383 28033 19395 28036
rect 19337 28027 19395 28033
rect 19426 28024 19432 28036
rect 19484 28064 19490 28076
rect 19978 28064 19984 28076
rect 19484 28036 19984 28064
rect 19484 28024 19490 28036
rect 19978 28024 19984 28036
rect 20036 28024 20042 28076
rect 20806 28064 20812 28076
rect 20767 28036 20812 28064
rect 20806 28024 20812 28036
rect 20864 28024 20870 28076
rect 20993 28067 21051 28073
rect 20993 28033 21005 28067
rect 21039 28064 21051 28067
rect 21818 28064 21824 28076
rect 21039 28036 21824 28064
rect 21039 28033 21051 28036
rect 20993 28027 21051 28033
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 22020 28073 22048 28104
rect 29730 28092 29736 28104
rect 29788 28092 29794 28144
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28033 22063 28067
rect 23014 28064 23020 28076
rect 22975 28036 23020 28064
rect 22005 28027 22063 28033
rect 23014 28024 23020 28036
rect 23072 28024 23078 28076
rect 25038 28064 25044 28076
rect 24999 28036 25044 28064
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 18138 27996 18144 28008
rect 16868 27968 17172 27996
rect 18099 27968 18144 27996
rect 13817 27931 13875 27937
rect 13817 27897 13829 27931
rect 13863 27897 13875 27931
rect 13817 27891 13875 27897
rect 15473 27931 15531 27937
rect 15473 27897 15485 27931
rect 15519 27928 15531 27931
rect 17034 27928 17040 27940
rect 15519 27900 17040 27928
rect 15519 27897 15531 27900
rect 15473 27891 15531 27897
rect 1949 27863 2007 27869
rect 1949 27829 1961 27863
rect 1995 27860 2007 27863
rect 3326 27860 3332 27872
rect 1995 27832 3332 27860
rect 1995 27829 2007 27832
rect 1949 27823 2007 27829
rect 3326 27820 3332 27832
rect 3384 27820 3390 27872
rect 5353 27863 5411 27869
rect 5353 27829 5365 27863
rect 5399 27860 5411 27863
rect 5902 27860 5908 27872
rect 5399 27832 5908 27860
rect 5399 27829 5411 27832
rect 5353 27823 5411 27829
rect 5902 27820 5908 27832
rect 5960 27820 5966 27872
rect 13832 27860 13860 27891
rect 17034 27888 17040 27900
rect 17092 27888 17098 27940
rect 17144 27928 17172 27968
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 18417 27999 18475 28005
rect 18417 27965 18429 27999
rect 18463 27965 18475 27999
rect 18417 27959 18475 27965
rect 23661 27999 23719 28005
rect 23661 27965 23673 27999
rect 23707 27965 23719 27999
rect 23842 27996 23848 28008
rect 23803 27968 23848 27996
rect 23661 27959 23719 27965
rect 18432 27928 18460 27959
rect 17144 27900 18460 27928
rect 23676 27928 23704 27959
rect 23842 27956 23848 27968
rect 23900 27956 23906 28008
rect 25222 27996 25228 28008
rect 25183 27968 25228 27996
rect 25222 27956 25228 27968
rect 25280 27956 25286 28008
rect 27154 27928 27160 27940
rect 23676 27900 27160 27928
rect 27154 27888 27160 27900
rect 27212 27888 27218 27940
rect 15746 27860 15752 27872
rect 13832 27832 15752 27860
rect 15746 27820 15752 27832
rect 15804 27820 15810 27872
rect 16209 27863 16267 27869
rect 16209 27829 16221 27863
rect 16255 27860 16267 27863
rect 17402 27860 17408 27872
rect 16255 27832 17408 27860
rect 16255 27829 16267 27832
rect 16209 27823 16267 27829
rect 17402 27820 17408 27832
rect 17460 27820 17466 27872
rect 20806 27820 20812 27872
rect 20864 27860 20870 27872
rect 22097 27863 22155 27869
rect 22097 27860 22109 27863
rect 20864 27832 22109 27860
rect 20864 27820 20870 27832
rect 22097 27829 22109 27832
rect 22143 27829 22155 27863
rect 22097 27823 22155 27829
rect 22833 27863 22891 27869
rect 22833 27829 22845 27863
rect 22879 27860 22891 27863
rect 23566 27860 23572 27872
rect 22879 27832 23572 27860
rect 22879 27829 22891 27832
rect 22833 27823 22891 27829
rect 23566 27820 23572 27832
rect 23624 27820 23630 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 11228 27659 11286 27665
rect 11228 27625 11240 27659
rect 11274 27656 11286 27659
rect 13722 27656 13728 27668
rect 11274 27628 13728 27656
rect 11274 27625 11286 27628
rect 11228 27619 11286 27625
rect 13722 27616 13728 27628
rect 13780 27616 13786 27668
rect 19426 27656 19432 27668
rect 13832 27628 19432 27656
rect 1581 27591 1639 27597
rect 1581 27557 1593 27591
rect 1627 27588 1639 27591
rect 3970 27588 3976 27600
rect 1627 27560 3976 27588
rect 1627 27557 1639 27560
rect 1581 27551 1639 27557
rect 3970 27548 3976 27560
rect 4028 27548 4034 27600
rect 12713 27591 12771 27597
rect 12713 27557 12725 27591
rect 12759 27588 12771 27591
rect 13832 27588 13860 27628
rect 19426 27616 19432 27628
rect 19484 27616 19490 27668
rect 21361 27659 21419 27665
rect 21361 27625 21373 27659
rect 21407 27656 21419 27659
rect 22002 27656 22008 27668
rect 21407 27628 22008 27656
rect 21407 27625 21419 27628
rect 21361 27619 21419 27625
rect 22002 27616 22008 27628
rect 22060 27616 22066 27668
rect 23934 27616 23940 27668
rect 23992 27656 23998 27668
rect 24578 27656 24584 27668
rect 23992 27628 24584 27656
rect 23992 27616 23998 27628
rect 24578 27616 24584 27628
rect 24636 27656 24642 27668
rect 24673 27659 24731 27665
rect 24673 27656 24685 27659
rect 24636 27628 24685 27656
rect 24636 27616 24642 27628
rect 24673 27625 24685 27628
rect 24719 27625 24731 27659
rect 24673 27619 24731 27625
rect 25222 27616 25228 27668
rect 25280 27656 25286 27668
rect 25317 27659 25375 27665
rect 25317 27656 25329 27659
rect 25280 27628 25329 27656
rect 25280 27616 25286 27628
rect 25317 27625 25329 27628
rect 25363 27625 25375 27659
rect 25317 27619 25375 27625
rect 12759 27560 13860 27588
rect 12759 27557 12771 27560
rect 12713 27551 12771 27557
rect 4709 27523 4767 27529
rect 4709 27489 4721 27523
rect 4755 27520 4767 27523
rect 5626 27520 5632 27532
rect 4755 27492 5632 27520
rect 4755 27489 4767 27492
rect 4709 27483 4767 27489
rect 5626 27480 5632 27492
rect 5684 27480 5690 27532
rect 5810 27520 5816 27532
rect 5771 27492 5816 27520
rect 5810 27480 5816 27492
rect 5868 27480 5874 27532
rect 12728 27520 12756 27551
rect 19334 27548 19340 27600
rect 19392 27588 19398 27600
rect 19797 27591 19855 27597
rect 19797 27588 19809 27591
rect 19392 27560 19809 27588
rect 19392 27548 19398 27560
rect 19797 27557 19809 27560
rect 19843 27588 19855 27591
rect 19978 27588 19984 27600
rect 19843 27560 19984 27588
rect 19843 27557 19855 27560
rect 19797 27551 19855 27557
rect 19978 27548 19984 27560
rect 20036 27548 20042 27600
rect 20530 27588 20536 27600
rect 20491 27560 20536 27588
rect 20530 27548 20536 27560
rect 20588 27548 20594 27600
rect 23385 27591 23443 27597
rect 23385 27557 23397 27591
rect 23431 27588 23443 27591
rect 23842 27588 23848 27600
rect 23431 27560 23848 27588
rect 23431 27557 23443 27560
rect 23385 27551 23443 27557
rect 23842 27548 23848 27560
rect 23900 27548 23906 27600
rect 30374 27588 30380 27600
rect 24596 27560 30380 27588
rect 12544 27492 12756 27520
rect 1762 27452 1768 27464
rect 1723 27424 1768 27452
rect 1762 27412 1768 27424
rect 1820 27412 1826 27464
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 10965 27455 11023 27461
rect 10965 27452 10977 27455
rect 9180 27424 10977 27452
rect 9180 27412 9186 27424
rect 10965 27421 10977 27424
rect 11011 27421 11023 27455
rect 10965 27415 11023 27421
rect 4062 27384 4068 27396
rect 4023 27356 4068 27384
rect 4062 27344 4068 27356
rect 4120 27344 4126 27396
rect 4157 27387 4215 27393
rect 4157 27353 4169 27387
rect 4203 27384 4215 27387
rect 4338 27384 4344 27396
rect 4203 27356 4344 27384
rect 4203 27353 4215 27356
rect 4157 27347 4215 27353
rect 4338 27344 4344 27356
rect 4396 27344 4402 27396
rect 5902 27344 5908 27396
rect 5960 27384 5966 27396
rect 5960 27356 6005 27384
rect 5960 27344 5966 27356
rect 6178 27344 6184 27396
rect 6236 27384 6242 27396
rect 6454 27384 6460 27396
rect 6236 27356 6460 27384
rect 6236 27344 6242 27356
rect 6454 27344 6460 27356
rect 6512 27344 6518 27396
rect 11882 27344 11888 27396
rect 11940 27344 11946 27396
rect 4246 27276 4252 27328
rect 4304 27316 4310 27328
rect 12158 27316 12164 27328
rect 4304 27288 12164 27316
rect 4304 27276 4310 27288
rect 12158 27276 12164 27288
rect 12216 27316 12222 27328
rect 12544 27316 12572 27492
rect 14642 27480 14648 27532
rect 14700 27520 14706 27532
rect 14700 27492 17172 27520
rect 14700 27480 14706 27492
rect 16393 27455 16451 27461
rect 16393 27421 16405 27455
rect 16439 27452 16451 27455
rect 16482 27452 16488 27464
rect 16439 27424 16488 27452
rect 16439 27421 16451 27424
rect 16393 27415 16451 27421
rect 16482 27412 16488 27424
rect 16540 27412 16546 27464
rect 17034 27452 17040 27464
rect 16995 27424 17040 27452
rect 17034 27412 17040 27424
rect 17092 27412 17098 27464
rect 17144 27452 17172 27492
rect 17402 27480 17408 27532
rect 17460 27520 17466 27532
rect 17460 27492 18000 27520
rect 17460 27480 17466 27492
rect 17497 27455 17555 27461
rect 17497 27452 17509 27455
rect 17144 27424 17509 27452
rect 17497 27421 17509 27424
rect 17543 27421 17555 27455
rect 17972 27452 18000 27492
rect 18138 27480 18144 27532
rect 18196 27520 18202 27532
rect 18233 27523 18291 27529
rect 18233 27520 18245 27523
rect 18196 27492 18245 27520
rect 18196 27480 18202 27492
rect 18233 27489 18245 27492
rect 18279 27489 18291 27523
rect 18233 27483 18291 27489
rect 19429 27523 19487 27529
rect 19429 27489 19441 27523
rect 19475 27520 19487 27523
rect 20806 27520 20812 27532
rect 19475 27492 20812 27520
rect 19475 27489 19487 27492
rect 19429 27483 19487 27489
rect 20806 27480 20812 27492
rect 20864 27480 20870 27532
rect 19613 27455 19671 27461
rect 19613 27452 19625 27455
rect 17972 27424 19625 27452
rect 17497 27415 17555 27421
rect 19613 27421 19625 27424
rect 19659 27421 19671 27455
rect 20714 27452 20720 27464
rect 20675 27424 20720 27452
rect 19613 27415 19671 27421
rect 20714 27412 20720 27424
rect 20772 27412 20778 27464
rect 21174 27412 21180 27464
rect 21232 27452 21238 27464
rect 21545 27455 21603 27461
rect 21545 27452 21557 27455
rect 21232 27424 21557 27452
rect 21232 27412 21238 27424
rect 21545 27421 21557 27424
rect 21591 27421 21603 27455
rect 23566 27452 23572 27464
rect 23527 27424 23572 27452
rect 21545 27415 21603 27421
rect 23566 27412 23572 27424
rect 23624 27412 23630 27464
rect 24596 27461 24624 27560
rect 30374 27548 30380 27560
rect 30432 27548 30438 27600
rect 26528 27492 35894 27520
rect 24581 27455 24639 27461
rect 24581 27421 24593 27455
rect 24627 27421 24639 27455
rect 25222 27452 25228 27464
rect 25183 27424 25228 27452
rect 24581 27415 24639 27421
rect 25222 27412 25228 27424
rect 25280 27412 25286 27464
rect 26528 27461 26556 27492
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27421 26111 27455
rect 26053 27415 26111 27421
rect 26513 27455 26571 27461
rect 26513 27421 26525 27455
rect 26559 27421 26571 27455
rect 27430 27452 27436 27464
rect 27391 27424 27436 27452
rect 26513 27415 26571 27421
rect 14918 27344 14924 27396
rect 14976 27384 14982 27396
rect 17589 27387 17647 27393
rect 17589 27384 17601 27387
rect 14976 27356 17601 27384
rect 14976 27344 14982 27356
rect 17589 27353 17601 27356
rect 17635 27353 17647 27387
rect 26068 27384 26096 27415
rect 27430 27412 27436 27424
rect 27488 27412 27494 27464
rect 35866 27452 35894 27492
rect 37734 27452 37740 27464
rect 35866 27424 37740 27452
rect 37734 27412 37740 27424
rect 37792 27412 37798 27464
rect 17589 27347 17647 27353
rect 24596 27356 26096 27384
rect 24596 27328 24624 27356
rect 26234 27344 26240 27396
rect 26292 27384 26298 27396
rect 27525 27387 27583 27393
rect 27525 27384 27537 27387
rect 26292 27356 27537 27384
rect 26292 27344 26298 27356
rect 27525 27353 27537 27356
rect 27571 27353 27583 27387
rect 27525 27347 27583 27353
rect 12216 27288 12572 27316
rect 12216 27276 12222 27288
rect 12802 27276 12808 27328
rect 12860 27316 12866 27328
rect 13998 27316 14004 27328
rect 12860 27288 14004 27316
rect 12860 27276 12866 27288
rect 13998 27276 14004 27288
rect 14056 27276 14062 27328
rect 16206 27316 16212 27328
rect 16167 27288 16212 27316
rect 16206 27276 16212 27288
rect 16264 27276 16270 27328
rect 16850 27316 16856 27328
rect 16811 27288 16856 27316
rect 16850 27276 16856 27288
rect 16908 27276 16914 27328
rect 24578 27276 24584 27328
rect 24636 27276 24642 27328
rect 24762 27276 24768 27328
rect 24820 27316 24826 27328
rect 25869 27319 25927 27325
rect 25869 27316 25881 27319
rect 24820 27288 25881 27316
rect 24820 27276 24826 27288
rect 25869 27285 25881 27288
rect 25915 27285 25927 27319
rect 25869 27279 25927 27285
rect 26605 27319 26663 27325
rect 26605 27285 26617 27319
rect 26651 27316 26663 27319
rect 27246 27316 27252 27328
rect 26651 27288 27252 27316
rect 26651 27285 26663 27288
rect 26605 27279 26663 27285
rect 27246 27276 27252 27288
rect 27304 27276 27310 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 4338 27112 4344 27124
rect 4299 27084 4344 27112
rect 4338 27072 4344 27084
rect 4396 27072 4402 27124
rect 12710 27112 12716 27124
rect 8312 27084 12716 27112
rect 6638 27004 6644 27056
rect 6696 27044 6702 27056
rect 8312 27053 8340 27084
rect 12710 27072 12716 27084
rect 12768 27072 12774 27124
rect 14550 27112 14556 27124
rect 12912 27084 14556 27112
rect 8297 27047 8355 27053
rect 8297 27044 8309 27047
rect 6696 27016 8309 27044
rect 6696 27004 6702 27016
rect 8297 27013 8309 27016
rect 8343 27013 8355 27047
rect 10962 27044 10968 27056
rect 9522 27016 10968 27044
rect 8297 27007 8355 27013
rect 10962 27004 10968 27016
rect 11020 27004 11026 27056
rect 11146 27004 11152 27056
rect 11204 27044 11210 27056
rect 11977 27047 12035 27053
rect 11977 27044 11989 27047
rect 11204 27016 11989 27044
rect 11204 27004 11210 27016
rect 11977 27013 11989 27016
rect 12023 27013 12035 27047
rect 12526 27044 12532 27056
rect 12487 27016 12532 27044
rect 11977 27007 12035 27013
rect 12526 27004 12532 27016
rect 12584 27004 12590 27056
rect 1670 26936 1676 26988
rect 1728 26976 1734 26988
rect 1857 26979 1915 26985
rect 1857 26976 1869 26979
rect 1728 26948 1869 26976
rect 1728 26936 1734 26948
rect 1857 26945 1869 26948
rect 1903 26945 1915 26979
rect 4246 26976 4252 26988
rect 4207 26948 4252 26976
rect 1857 26939 1915 26945
rect 4246 26936 4252 26948
rect 4304 26936 4310 26988
rect 12802 26976 12808 26988
rect 12544 26948 12808 26976
rect 8021 26911 8079 26917
rect 8021 26877 8033 26911
rect 8067 26908 8079 26911
rect 10042 26908 10048 26920
rect 8067 26880 8156 26908
rect 10003 26880 10048 26908
rect 8067 26877 8079 26880
rect 8021 26871 8079 26877
rect 1854 26772 1860 26784
rect 1815 26744 1860 26772
rect 1854 26732 1860 26744
rect 1912 26732 1918 26784
rect 8128 26772 8156 26880
rect 10042 26868 10048 26880
rect 10100 26868 10106 26920
rect 11885 26911 11943 26917
rect 11885 26877 11897 26911
rect 11931 26908 11943 26911
rect 12544 26908 12572 26948
rect 12802 26936 12808 26948
rect 12860 26936 12866 26988
rect 11931 26880 12572 26908
rect 11931 26877 11943 26880
rect 11885 26871 11943 26877
rect 9306 26800 9312 26852
rect 9364 26840 9370 26852
rect 12912 26840 12940 27084
rect 14550 27072 14556 27084
rect 14608 27072 14614 27124
rect 19337 27115 19395 27121
rect 19337 27081 19349 27115
rect 19383 27112 19395 27115
rect 20714 27112 20720 27124
rect 19383 27084 20720 27112
rect 19383 27081 19395 27084
rect 19337 27075 19395 27081
rect 20714 27072 20720 27084
rect 20772 27072 20778 27124
rect 22554 27072 22560 27124
rect 22612 27112 22618 27124
rect 25222 27112 25228 27124
rect 22612 27084 25228 27112
rect 22612 27072 22618 27084
rect 25222 27072 25228 27084
rect 25280 27072 25286 27124
rect 15930 27044 15936 27056
rect 14490 27016 15936 27044
rect 15930 27004 15936 27016
rect 15988 27004 15994 27056
rect 22922 27044 22928 27056
rect 19306 27016 22928 27044
rect 16117 26979 16175 26985
rect 16117 26945 16129 26979
rect 16163 26976 16175 26979
rect 16390 26976 16396 26988
rect 16163 26948 16396 26976
rect 16163 26945 16175 26948
rect 16117 26939 16175 26945
rect 16390 26936 16396 26948
rect 16448 26936 16454 26988
rect 19306 26976 19334 27016
rect 22922 27004 22928 27016
rect 22980 27004 22986 27056
rect 24762 27044 24768 27056
rect 24723 27016 24768 27044
rect 24762 27004 24768 27016
rect 24820 27004 24826 27056
rect 16500 26948 19334 26976
rect 12986 26868 12992 26920
rect 13044 26908 13050 26920
rect 13262 26908 13268 26920
rect 13044 26880 13089 26908
rect 13223 26880 13268 26908
rect 13044 26868 13050 26880
rect 13262 26868 13268 26880
rect 13320 26868 13326 26920
rect 13722 26868 13728 26920
rect 13780 26908 13786 26920
rect 13780 26880 14320 26908
rect 13780 26868 13786 26880
rect 9364 26812 12940 26840
rect 14292 26840 14320 26880
rect 14550 26868 14556 26920
rect 14608 26908 14614 26920
rect 16500 26908 16528 26948
rect 19426 26936 19432 26988
rect 19484 26976 19490 26988
rect 19521 26979 19579 26985
rect 19521 26976 19533 26979
rect 19484 26948 19533 26976
rect 19484 26936 19490 26948
rect 19521 26945 19533 26948
rect 19567 26945 19579 26979
rect 20254 26976 20260 26988
rect 20215 26948 20260 26976
rect 19521 26939 19579 26945
rect 20254 26936 20260 26948
rect 20312 26936 20318 26988
rect 20993 26979 21051 26985
rect 20993 26945 21005 26979
rect 21039 26976 21051 26979
rect 21082 26976 21088 26988
rect 21039 26948 21088 26976
rect 21039 26945 21051 26948
rect 20993 26939 21051 26945
rect 21082 26936 21088 26948
rect 21140 26936 21146 26988
rect 27525 26979 27583 26985
rect 27525 26945 27537 26979
rect 27571 26976 27583 26979
rect 37274 26976 37280 26988
rect 27571 26948 37280 26976
rect 27571 26945 27583 26948
rect 27525 26939 27583 26945
rect 37274 26936 37280 26948
rect 37332 26936 37338 26988
rect 38286 26976 38292 26988
rect 38247 26948 38292 26976
rect 38286 26936 38292 26948
rect 38344 26936 38350 26988
rect 17310 26908 17316 26920
rect 14608 26880 16528 26908
rect 17271 26880 17316 26908
rect 14608 26868 14614 26880
rect 17310 26868 17316 26880
rect 17368 26868 17374 26920
rect 17402 26868 17408 26920
rect 17460 26908 17466 26920
rect 20714 26908 20720 26920
rect 17460 26880 20720 26908
rect 17460 26868 17466 26880
rect 20714 26868 20720 26880
rect 20772 26868 20778 26920
rect 24486 26908 24492 26920
rect 22066 26880 24492 26908
rect 16114 26840 16120 26852
rect 14292 26812 16120 26840
rect 9364 26800 9370 26812
rect 16114 26800 16120 26812
rect 16172 26840 16178 26852
rect 22066 26840 22094 26880
rect 24486 26868 24492 26880
rect 24544 26868 24550 26920
rect 24670 26908 24676 26920
rect 24631 26880 24676 26908
rect 24670 26868 24676 26880
rect 24728 26868 24734 26920
rect 24949 26911 25007 26917
rect 24949 26877 24961 26911
rect 24995 26877 25007 26911
rect 24949 26871 25007 26877
rect 16172 26812 22094 26840
rect 16172 26800 16178 26812
rect 24118 26800 24124 26852
rect 24176 26840 24182 26852
rect 24964 26840 24992 26871
rect 31754 26840 31760 26852
rect 24176 26812 31760 26840
rect 24176 26800 24182 26812
rect 31754 26800 31760 26812
rect 31812 26800 31818 26852
rect 8294 26772 8300 26784
rect 8128 26744 8300 26772
rect 8294 26732 8300 26744
rect 8352 26732 8358 26784
rect 10778 26732 10784 26784
rect 10836 26772 10842 26784
rect 13814 26772 13820 26784
rect 10836 26744 13820 26772
rect 10836 26732 10842 26744
rect 13814 26732 13820 26744
rect 13872 26732 13878 26784
rect 14734 26772 14740 26784
rect 14695 26744 14740 26772
rect 14734 26732 14740 26744
rect 14792 26732 14798 26784
rect 14826 26732 14832 26784
rect 14884 26772 14890 26784
rect 16209 26775 16267 26781
rect 16209 26772 16221 26775
rect 14884 26744 16221 26772
rect 14884 26732 14890 26744
rect 16209 26741 16221 26744
rect 16255 26741 16267 26775
rect 16209 26735 16267 26741
rect 19610 26732 19616 26784
rect 19668 26772 19674 26784
rect 20073 26775 20131 26781
rect 20073 26772 20085 26775
rect 19668 26744 20085 26772
rect 19668 26732 19674 26744
rect 20073 26741 20085 26744
rect 20119 26741 20131 26775
rect 20073 26735 20131 26741
rect 20806 26732 20812 26784
rect 20864 26772 20870 26784
rect 21085 26775 21143 26781
rect 21085 26772 21097 26775
rect 20864 26744 21097 26772
rect 20864 26732 20870 26744
rect 21085 26741 21097 26744
rect 21131 26741 21143 26775
rect 21085 26735 21143 26741
rect 25958 26732 25964 26784
rect 26016 26772 26022 26784
rect 27617 26775 27675 26781
rect 27617 26772 27629 26775
rect 26016 26744 27629 26772
rect 26016 26732 26022 26744
rect 27617 26741 27629 26744
rect 27663 26741 27675 26775
rect 27617 26735 27675 26741
rect 37274 26732 37280 26784
rect 37332 26772 37338 26784
rect 38105 26775 38163 26781
rect 38105 26772 38117 26775
rect 37332 26744 38117 26772
rect 37332 26732 37338 26744
rect 38105 26741 38117 26744
rect 38151 26741 38163 26775
rect 38105 26735 38163 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 2501 26571 2559 26577
rect 2501 26537 2513 26571
rect 2547 26568 2559 26571
rect 3050 26568 3056 26580
rect 2547 26540 3056 26568
rect 2547 26537 2559 26540
rect 2501 26531 2559 26537
rect 3050 26528 3056 26540
rect 3108 26528 3114 26580
rect 5629 26571 5687 26577
rect 5629 26537 5641 26571
rect 5675 26568 5687 26571
rect 6168 26571 6226 26577
rect 6168 26568 6180 26571
rect 5675 26540 6180 26568
rect 5675 26537 5687 26540
rect 5629 26531 5687 26537
rect 6168 26537 6180 26540
rect 6214 26568 6226 26571
rect 26237 26571 26295 26577
rect 6214 26540 24716 26568
rect 6214 26537 6226 26540
rect 6168 26531 6226 26537
rect 16482 26500 16488 26512
rect 16443 26472 16488 26500
rect 16482 26460 16488 26472
rect 16540 26460 16546 26512
rect 18690 26500 18696 26512
rect 16684 26472 18696 26500
rect 1854 26432 1860 26444
rect 1815 26404 1860 26432
rect 1854 26392 1860 26404
rect 1912 26392 1918 26444
rect 2041 26435 2099 26441
rect 2041 26401 2053 26435
rect 2087 26432 2099 26435
rect 2498 26432 2504 26444
rect 2087 26404 2504 26432
rect 2087 26401 2099 26404
rect 2041 26395 2099 26401
rect 2498 26392 2504 26404
rect 2556 26392 2562 26444
rect 5905 26435 5963 26441
rect 5905 26401 5917 26435
rect 5951 26432 5963 26435
rect 8294 26432 8300 26444
rect 5951 26404 8300 26432
rect 5951 26401 5963 26404
rect 5905 26395 5963 26401
rect 8294 26392 8300 26404
rect 8352 26432 8358 26444
rect 9122 26432 9128 26444
rect 8352 26404 9128 26432
rect 8352 26392 8358 26404
rect 9122 26392 9128 26404
rect 9180 26432 9186 26444
rect 9401 26435 9459 26441
rect 9401 26432 9413 26435
rect 9180 26404 9413 26432
rect 9180 26392 9186 26404
rect 9401 26401 9413 26404
rect 9447 26432 9459 26435
rect 11885 26435 11943 26441
rect 11885 26432 11897 26435
rect 9447 26404 11897 26432
rect 9447 26401 9459 26404
rect 9401 26395 9459 26401
rect 11885 26401 11897 26404
rect 11931 26432 11943 26435
rect 13170 26432 13176 26444
rect 11931 26404 13176 26432
rect 11931 26401 11943 26404
rect 11885 26395 11943 26401
rect 13170 26392 13176 26404
rect 13228 26432 13234 26444
rect 14277 26435 14335 26441
rect 14277 26432 14289 26435
rect 13228 26404 14289 26432
rect 13228 26392 13234 26404
rect 14277 26401 14289 26404
rect 14323 26401 14335 26435
rect 14550 26432 14556 26444
rect 14511 26404 14556 26432
rect 14277 26395 14335 26401
rect 14550 26392 14556 26404
rect 14608 26392 14614 26444
rect 3142 26364 3148 26376
rect 3103 26336 3148 26364
rect 3142 26324 3148 26336
rect 3200 26324 3206 26376
rect 7929 26367 7987 26373
rect 7929 26333 7941 26367
rect 7975 26364 7987 26367
rect 9306 26364 9312 26376
rect 7975 26336 9312 26364
rect 7975 26333 7987 26336
rect 7929 26327 7987 26333
rect 9306 26324 9312 26336
rect 9364 26324 9370 26376
rect 10778 26324 10784 26376
rect 10836 26324 10842 26376
rect 16574 26364 16580 26376
rect 10980 26336 11928 26364
rect 9677 26299 9735 26305
rect 7406 26268 9628 26296
rect 2958 26228 2964 26240
rect 2919 26200 2964 26228
rect 2958 26188 2964 26200
rect 3016 26188 3022 26240
rect 9600 26228 9628 26268
rect 9677 26265 9689 26299
rect 9723 26296 9735 26299
rect 9723 26268 10088 26296
rect 9723 26265 9735 26268
rect 9677 26259 9735 26265
rect 9766 26228 9772 26240
rect 9600 26200 9772 26228
rect 9766 26188 9772 26200
rect 9824 26188 9830 26240
rect 10060 26228 10088 26268
rect 10980 26228 11008 26336
rect 11422 26296 11428 26308
rect 11383 26268 11428 26296
rect 11422 26256 11428 26268
rect 11480 26256 11486 26308
rect 11900 26296 11928 26336
rect 15856 26336 16580 26364
rect 11900 26268 12112 26296
rect 10060 26200 11008 26228
rect 12084 26228 12112 26268
rect 12158 26256 12164 26308
rect 12216 26296 12222 26308
rect 12216 26268 12261 26296
rect 12216 26256 12222 26268
rect 12894 26256 12900 26308
rect 12952 26256 12958 26308
rect 13648 26268 14964 26296
rect 13648 26237 13676 26268
rect 13633 26231 13691 26237
rect 13633 26228 13645 26231
rect 12084 26200 13645 26228
rect 13633 26197 13645 26200
rect 13679 26197 13691 26231
rect 14936 26228 14964 26268
rect 15010 26256 15016 26308
rect 15068 26256 15074 26308
rect 15856 26228 15884 26336
rect 16574 26324 16580 26336
rect 16632 26324 16638 26376
rect 16684 26373 16712 26472
rect 18690 26460 18696 26472
rect 18748 26460 18754 26512
rect 19426 26460 19432 26512
rect 19484 26500 19490 26512
rect 20073 26503 20131 26509
rect 20073 26500 20085 26503
rect 19484 26472 20085 26500
rect 19484 26460 19490 26472
rect 20073 26469 20085 26472
rect 20119 26469 20131 26503
rect 20073 26463 20131 26469
rect 22557 26503 22615 26509
rect 22557 26469 22569 26503
rect 22603 26500 22615 26503
rect 22738 26500 22744 26512
rect 22603 26472 22744 26500
rect 22603 26469 22615 26472
rect 22557 26463 22615 26469
rect 22738 26460 22744 26472
rect 22796 26460 22802 26512
rect 24578 26500 24584 26512
rect 24539 26472 24584 26500
rect 24578 26460 24584 26472
rect 24636 26460 24642 26512
rect 24688 26500 24716 26540
rect 26237 26537 26249 26571
rect 26283 26568 26295 26571
rect 27798 26568 27804 26580
rect 26283 26540 27804 26568
rect 26283 26537 26295 26540
rect 26237 26531 26295 26537
rect 27798 26528 27804 26540
rect 27856 26528 27862 26580
rect 24688 26472 35894 26500
rect 17310 26432 17316 26444
rect 17271 26404 17316 26432
rect 17310 26392 17316 26404
rect 17368 26392 17374 26444
rect 17586 26432 17592 26444
rect 17547 26404 17592 26432
rect 17586 26392 17592 26404
rect 17644 26392 17650 26444
rect 19521 26435 19579 26441
rect 19521 26401 19533 26435
rect 19567 26432 19579 26435
rect 19567 26404 20576 26432
rect 19567 26401 19579 26404
rect 19521 26395 19579 26401
rect 16669 26367 16727 26373
rect 16669 26333 16681 26367
rect 16715 26333 16727 26367
rect 16669 26327 16727 26333
rect 16114 26296 16120 26308
rect 16040 26268 16120 26296
rect 16040 26237 16068 26268
rect 16114 26256 16120 26268
rect 16172 26256 16178 26308
rect 16206 26256 16212 26308
rect 16264 26296 16270 26308
rect 17405 26299 17463 26305
rect 17405 26296 17417 26299
rect 16264 26268 17417 26296
rect 16264 26256 16270 26268
rect 17405 26265 17417 26268
rect 17451 26265 17463 26299
rect 17405 26259 17463 26265
rect 19610 26256 19616 26308
rect 19668 26296 19674 26308
rect 20548 26296 20576 26404
rect 20622 26392 20628 26444
rect 20680 26432 20686 26444
rect 20806 26432 20812 26444
rect 20680 26404 20725 26432
rect 20767 26404 20812 26432
rect 20680 26392 20686 26404
rect 20806 26392 20812 26404
rect 20864 26392 20870 26444
rect 27890 26432 27896 26444
rect 27851 26404 27896 26432
rect 27890 26392 27896 26404
rect 27948 26392 27954 26444
rect 28077 26435 28135 26441
rect 28077 26401 28089 26435
rect 28123 26432 28135 26435
rect 29089 26435 29147 26441
rect 29089 26432 29101 26435
rect 28123 26404 29101 26432
rect 28123 26401 28135 26404
rect 28077 26395 28135 26401
rect 29089 26401 29101 26404
rect 29135 26401 29147 26435
rect 35866 26432 35894 26472
rect 37366 26432 37372 26444
rect 35866 26404 37372 26432
rect 29089 26395 29147 26401
rect 37366 26392 37372 26404
rect 37424 26392 37430 26444
rect 21266 26364 21272 26376
rect 21227 26336 21272 26364
rect 21266 26324 21272 26336
rect 21324 26364 21330 26376
rect 21913 26367 21971 26373
rect 21913 26364 21925 26367
rect 21324 26336 21925 26364
rect 21324 26324 21330 26336
rect 21913 26333 21925 26336
rect 21959 26333 21971 26367
rect 22094 26364 22100 26376
rect 22055 26336 22100 26364
rect 21913 26327 21971 26333
rect 22094 26324 22100 26336
rect 22152 26324 22158 26376
rect 22278 26324 22284 26376
rect 22336 26364 22342 26376
rect 24765 26367 24823 26373
rect 24765 26364 24777 26367
rect 22336 26336 24777 26364
rect 22336 26324 22342 26336
rect 24765 26333 24777 26336
rect 24811 26333 24823 26367
rect 26421 26367 26479 26373
rect 26421 26364 26433 26367
rect 24765 26327 24823 26333
rect 26206 26336 26433 26364
rect 22186 26296 22192 26308
rect 19668 26268 19713 26296
rect 20548 26268 22192 26296
rect 19668 26256 19674 26268
rect 22186 26256 22192 26268
rect 22244 26256 22250 26308
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 26206 26296 26234 26336
rect 26421 26333 26433 26336
rect 26467 26333 26479 26367
rect 26421 26327 26479 26333
rect 27338 26324 27344 26376
rect 27396 26364 27402 26376
rect 28997 26367 29055 26373
rect 28997 26364 29009 26367
rect 27396 26336 29009 26364
rect 27396 26324 27402 26336
rect 28997 26333 29009 26336
rect 29043 26333 29055 26367
rect 28997 26327 29055 26333
rect 24544 26268 26234 26296
rect 24544 26256 24550 26268
rect 14936 26200 15884 26228
rect 16025 26231 16083 26237
rect 13633 26191 13691 26197
rect 16025 26197 16037 26231
rect 16071 26197 16083 26231
rect 16025 26191 16083 26197
rect 27614 26188 27620 26240
rect 27672 26228 27678 26240
rect 28537 26231 28595 26237
rect 28537 26228 28549 26231
rect 27672 26200 28549 26228
rect 27672 26188 27678 26200
rect 28537 26197 28549 26200
rect 28583 26197 28595 26231
rect 28537 26191 28595 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 2501 26027 2559 26033
rect 2501 25993 2513 26027
rect 2547 26024 2559 26027
rect 3050 26024 3056 26036
rect 2547 25996 3056 26024
rect 2547 25993 2559 25996
rect 2501 25987 2559 25993
rect 3050 25984 3056 25996
rect 3108 25984 3114 26036
rect 5258 26024 5264 26036
rect 3344 25996 5264 26024
rect 2041 25891 2099 25897
rect 2041 25857 2053 25891
rect 2087 25888 2099 25891
rect 2406 25888 2412 25900
rect 2087 25860 2412 25888
rect 2087 25857 2099 25860
rect 2041 25851 2099 25857
rect 2406 25848 2412 25860
rect 2464 25848 2470 25900
rect 3344 25897 3372 25996
rect 5258 25984 5264 25996
rect 5316 26024 5322 26036
rect 5316 25996 5580 26024
rect 5316 25984 5322 25996
rect 3329 25891 3387 25897
rect 3329 25857 3341 25891
rect 3375 25857 3387 25891
rect 3329 25851 3387 25857
rect 5350 25848 5356 25900
rect 5408 25848 5414 25900
rect 5552 25888 5580 25996
rect 9030 25984 9036 26036
rect 9088 26024 9094 26036
rect 11422 26024 11428 26036
rect 9088 25996 11428 26024
rect 9088 25984 9094 25996
rect 11422 25984 11428 25996
rect 11480 26024 11486 26036
rect 12342 26024 12348 26036
rect 11480 25996 12348 26024
rect 11480 25984 11486 25996
rect 12342 25984 12348 25996
rect 12400 25984 12406 26036
rect 13265 26027 13323 26033
rect 13265 25993 13277 26027
rect 13311 26024 13323 26027
rect 15010 26024 15016 26036
rect 13311 25996 15016 26024
rect 13311 25993 13323 25996
rect 13265 25987 13323 25993
rect 15010 25984 15016 25996
rect 15068 25984 15074 26036
rect 21361 26027 21419 26033
rect 21361 25993 21373 26027
rect 21407 26024 21419 26027
rect 22094 26024 22100 26036
rect 21407 25996 22100 26024
rect 21407 25993 21419 25996
rect 21361 25987 21419 25993
rect 22094 25984 22100 25996
rect 22152 25984 22158 26036
rect 8202 25916 8208 25968
rect 8260 25956 8266 25968
rect 14366 25956 14372 25968
rect 8260 25928 14372 25956
rect 8260 25916 8266 25928
rect 14366 25916 14372 25928
rect 14424 25956 14430 25968
rect 14642 25956 14648 25968
rect 14424 25928 14648 25956
rect 14424 25916 14430 25928
rect 14642 25916 14648 25928
rect 14700 25916 14706 25968
rect 16850 25916 16856 25968
rect 16908 25956 16914 25968
rect 17773 25959 17831 25965
rect 17773 25956 17785 25959
rect 16908 25928 17785 25956
rect 16908 25916 16914 25928
rect 17773 25925 17785 25928
rect 17819 25925 17831 25959
rect 19334 25956 19340 25968
rect 19295 25928 19340 25956
rect 17773 25919 17831 25925
rect 19334 25916 19340 25928
rect 19392 25916 19398 25968
rect 28534 25956 28540 25968
rect 27172 25928 28540 25956
rect 27172 25900 27200 25928
rect 28534 25916 28540 25928
rect 28592 25956 28598 25968
rect 28905 25959 28963 25965
rect 28905 25956 28917 25959
rect 28592 25928 28917 25956
rect 28592 25916 28598 25928
rect 28905 25925 28917 25928
rect 28951 25925 28963 25959
rect 28905 25919 28963 25925
rect 10042 25888 10048 25900
rect 5552 25860 10048 25888
rect 10042 25848 10048 25860
rect 10100 25848 10106 25900
rect 13173 25891 13231 25897
rect 13173 25857 13185 25891
rect 13219 25888 13231 25891
rect 16206 25888 16212 25900
rect 13219 25860 16212 25888
rect 13219 25857 13231 25860
rect 13173 25851 13231 25857
rect 1854 25820 1860 25832
rect 1815 25792 1860 25820
rect 1854 25780 1860 25792
rect 1912 25820 1918 25832
rect 2222 25820 2228 25832
rect 1912 25792 2228 25820
rect 1912 25780 1918 25792
rect 2222 25780 2228 25792
rect 2280 25780 2286 25832
rect 3970 25820 3976 25832
rect 3931 25792 3976 25820
rect 3970 25780 3976 25792
rect 4028 25780 4034 25832
rect 4249 25823 4307 25829
rect 4249 25789 4261 25823
rect 4295 25820 4307 25823
rect 10594 25820 10600 25832
rect 4295 25792 10600 25820
rect 4295 25789 4307 25792
rect 4249 25783 4307 25789
rect 10594 25780 10600 25792
rect 10652 25780 10658 25832
rect 11698 25780 11704 25832
rect 11756 25820 11762 25832
rect 13188 25820 13216 25851
rect 16206 25848 16212 25860
rect 16264 25888 16270 25900
rect 16390 25888 16396 25900
rect 16264 25860 16396 25888
rect 16264 25848 16270 25860
rect 16390 25848 16396 25860
rect 16448 25888 16454 25900
rect 16945 25891 17003 25897
rect 16945 25888 16957 25891
rect 16448 25860 16957 25888
rect 16448 25848 16454 25860
rect 16945 25857 16957 25860
rect 16991 25857 17003 25891
rect 16945 25851 17003 25857
rect 20714 25848 20720 25900
rect 20772 25888 20778 25900
rect 20809 25891 20867 25897
rect 20809 25888 20821 25891
rect 20772 25860 20821 25888
rect 20772 25848 20778 25860
rect 20809 25857 20821 25860
rect 20855 25857 20867 25891
rect 20809 25851 20867 25857
rect 21174 25848 21180 25900
rect 21232 25888 21238 25900
rect 21269 25891 21327 25897
rect 21269 25888 21281 25891
rect 21232 25860 21281 25888
rect 21232 25848 21238 25860
rect 21269 25857 21281 25860
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 22370 25848 22376 25900
rect 22428 25888 22434 25900
rect 23293 25891 23351 25897
rect 23293 25888 23305 25891
rect 22428 25860 23305 25888
rect 22428 25848 22434 25860
rect 23293 25857 23305 25860
rect 23339 25857 23351 25891
rect 23293 25851 23351 25857
rect 26605 25891 26663 25897
rect 26605 25857 26617 25891
rect 26651 25888 26663 25891
rect 27062 25888 27068 25900
rect 26651 25860 27068 25888
rect 26651 25857 26663 25860
rect 26605 25851 26663 25857
rect 27062 25848 27068 25860
rect 27120 25848 27126 25900
rect 27154 25848 27160 25900
rect 27212 25888 27218 25900
rect 28813 25891 28871 25897
rect 27212 25860 27257 25888
rect 27212 25848 27218 25860
rect 28813 25857 28825 25891
rect 28859 25857 28871 25891
rect 29454 25888 29460 25900
rect 29415 25860 29460 25888
rect 28813 25851 28871 25857
rect 17681 25823 17739 25829
rect 17681 25820 17693 25823
rect 11756 25792 13216 25820
rect 17604 25792 17693 25820
rect 11756 25780 11762 25792
rect 17604 25764 17632 25792
rect 17681 25789 17693 25792
rect 17727 25789 17739 25823
rect 18506 25820 18512 25832
rect 18467 25792 18512 25820
rect 17681 25783 17739 25789
rect 18506 25780 18512 25792
rect 18564 25780 18570 25832
rect 19242 25820 19248 25832
rect 19203 25792 19248 25820
rect 19242 25780 19248 25792
rect 19300 25780 19306 25832
rect 19518 25820 19524 25832
rect 19479 25792 19524 25820
rect 19518 25780 19524 25792
rect 19576 25780 19582 25832
rect 27341 25823 27399 25829
rect 27341 25789 27353 25823
rect 27387 25789 27399 25823
rect 28828 25820 28856 25851
rect 29454 25848 29460 25860
rect 29512 25848 29518 25900
rect 38102 25820 38108 25832
rect 28828 25792 38108 25820
rect 27341 25783 27399 25789
rect 17586 25712 17592 25764
rect 17644 25712 17650 25764
rect 26421 25755 26479 25761
rect 26421 25721 26433 25755
rect 26467 25752 26479 25755
rect 27356 25752 27384 25783
rect 38102 25780 38108 25792
rect 38160 25780 38166 25832
rect 26467 25724 27384 25752
rect 26467 25721 26479 25724
rect 26421 25715 26479 25721
rect 3418 25684 3424 25696
rect 3379 25656 3424 25684
rect 3418 25644 3424 25656
rect 3476 25644 3482 25696
rect 5721 25687 5779 25693
rect 5721 25653 5733 25687
rect 5767 25684 5779 25687
rect 11146 25684 11152 25696
rect 5767 25656 11152 25684
rect 5767 25653 5779 25656
rect 5721 25647 5779 25653
rect 11146 25644 11152 25656
rect 11204 25644 11210 25696
rect 16022 25644 16028 25696
rect 16080 25684 16086 25696
rect 17037 25687 17095 25693
rect 17037 25684 17049 25687
rect 16080 25656 17049 25684
rect 16080 25644 16086 25656
rect 17037 25653 17049 25656
rect 17083 25653 17095 25687
rect 20622 25684 20628 25696
rect 20583 25656 20628 25684
rect 17037 25647 17095 25653
rect 20622 25644 20628 25656
rect 20680 25644 20686 25696
rect 23109 25687 23167 25693
rect 23109 25653 23121 25687
rect 23155 25684 23167 25687
rect 23474 25684 23480 25696
rect 23155 25656 23480 25684
rect 23155 25653 23167 25656
rect 23109 25647 23167 25653
rect 23474 25644 23480 25656
rect 23532 25644 23538 25696
rect 27614 25684 27620 25696
rect 27575 25656 27620 25684
rect 27614 25644 27620 25656
rect 27672 25644 27678 25696
rect 28166 25644 28172 25696
rect 28224 25684 28230 25696
rect 29549 25687 29607 25693
rect 29549 25684 29561 25687
rect 28224 25656 29561 25684
rect 28224 25644 28230 25656
rect 29549 25653 29561 25656
rect 29595 25653 29607 25687
rect 29549 25647 29607 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 3329 25483 3387 25489
rect 3329 25449 3341 25483
rect 3375 25480 3387 25483
rect 3786 25480 3792 25492
rect 3375 25452 3792 25480
rect 3375 25449 3387 25452
rect 3329 25443 3387 25449
rect 3786 25440 3792 25452
rect 3844 25440 3850 25492
rect 5350 25440 5356 25492
rect 5408 25480 5414 25492
rect 13722 25480 13728 25492
rect 5408 25452 13728 25480
rect 5408 25440 5414 25452
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 19981 25483 20039 25489
rect 19981 25449 19993 25483
rect 20027 25480 20039 25483
rect 20254 25480 20260 25492
rect 20027 25452 20260 25480
rect 20027 25449 20039 25452
rect 19981 25443 20039 25449
rect 20254 25440 20260 25452
rect 20312 25440 20318 25492
rect 22370 25480 22376 25492
rect 22331 25452 22376 25480
rect 22370 25440 22376 25452
rect 22428 25440 22434 25492
rect 27062 25480 27068 25492
rect 27023 25452 27068 25480
rect 27062 25440 27068 25452
rect 27120 25440 27126 25492
rect 32953 25483 33011 25489
rect 32953 25449 32965 25483
rect 32999 25480 33011 25483
rect 36630 25480 36636 25492
rect 32999 25452 36636 25480
rect 32999 25449 33011 25452
rect 32953 25443 33011 25449
rect 36630 25440 36636 25452
rect 36688 25440 36694 25492
rect 38102 25480 38108 25492
rect 38063 25452 38108 25480
rect 38102 25440 38108 25452
rect 38160 25440 38166 25492
rect 2041 25415 2099 25421
rect 2041 25381 2053 25415
rect 2087 25412 2099 25415
rect 3510 25412 3516 25424
rect 2087 25384 3516 25412
rect 2087 25381 2099 25384
rect 2041 25375 2099 25381
rect 3510 25372 3516 25384
rect 3568 25372 3574 25424
rect 4617 25415 4675 25421
rect 4617 25381 4629 25415
rect 4663 25412 4675 25415
rect 4663 25384 9260 25412
rect 4663 25381 4675 25384
rect 4617 25375 4675 25381
rect 2958 25344 2964 25356
rect 1964 25316 2964 25344
rect 1964 25285 1992 25316
rect 2958 25304 2964 25316
rect 3016 25304 3022 25356
rect 3326 25304 3332 25356
rect 3384 25344 3390 25356
rect 4065 25347 4123 25353
rect 4065 25344 4077 25347
rect 3384 25316 4077 25344
rect 3384 25304 3390 25316
rect 4065 25313 4077 25316
rect 4111 25313 4123 25347
rect 9122 25344 9128 25356
rect 9083 25316 9128 25344
rect 4065 25307 4123 25313
rect 9122 25304 9128 25316
rect 9180 25304 9186 25356
rect 9232 25344 9260 25384
rect 10962 25372 10968 25424
rect 11020 25412 11026 25424
rect 16393 25415 16451 25421
rect 16393 25412 16405 25415
rect 11020 25384 16405 25412
rect 11020 25372 11026 25384
rect 16393 25381 16405 25384
rect 16439 25381 16451 25415
rect 19518 25412 19524 25424
rect 16393 25375 16451 25381
rect 18340 25384 19524 25412
rect 18340 25344 18368 25384
rect 19518 25372 19524 25384
rect 19576 25372 19582 25424
rect 9232 25316 18368 25344
rect 18417 25347 18475 25353
rect 18417 25313 18429 25347
rect 18463 25344 18475 25347
rect 19242 25344 19248 25356
rect 18463 25316 19248 25344
rect 18463 25313 18475 25316
rect 18417 25307 18475 25313
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 23385 25347 23443 25353
rect 23385 25313 23397 25347
rect 23431 25344 23443 25347
rect 26234 25344 26240 25356
rect 23431 25316 26240 25344
rect 23431 25313 23443 25316
rect 23385 25307 23443 25313
rect 26234 25304 26240 25316
rect 26292 25304 26298 25356
rect 28534 25344 28540 25356
rect 28495 25316 28540 25344
rect 28534 25304 28540 25316
rect 28592 25304 28598 25356
rect 1949 25279 2007 25285
rect 1949 25245 1961 25279
rect 1995 25245 2007 25279
rect 1949 25239 2007 25245
rect 2498 25236 2504 25288
rect 2556 25276 2562 25288
rect 2593 25279 2651 25285
rect 2593 25276 2605 25279
rect 2556 25248 2605 25276
rect 2556 25236 2562 25248
rect 2593 25245 2605 25248
rect 2639 25245 2651 25279
rect 2593 25239 2651 25245
rect 3237 25279 3295 25285
rect 3237 25245 3249 25279
rect 3283 25245 3295 25279
rect 3237 25239 3295 25245
rect 3252 25208 3280 25239
rect 8202 25236 8208 25288
rect 8260 25276 8266 25288
rect 8389 25279 8447 25285
rect 8389 25276 8401 25279
rect 8260 25248 8401 25276
rect 8260 25236 8266 25248
rect 8389 25245 8401 25248
rect 8435 25245 8447 25279
rect 8389 25239 8447 25245
rect 16301 25279 16359 25285
rect 16301 25245 16313 25279
rect 16347 25276 16359 25279
rect 16390 25276 16396 25288
rect 16347 25248 16396 25276
rect 16347 25245 16359 25248
rect 16301 25239 16359 25245
rect 16390 25236 16396 25248
rect 16448 25236 16454 25288
rect 20165 25279 20223 25285
rect 20165 25245 20177 25279
rect 20211 25276 20223 25279
rect 20530 25276 20536 25288
rect 20211 25248 20536 25276
rect 20211 25245 20223 25248
rect 20165 25239 20223 25245
rect 20530 25236 20536 25248
rect 20588 25236 20594 25288
rect 20898 25276 20904 25288
rect 20859 25248 20904 25276
rect 20898 25236 20904 25248
rect 20956 25236 20962 25288
rect 22557 25279 22615 25285
rect 22557 25245 22569 25279
rect 22603 25276 22615 25279
rect 22922 25276 22928 25288
rect 22603 25248 22928 25276
rect 22603 25245 22615 25248
rect 22557 25239 22615 25245
rect 22922 25236 22928 25248
rect 22980 25236 22986 25288
rect 23566 25276 23572 25288
rect 23527 25248 23572 25276
rect 23566 25236 23572 25248
rect 23624 25236 23630 25288
rect 24486 25236 24492 25288
rect 24544 25276 24550 25288
rect 24581 25279 24639 25285
rect 24581 25276 24593 25279
rect 24544 25248 24593 25276
rect 24544 25236 24550 25248
rect 24581 25245 24593 25248
rect 24627 25245 24639 25279
rect 24581 25239 24639 25245
rect 27154 25236 27160 25288
rect 27212 25276 27218 25288
rect 27249 25279 27307 25285
rect 27249 25276 27261 25279
rect 27212 25248 27261 25276
rect 27212 25236 27218 25248
rect 27249 25245 27261 25248
rect 27295 25276 27307 25279
rect 27338 25276 27344 25288
rect 27295 25248 27344 25276
rect 27295 25245 27307 25248
rect 27249 25239 27307 25245
rect 27338 25236 27344 25248
rect 27396 25236 27402 25288
rect 27798 25236 27804 25288
rect 27856 25276 27862 25288
rect 27893 25279 27951 25285
rect 27893 25276 27905 25279
rect 27856 25248 27905 25276
rect 27856 25236 27862 25248
rect 27893 25245 27905 25248
rect 27939 25245 27951 25279
rect 27893 25239 27951 25245
rect 28721 25279 28779 25285
rect 28721 25245 28733 25279
rect 28767 25276 28779 25279
rect 28994 25276 29000 25288
rect 28767 25248 29000 25276
rect 28767 25245 28779 25248
rect 28721 25239 28779 25245
rect 28994 25236 29000 25248
rect 29052 25236 29058 25288
rect 32309 25279 32367 25285
rect 32309 25245 32321 25279
rect 32355 25245 32367 25279
rect 32309 25239 32367 25245
rect 32401 25279 32459 25285
rect 32401 25245 32413 25279
rect 32447 25276 32459 25279
rect 33137 25279 33195 25285
rect 33137 25276 33149 25279
rect 32447 25248 33149 25276
rect 32447 25245 32459 25248
rect 32401 25239 32459 25245
rect 33137 25245 33149 25248
rect 33183 25245 33195 25279
rect 38286 25276 38292 25288
rect 38247 25248 38292 25276
rect 33137 25239 33195 25245
rect 3326 25208 3332 25220
rect 3252 25180 3332 25208
rect 3326 25168 3332 25180
rect 3384 25208 3390 25220
rect 3694 25208 3700 25220
rect 3384 25180 3700 25208
rect 3384 25168 3390 25180
rect 3694 25168 3700 25180
rect 3752 25168 3758 25220
rect 4157 25211 4215 25217
rect 4157 25177 4169 25211
rect 4203 25177 4215 25211
rect 4157 25171 4215 25177
rect 2682 25140 2688 25152
rect 2643 25112 2688 25140
rect 2682 25100 2688 25112
rect 2740 25100 2746 25152
rect 3418 25100 3424 25152
rect 3476 25140 3482 25152
rect 4172 25140 4200 25171
rect 9030 25168 9036 25220
rect 9088 25208 9094 25220
rect 9401 25211 9459 25217
rect 9401 25208 9413 25211
rect 9088 25180 9413 25208
rect 9088 25168 9094 25180
rect 9401 25177 9413 25180
rect 9447 25177 9459 25211
rect 14826 25208 14832 25220
rect 10626 25180 14832 25208
rect 9401 25171 9459 25177
rect 14826 25168 14832 25180
rect 14884 25168 14890 25220
rect 28902 25168 28908 25220
rect 28960 25208 28966 25220
rect 32324 25208 32352 25239
rect 38286 25236 38292 25248
rect 38344 25236 38350 25288
rect 28960 25180 32352 25208
rect 28960 25168 28966 25180
rect 3476 25112 4200 25140
rect 3476 25100 3482 25112
rect 5442 25100 5448 25152
rect 5500 25140 5506 25152
rect 8481 25143 8539 25149
rect 8481 25140 8493 25143
rect 5500 25112 8493 25140
rect 5500 25100 5506 25112
rect 8481 25109 8493 25112
rect 8527 25109 8539 25143
rect 10870 25140 10876 25152
rect 10831 25112 10876 25140
rect 8481 25103 8539 25109
rect 10870 25100 10876 25112
rect 10928 25100 10934 25152
rect 20717 25143 20775 25149
rect 20717 25109 20729 25143
rect 20763 25140 20775 25143
rect 20990 25140 20996 25152
rect 20763 25112 20996 25140
rect 20763 25109 20775 25112
rect 20717 25103 20775 25109
rect 20990 25100 20996 25112
rect 21048 25100 21054 25152
rect 24026 25140 24032 25152
rect 23987 25112 24032 25140
rect 24026 25100 24032 25112
rect 24084 25100 24090 25152
rect 24673 25143 24731 25149
rect 24673 25109 24685 25143
rect 24719 25140 24731 25143
rect 25314 25140 25320 25152
rect 24719 25112 25320 25140
rect 24719 25109 24731 25112
rect 24673 25103 24731 25109
rect 25314 25100 25320 25112
rect 25372 25100 25378 25152
rect 27706 25140 27712 25152
rect 27667 25112 27712 25140
rect 27706 25100 27712 25112
rect 27764 25100 27770 25152
rect 29181 25143 29239 25149
rect 29181 25109 29193 25143
rect 29227 25140 29239 25143
rect 29822 25140 29828 25152
rect 29227 25112 29828 25140
rect 29227 25109 29239 25112
rect 29181 25103 29239 25109
rect 29822 25100 29828 25112
rect 29880 25100 29886 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19705 24939 19763 24945
rect 19705 24936 19717 24939
rect 19392 24908 19717 24936
rect 19392 24896 19398 24908
rect 19705 24905 19717 24908
rect 19751 24905 19763 24939
rect 19705 24899 19763 24905
rect 23937 24939 23995 24945
rect 23937 24905 23949 24939
rect 23983 24936 23995 24939
rect 24026 24936 24032 24948
rect 23983 24908 24032 24936
rect 23983 24905 23995 24908
rect 23937 24899 23995 24905
rect 24026 24896 24032 24908
rect 24084 24896 24090 24948
rect 17218 24868 17224 24880
rect 17179 24840 17224 24868
rect 17218 24828 17224 24840
rect 17276 24828 17282 24880
rect 25314 24868 25320 24880
rect 25275 24840 25320 24868
rect 25314 24828 25320 24840
rect 25372 24828 25378 24880
rect 30285 24871 30343 24877
rect 30285 24868 30297 24871
rect 30024 24840 30297 24868
rect 7558 24800 7564 24812
rect 3174 24772 7564 24800
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 10873 24803 10931 24809
rect 10873 24769 10885 24803
rect 10919 24800 10931 24803
rect 11698 24800 11704 24812
rect 10919 24772 11704 24800
rect 10919 24769 10931 24772
rect 10873 24763 10931 24769
rect 11698 24760 11704 24772
rect 11756 24760 11762 24812
rect 16022 24800 16028 24812
rect 14858 24772 16028 24800
rect 16022 24760 16028 24772
rect 16080 24760 16086 24812
rect 16114 24760 16120 24812
rect 16172 24800 16178 24812
rect 19889 24803 19947 24809
rect 16172 24772 16217 24800
rect 16172 24760 16178 24772
rect 19889 24769 19901 24803
rect 19935 24800 19947 24803
rect 20622 24800 20628 24812
rect 19935 24772 20628 24800
rect 19935 24769 19947 24772
rect 19889 24763 19947 24769
rect 20622 24760 20628 24772
rect 20680 24760 20686 24812
rect 20990 24800 20996 24812
rect 20951 24772 20996 24800
rect 20990 24760 20996 24772
rect 21048 24760 21054 24812
rect 22649 24803 22707 24809
rect 22649 24769 22661 24803
rect 22695 24800 22707 24803
rect 22922 24800 22928 24812
rect 22695 24772 22928 24800
rect 22695 24769 22707 24772
rect 22649 24763 22707 24769
rect 22922 24760 22928 24772
rect 22980 24760 22986 24812
rect 23474 24800 23480 24812
rect 23435 24772 23480 24800
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 25869 24803 25927 24809
rect 25869 24769 25881 24803
rect 25915 24800 25927 24803
rect 27982 24800 27988 24812
rect 25915 24772 27988 24800
rect 25915 24769 25927 24772
rect 25869 24763 25927 24769
rect 27982 24760 27988 24772
rect 28040 24760 28046 24812
rect 28350 24760 28356 24812
rect 28408 24800 28414 24812
rect 28537 24803 28595 24809
rect 28537 24800 28549 24803
rect 28408 24772 28549 24800
rect 28408 24760 28414 24772
rect 28537 24769 28549 24772
rect 28583 24769 28595 24803
rect 28537 24763 28595 24769
rect 28626 24760 28632 24812
rect 28684 24800 28690 24812
rect 28997 24803 29055 24809
rect 28997 24800 29009 24803
rect 28684 24772 29009 24800
rect 28684 24760 28690 24772
rect 28997 24769 29009 24772
rect 29043 24769 29055 24803
rect 28997 24763 29055 24769
rect 29089 24803 29147 24809
rect 29089 24769 29101 24803
rect 29135 24800 29147 24803
rect 30024 24800 30052 24840
rect 30285 24837 30297 24840
rect 30331 24837 30343 24871
rect 30285 24831 30343 24837
rect 29135 24772 30052 24800
rect 29135 24769 29147 24772
rect 29089 24763 29147 24769
rect 1765 24735 1823 24741
rect 1765 24701 1777 24735
rect 1811 24732 1823 24735
rect 2041 24735 2099 24741
rect 1811 24704 1900 24732
rect 1811 24701 1823 24704
rect 1765 24695 1823 24701
rect 1872 24596 1900 24704
rect 2041 24701 2053 24735
rect 2087 24732 2099 24735
rect 2590 24732 2596 24744
rect 2087 24704 2596 24732
rect 2087 24701 2099 24704
rect 2041 24695 2099 24701
rect 2590 24692 2596 24704
rect 2648 24692 2654 24744
rect 9766 24692 9772 24744
rect 9824 24732 9830 24744
rect 10965 24735 11023 24741
rect 10965 24732 10977 24735
rect 9824 24704 10977 24732
rect 9824 24692 9830 24704
rect 10965 24701 10977 24704
rect 11011 24701 11023 24735
rect 10965 24695 11023 24701
rect 13170 24692 13176 24744
rect 13228 24732 13234 24744
rect 13449 24735 13507 24741
rect 13449 24732 13461 24735
rect 13228 24704 13461 24732
rect 13228 24692 13234 24704
rect 13449 24701 13461 24704
rect 13495 24701 13507 24735
rect 13725 24735 13783 24741
rect 13725 24732 13737 24735
rect 13449 24695 13507 24701
rect 13556 24704 13737 24732
rect 12986 24624 12992 24676
rect 13044 24664 13050 24676
rect 13556 24664 13584 24704
rect 13725 24701 13737 24704
rect 13771 24701 13783 24735
rect 13725 24695 13783 24701
rect 15930 24692 15936 24744
rect 15988 24732 15994 24744
rect 16209 24735 16267 24741
rect 16209 24732 16221 24735
rect 15988 24704 16221 24732
rect 15988 24692 15994 24704
rect 16209 24701 16221 24704
rect 16255 24701 16267 24735
rect 17129 24735 17187 24741
rect 17129 24732 17141 24735
rect 16209 24695 16267 24701
rect 16316 24704 17141 24732
rect 13044 24636 13584 24664
rect 13044 24624 13050 24636
rect 15654 24624 15660 24676
rect 15712 24664 15718 24676
rect 16316 24664 16344 24704
rect 17129 24701 17141 24704
rect 17175 24701 17187 24735
rect 17129 24695 17187 24701
rect 17405 24735 17463 24741
rect 17405 24701 17417 24735
rect 17451 24701 17463 24735
rect 17405 24695 17463 24701
rect 23293 24735 23351 24741
rect 23293 24701 23305 24735
rect 23339 24732 23351 24735
rect 23382 24732 23388 24744
rect 23339 24704 23388 24732
rect 23339 24701 23351 24704
rect 23293 24695 23351 24701
rect 15712 24636 16344 24664
rect 15712 24624 15718 24636
rect 17034 24624 17040 24676
rect 17092 24664 17098 24676
rect 17420 24664 17448 24695
rect 23382 24692 23388 24704
rect 23440 24732 23446 24744
rect 23934 24732 23940 24744
rect 23440 24704 23940 24732
rect 23440 24692 23446 24704
rect 23934 24692 23940 24704
rect 23992 24692 23998 24744
rect 24026 24692 24032 24744
rect 24084 24732 24090 24744
rect 25225 24735 25283 24741
rect 25225 24732 25237 24735
rect 24084 24704 25237 24732
rect 24084 24692 24090 24704
rect 25225 24701 25237 24704
rect 25271 24701 25283 24735
rect 25225 24695 25283 24701
rect 29546 24692 29552 24744
rect 29604 24732 29610 24744
rect 30193 24735 30251 24741
rect 30193 24732 30205 24735
rect 29604 24704 30205 24732
rect 29604 24692 29610 24704
rect 30193 24701 30205 24704
rect 30239 24701 30251 24735
rect 30466 24732 30472 24744
rect 30427 24704 30472 24732
rect 30193 24695 30251 24701
rect 30466 24692 30472 24704
rect 30524 24692 30530 24744
rect 17092 24636 17448 24664
rect 22741 24667 22799 24673
rect 17092 24624 17098 24636
rect 22741 24633 22753 24667
rect 22787 24664 22799 24667
rect 23566 24664 23572 24676
rect 22787 24636 23572 24664
rect 22787 24633 22799 24636
rect 22741 24627 22799 24633
rect 23566 24624 23572 24636
rect 23624 24624 23630 24676
rect 2774 24596 2780 24608
rect 1872 24568 2780 24596
rect 2774 24556 2780 24568
rect 2832 24556 2838 24608
rect 3510 24596 3516 24608
rect 3471 24568 3516 24596
rect 3510 24556 3516 24568
rect 3568 24556 3574 24608
rect 15197 24599 15255 24605
rect 15197 24565 15209 24599
rect 15243 24596 15255 24599
rect 15930 24596 15936 24608
rect 15243 24568 15936 24596
rect 15243 24565 15255 24568
rect 15197 24559 15255 24565
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 20806 24596 20812 24608
rect 20767 24568 20812 24596
rect 20806 24556 20812 24568
rect 20864 24556 20870 24608
rect 28353 24599 28411 24605
rect 28353 24565 28365 24599
rect 28399 24596 28411 24599
rect 29914 24596 29920 24608
rect 28399 24568 29920 24596
rect 28399 24565 28411 24568
rect 28353 24559 28411 24565
rect 29914 24556 29920 24568
rect 29972 24556 29978 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1762 24392 1768 24404
rect 1723 24364 1768 24392
rect 1762 24352 1768 24364
rect 1820 24352 1826 24404
rect 4062 24392 4068 24404
rect 4023 24364 4068 24392
rect 4062 24352 4068 24364
rect 4120 24352 4126 24404
rect 5902 24352 5908 24404
rect 5960 24392 5966 24404
rect 13630 24392 13636 24404
rect 5960 24364 13636 24392
rect 5960 24352 5966 24364
rect 13630 24352 13636 24364
rect 13688 24352 13694 24404
rect 13722 24352 13728 24404
rect 13780 24392 13786 24404
rect 15841 24395 15899 24401
rect 15841 24392 15853 24395
rect 13780 24364 15853 24392
rect 13780 24352 13786 24364
rect 15841 24361 15853 24364
rect 15887 24361 15899 24395
rect 15841 24355 15899 24361
rect 15930 24352 15936 24404
rect 15988 24392 15994 24404
rect 22278 24392 22284 24404
rect 15988 24364 22284 24392
rect 15988 24352 15994 24364
rect 22278 24352 22284 24364
rect 22336 24352 22342 24404
rect 28994 24392 29000 24404
rect 27448 24364 27752 24392
rect 28955 24364 29000 24392
rect 6638 24324 6644 24336
rect 6599 24296 6644 24324
rect 6638 24284 6644 24296
rect 6696 24284 6702 24336
rect 1854 24216 1860 24268
rect 1912 24256 1918 24268
rect 20346 24256 20352 24268
rect 1912 24228 20352 24256
rect 1912 24216 1918 24228
rect 20346 24216 20352 24228
rect 20404 24216 20410 24268
rect 20806 24256 20812 24268
rect 20767 24228 20812 24256
rect 20806 24216 20812 24228
rect 20864 24216 20870 24268
rect 20898 24216 20904 24268
rect 20956 24256 20962 24268
rect 21542 24256 21548 24268
rect 20956 24228 21548 24256
rect 20956 24216 20962 24228
rect 21542 24216 21548 24228
rect 21600 24256 21606 24268
rect 21600 24228 23152 24256
rect 21600 24216 21606 24228
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24188 1639 24191
rect 1946 24188 1952 24200
rect 1627 24160 1952 24188
rect 1627 24157 1639 24160
rect 1581 24151 1639 24157
rect 1946 24148 1952 24160
rect 2004 24148 2010 24200
rect 2866 24148 2872 24200
rect 2924 24188 2930 24200
rect 3973 24191 4031 24197
rect 3973 24188 3985 24191
rect 2924 24160 3985 24188
rect 2924 24148 2930 24160
rect 3973 24157 3985 24160
rect 4019 24157 4031 24191
rect 3973 24151 4031 24157
rect 4062 24148 4068 24200
rect 4120 24188 4126 24200
rect 4893 24191 4951 24197
rect 4893 24188 4905 24191
rect 4120 24160 4905 24188
rect 4120 24148 4126 24160
rect 4893 24157 4905 24160
rect 4939 24157 4951 24191
rect 4893 24151 4951 24157
rect 7742 24148 7748 24200
rect 7800 24188 7806 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 7800 24160 9137 24188
rect 7800 24148 7806 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9125 24151 9183 24157
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24188 14611 24191
rect 15286 24188 15292 24200
rect 14599 24160 15292 24188
rect 14599 24157 14611 24160
rect 14553 24151 14611 24157
rect 15286 24148 15292 24160
rect 15344 24188 15350 24200
rect 15749 24191 15807 24197
rect 15749 24188 15761 24191
rect 15344 24160 15761 24188
rect 15344 24148 15350 24160
rect 15749 24157 15761 24160
rect 15795 24188 15807 24191
rect 16114 24188 16120 24200
rect 15795 24160 16120 24188
rect 15795 24157 15807 24160
rect 15749 24151 15807 24157
rect 16114 24148 16120 24160
rect 16172 24148 16178 24200
rect 16390 24188 16396 24200
rect 16351 24160 16396 24188
rect 16390 24148 16396 24160
rect 16448 24148 16454 24200
rect 18690 24188 18696 24200
rect 18651 24160 18696 24188
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 23124 24197 23152 24228
rect 20625 24191 20683 24197
rect 20625 24157 20637 24191
rect 20671 24157 20683 24191
rect 20625 24151 20683 24157
rect 23109 24191 23167 24197
rect 23109 24157 23121 24191
rect 23155 24157 23167 24191
rect 25406 24188 25412 24200
rect 25367 24160 25412 24188
rect 23109 24151 23167 24157
rect 5169 24123 5227 24129
rect 5169 24089 5181 24123
rect 5215 24089 5227 24123
rect 16485 24123 16543 24129
rect 16485 24120 16497 24123
rect 6394 24092 16497 24120
rect 5169 24083 5227 24089
rect 16485 24089 16497 24092
rect 16531 24089 16543 24123
rect 16485 24083 16543 24089
rect 5184 24052 5212 24083
rect 17862 24080 17868 24132
rect 17920 24120 17926 24132
rect 20640 24120 20668 24151
rect 25406 24148 25412 24160
rect 25464 24188 25470 24200
rect 27154 24188 27160 24200
rect 25464 24160 27160 24188
rect 25464 24148 25470 24160
rect 27154 24148 27160 24160
rect 27212 24148 27218 24200
rect 17920 24092 20668 24120
rect 22005 24123 22063 24129
rect 17920 24080 17926 24092
rect 22005 24089 22017 24123
rect 22051 24089 22063 24123
rect 22005 24083 22063 24089
rect 5534 24052 5540 24064
rect 5184 24024 5540 24052
rect 5534 24012 5540 24024
rect 5592 24052 5598 24064
rect 6178 24052 6184 24064
rect 5592 24024 6184 24052
rect 5592 24012 5598 24024
rect 6178 24012 6184 24024
rect 6236 24012 6242 24064
rect 9217 24055 9275 24061
rect 9217 24021 9229 24055
rect 9263 24052 9275 24055
rect 10778 24052 10784 24064
rect 9263 24024 10784 24052
rect 9263 24021 9275 24024
rect 9217 24015 9275 24021
rect 10778 24012 10784 24024
rect 10836 24012 10842 24064
rect 14550 24012 14556 24064
rect 14608 24052 14614 24064
rect 14645 24055 14703 24061
rect 14645 24052 14657 24055
rect 14608 24024 14657 24052
rect 14608 24012 14614 24024
rect 14645 24021 14657 24024
rect 14691 24021 14703 24055
rect 14645 24015 14703 24021
rect 15562 24012 15568 24064
rect 15620 24052 15626 24064
rect 16114 24052 16120 24064
rect 15620 24024 16120 24052
rect 15620 24012 15626 24024
rect 16114 24012 16120 24024
rect 16172 24012 16178 24064
rect 18046 24012 18052 24064
rect 18104 24052 18110 24064
rect 18509 24055 18567 24061
rect 18509 24052 18521 24055
rect 18104 24024 18521 24052
rect 18104 24012 18110 24024
rect 18509 24021 18521 24024
rect 18555 24021 18567 24055
rect 18509 24015 18567 24021
rect 21269 24055 21327 24061
rect 21269 24021 21281 24055
rect 21315 24052 21327 24055
rect 21358 24052 21364 24064
rect 21315 24024 21364 24052
rect 21315 24021 21327 24024
rect 21269 24015 21327 24021
rect 21358 24012 21364 24024
rect 21416 24052 21422 24064
rect 22020 24052 22048 24083
rect 22094 24080 22100 24132
rect 22152 24120 22158 24132
rect 22649 24123 22707 24129
rect 22152 24092 22197 24120
rect 22152 24080 22158 24092
rect 22649 24089 22661 24123
rect 22695 24120 22707 24123
rect 26326 24120 26332 24132
rect 22695 24092 26332 24120
rect 22695 24089 22707 24092
rect 22649 24083 22707 24089
rect 26326 24080 26332 24092
rect 26384 24120 26390 24132
rect 27448 24120 27476 24364
rect 27617 24327 27675 24333
rect 27617 24293 27629 24327
rect 27663 24293 27675 24327
rect 27724 24324 27752 24364
rect 28994 24352 29000 24364
rect 29052 24352 29058 24404
rect 33318 24324 33324 24336
rect 27724 24296 33324 24324
rect 27617 24287 27675 24293
rect 27632 24256 27660 24287
rect 33318 24284 33324 24296
rect 33376 24284 33382 24336
rect 27632 24228 28488 24256
rect 27522 24148 27528 24200
rect 27580 24188 27586 24200
rect 28460 24197 28488 24228
rect 27801 24191 27859 24197
rect 27801 24188 27813 24191
rect 27580 24160 27813 24188
rect 27580 24148 27586 24160
rect 27801 24157 27813 24160
rect 27847 24157 27859 24191
rect 27801 24151 27859 24157
rect 28445 24191 28503 24197
rect 28445 24157 28457 24191
rect 28491 24157 28503 24191
rect 28445 24151 28503 24157
rect 28905 24191 28963 24197
rect 28905 24157 28917 24191
rect 28951 24157 28963 24191
rect 28905 24151 28963 24157
rect 26384 24092 27476 24120
rect 27816 24120 27844 24151
rect 28920 24120 28948 24151
rect 27816 24092 28948 24120
rect 26384 24080 26390 24092
rect 21416 24024 22048 24052
rect 21416 24012 21422 24024
rect 22278 24012 22284 24064
rect 22336 24052 22342 24064
rect 23201 24055 23259 24061
rect 23201 24052 23213 24055
rect 22336 24024 23213 24052
rect 22336 24012 22342 24024
rect 23201 24021 23213 24024
rect 23247 24021 23259 24055
rect 23201 24015 23259 24021
rect 25130 24012 25136 24064
rect 25188 24052 25194 24064
rect 25225 24055 25283 24061
rect 25225 24052 25237 24055
rect 25188 24024 25237 24052
rect 25188 24012 25194 24024
rect 25225 24021 25237 24024
rect 25271 24021 25283 24055
rect 28258 24052 28264 24064
rect 28219 24024 28264 24052
rect 25225 24015 25283 24021
rect 28258 24012 28264 24024
rect 28316 24012 28322 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 5902 23848 5908 23860
rect 2240 23820 5908 23848
rect 2240 23789 2268 23820
rect 5902 23808 5908 23820
rect 5960 23808 5966 23860
rect 13630 23808 13636 23860
rect 13688 23848 13694 23860
rect 15013 23851 15071 23857
rect 15013 23848 15025 23851
rect 13688 23820 15025 23848
rect 13688 23808 13694 23820
rect 15013 23817 15025 23820
rect 15059 23848 15071 23851
rect 21174 23848 21180 23860
rect 15059 23820 21180 23848
rect 15059 23817 15071 23820
rect 15013 23811 15071 23817
rect 21174 23808 21180 23820
rect 21232 23808 21238 23860
rect 21358 23848 21364 23860
rect 21319 23820 21364 23848
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 22094 23848 22100 23860
rect 22055 23820 22100 23848
rect 22094 23808 22100 23820
rect 22152 23808 22158 23860
rect 27522 23848 27528 23860
rect 22204 23820 27528 23848
rect 2225 23783 2283 23789
rect 2225 23749 2237 23783
rect 2271 23749 2283 23783
rect 5442 23780 5448 23792
rect 3450 23752 5448 23780
rect 2225 23743 2283 23749
rect 5442 23740 5448 23752
rect 5500 23740 5506 23792
rect 6733 23783 6791 23789
rect 6733 23749 6745 23783
rect 6779 23780 6791 23783
rect 6822 23780 6828 23792
rect 6779 23752 6828 23780
rect 6779 23749 6791 23752
rect 6733 23743 6791 23749
rect 6822 23740 6828 23752
rect 6880 23740 6886 23792
rect 7285 23783 7343 23789
rect 7285 23749 7297 23783
rect 7331 23780 7343 23783
rect 10686 23780 10692 23792
rect 7331 23752 10692 23780
rect 7331 23749 7343 23752
rect 7285 23743 7343 23749
rect 10686 23740 10692 23752
rect 10744 23740 10750 23792
rect 14918 23780 14924 23792
rect 14766 23752 14924 23780
rect 14918 23740 14924 23752
rect 14976 23740 14982 23792
rect 22204 23780 22232 23820
rect 27522 23808 27528 23820
rect 27580 23808 27586 23860
rect 28350 23848 28356 23860
rect 28311 23820 28356 23848
rect 28350 23808 28356 23820
rect 28408 23808 28414 23860
rect 15028 23752 22232 23780
rect 25777 23783 25835 23789
rect 7742 23712 7748 23724
rect 7703 23684 7748 23712
rect 7742 23672 7748 23684
rect 7800 23672 7806 23724
rect 1949 23647 2007 23653
rect 1949 23613 1961 23647
rect 1995 23644 2007 23647
rect 2774 23644 2780 23656
rect 1995 23616 2780 23644
rect 1995 23613 2007 23616
rect 1949 23607 2007 23613
rect 2774 23604 2780 23616
rect 2832 23644 2838 23656
rect 3970 23644 3976 23656
rect 2832 23616 3976 23644
rect 2832 23604 2838 23616
rect 3970 23604 3976 23616
rect 4028 23604 4034 23656
rect 6641 23647 6699 23653
rect 6641 23613 6653 23647
rect 6687 23644 6699 23647
rect 12342 23644 12348 23656
rect 6687 23616 12348 23644
rect 6687 23613 6699 23616
rect 6641 23607 6699 23613
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 13170 23604 13176 23656
rect 13228 23644 13234 23656
rect 13265 23647 13323 23653
rect 13265 23644 13277 23647
rect 13228 23616 13277 23644
rect 13228 23604 13234 23616
rect 13265 23613 13277 23616
rect 13311 23613 13323 23647
rect 13265 23607 13323 23613
rect 13541 23647 13599 23653
rect 13541 23613 13553 23647
rect 13587 23644 13599 23647
rect 14826 23644 14832 23656
rect 13587 23616 14832 23644
rect 13587 23613 13599 23616
rect 13541 23607 13599 23613
rect 14826 23604 14832 23616
rect 14884 23604 14890 23656
rect 3510 23536 3516 23588
rect 3568 23576 3574 23588
rect 6730 23576 6736 23588
rect 3568 23548 6736 23576
rect 3568 23536 3574 23548
rect 6730 23536 6736 23548
rect 6788 23576 6794 23588
rect 10134 23576 10140 23588
rect 6788 23548 10140 23576
rect 6788 23536 6794 23548
rect 10134 23536 10140 23548
rect 10192 23536 10198 23588
rect 15028 23576 15056 23752
rect 25777 23749 25789 23783
rect 25823 23780 25835 23783
rect 26602 23780 26608 23792
rect 25823 23752 26608 23780
rect 25823 23749 25835 23752
rect 25777 23743 25835 23749
rect 26602 23740 26608 23752
rect 26660 23740 26666 23792
rect 27341 23783 27399 23789
rect 27341 23749 27353 23783
rect 27387 23780 27399 23783
rect 27706 23780 27712 23792
rect 27387 23752 27712 23780
rect 27387 23749 27399 23752
rect 27341 23743 27399 23749
rect 27706 23740 27712 23752
rect 27764 23740 27770 23792
rect 27893 23783 27951 23789
rect 27893 23749 27905 23783
rect 27939 23780 27951 23783
rect 27982 23780 27988 23792
rect 27939 23752 27988 23780
rect 27939 23749 27951 23752
rect 27893 23743 27951 23749
rect 27982 23740 27988 23752
rect 28040 23740 28046 23792
rect 29914 23780 29920 23792
rect 29875 23752 29920 23780
rect 29914 23740 29920 23752
rect 29972 23740 29978 23792
rect 30466 23780 30472 23792
rect 30427 23752 30472 23780
rect 30466 23740 30472 23752
rect 30524 23740 30530 23792
rect 15102 23672 15108 23724
rect 15160 23712 15166 23724
rect 16390 23712 16396 23724
rect 15160 23684 16396 23712
rect 15160 23672 15166 23684
rect 16390 23672 16396 23684
rect 16448 23712 16454 23724
rect 16853 23715 16911 23721
rect 16853 23712 16865 23715
rect 16448 23684 16865 23712
rect 16448 23672 16454 23684
rect 16853 23681 16865 23684
rect 16899 23681 16911 23715
rect 18046 23712 18052 23724
rect 18007 23684 18052 23712
rect 16853 23675 16911 23681
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 19889 23715 19947 23721
rect 19889 23681 19901 23715
rect 19935 23712 19947 23715
rect 19978 23712 19984 23724
rect 19935 23684 19984 23712
rect 19935 23681 19947 23684
rect 19889 23675 19947 23681
rect 19978 23672 19984 23684
rect 20036 23672 20042 23724
rect 20346 23712 20352 23724
rect 20307 23684 20352 23712
rect 20346 23672 20352 23684
rect 20404 23712 20410 23724
rect 20714 23712 20720 23724
rect 20404 23684 20720 23712
rect 20404 23672 20410 23684
rect 20714 23672 20720 23684
rect 20772 23672 20778 23724
rect 22002 23712 22008 23724
rect 21963 23684 22008 23712
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 25130 23712 25136 23724
rect 25091 23684 25136 23712
rect 25130 23672 25136 23684
rect 25188 23672 25194 23724
rect 26326 23672 26332 23724
rect 26384 23712 26390 23724
rect 28534 23712 28540 23724
rect 26384 23684 26429 23712
rect 28495 23684 28540 23712
rect 26384 23672 26390 23684
rect 28534 23672 28540 23684
rect 28592 23672 28598 23724
rect 38286 23712 38292 23724
rect 38247 23684 38292 23712
rect 38286 23672 38292 23684
rect 38344 23672 38350 23724
rect 16758 23604 16764 23656
rect 16816 23644 16822 23656
rect 16942 23644 16948 23656
rect 16816 23616 16948 23644
rect 16816 23604 16822 23616
rect 16942 23604 16948 23616
rect 17000 23644 17006 23656
rect 17862 23644 17868 23656
rect 17000 23616 17868 23644
rect 17000 23604 17006 23616
rect 17862 23604 17868 23616
rect 17920 23644 17926 23656
rect 18601 23647 18659 23653
rect 18601 23644 18613 23647
rect 17920 23616 18613 23644
rect 17920 23604 17926 23616
rect 18601 23613 18613 23616
rect 18647 23613 18659 23647
rect 18782 23644 18788 23656
rect 18743 23616 18788 23644
rect 18601 23607 18659 23613
rect 18782 23604 18788 23616
rect 18840 23604 18846 23656
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23644 20959 23647
rect 22278 23644 22284 23656
rect 20947 23616 22284 23644
rect 20947 23613 20959 23616
rect 20901 23607 20959 23613
rect 22278 23604 22284 23616
rect 22336 23604 22342 23656
rect 23290 23644 23296 23656
rect 23251 23616 23296 23644
rect 23290 23604 23296 23616
rect 23348 23604 23354 23656
rect 25222 23604 25228 23656
rect 25280 23644 25286 23656
rect 25685 23647 25743 23653
rect 25685 23644 25697 23647
rect 25280 23616 25697 23644
rect 25280 23604 25286 23616
rect 25685 23613 25697 23616
rect 25731 23613 25743 23647
rect 25685 23607 25743 23613
rect 27249 23647 27307 23653
rect 27249 23613 27261 23647
rect 27295 23613 27307 23647
rect 29822 23644 29828 23656
rect 29783 23616 29828 23644
rect 27249 23607 27307 23613
rect 21082 23576 21088 23588
rect 14936 23548 15056 23576
rect 15120 23548 21088 23576
rect 3694 23508 3700 23520
rect 3655 23480 3700 23508
rect 3694 23468 3700 23480
rect 3752 23508 3758 23520
rect 5166 23508 5172 23520
rect 3752 23480 5172 23508
rect 3752 23468 3758 23480
rect 5166 23468 5172 23480
rect 5224 23468 5230 23520
rect 7834 23508 7840 23520
rect 7795 23480 7840 23508
rect 7834 23468 7840 23480
rect 7892 23468 7898 23520
rect 10594 23468 10600 23520
rect 10652 23508 10658 23520
rect 14936 23508 14964 23548
rect 10652 23480 14964 23508
rect 10652 23468 10658 23480
rect 15010 23468 15016 23520
rect 15068 23508 15074 23520
rect 15120 23508 15148 23548
rect 21082 23536 21088 23548
rect 21140 23536 21146 23588
rect 27264 23576 27292 23607
rect 29822 23604 29828 23616
rect 29880 23604 29886 23656
rect 30098 23576 30104 23588
rect 27264 23548 30104 23576
rect 30098 23536 30104 23548
rect 30156 23536 30162 23588
rect 15068 23480 15148 23508
rect 15068 23468 15074 23480
rect 15194 23468 15200 23520
rect 15252 23508 15258 23520
rect 16945 23511 17003 23517
rect 16945 23508 16957 23511
rect 15252 23480 16957 23508
rect 15252 23468 15258 23480
rect 16945 23477 16957 23480
rect 16991 23477 17003 23511
rect 17862 23508 17868 23520
rect 17823 23480 17868 23508
rect 16945 23471 17003 23477
rect 17862 23468 17868 23480
rect 17920 23468 17926 23520
rect 18598 23468 18604 23520
rect 18656 23508 18662 23520
rect 18969 23511 19027 23517
rect 18969 23508 18981 23511
rect 18656 23480 18981 23508
rect 18656 23468 18662 23480
rect 18969 23477 18981 23480
rect 19015 23477 19027 23511
rect 19702 23508 19708 23520
rect 19663 23480 19708 23508
rect 18969 23471 19027 23477
rect 19702 23468 19708 23480
rect 19760 23468 19766 23520
rect 24946 23508 24952 23520
rect 24907 23480 24952 23508
rect 24946 23468 24952 23480
rect 25004 23468 25010 23520
rect 36446 23468 36452 23520
rect 36504 23508 36510 23520
rect 38105 23511 38163 23517
rect 38105 23508 38117 23511
rect 36504 23480 38117 23508
rect 36504 23468 36510 23480
rect 38105 23477 38117 23480
rect 38151 23477 38163 23511
rect 38105 23471 38163 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 5718 23304 5724 23316
rect 5679 23276 5724 23304
rect 5718 23264 5724 23276
rect 5776 23264 5782 23316
rect 7374 23264 7380 23316
rect 7432 23304 7438 23316
rect 18233 23307 18291 23313
rect 7432 23276 16436 23304
rect 7432 23264 7438 23276
rect 11146 23236 11152 23248
rect 11107 23208 11152 23236
rect 11146 23196 11152 23208
rect 11204 23196 11210 23248
rect 16408 23236 16436 23276
rect 18233 23273 18245 23307
rect 18279 23304 18291 23307
rect 18782 23304 18788 23316
rect 18279 23276 18788 23304
rect 18279 23273 18291 23276
rect 18233 23267 18291 23273
rect 18782 23264 18788 23276
rect 18840 23264 18846 23316
rect 26602 23304 26608 23316
rect 26563 23276 26608 23304
rect 26602 23264 26608 23276
rect 26660 23264 26666 23316
rect 27985 23307 28043 23313
rect 27985 23273 27997 23307
rect 28031 23304 28043 23307
rect 29822 23304 29828 23316
rect 28031 23276 29828 23304
rect 28031 23273 28043 23276
rect 27985 23267 28043 23273
rect 29822 23264 29828 23276
rect 29880 23264 29886 23316
rect 19426 23236 19432 23248
rect 16408 23208 19432 23236
rect 4249 23171 4307 23177
rect 4249 23137 4261 23171
rect 4295 23168 4307 23171
rect 4614 23168 4620 23180
rect 4295 23140 4620 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 4614 23128 4620 23140
rect 4672 23168 4678 23180
rect 4982 23168 4988 23180
rect 4672 23140 4988 23168
rect 4672 23128 4678 23140
rect 4982 23128 4988 23140
rect 5040 23128 5046 23180
rect 1578 23100 1584 23112
rect 1539 23072 1584 23100
rect 1578 23060 1584 23072
rect 1636 23060 1642 23112
rect 3970 23100 3976 23112
rect 3931 23072 3976 23100
rect 3970 23060 3976 23072
rect 4028 23060 4034 23112
rect 11164 23100 11192 23196
rect 11517 23171 11575 23177
rect 11517 23137 11529 23171
rect 11563 23168 11575 23171
rect 13170 23168 13176 23180
rect 11563 23140 13176 23168
rect 11563 23137 11575 23140
rect 11517 23131 11575 23137
rect 13170 23128 13176 23140
rect 13228 23128 13234 23180
rect 13262 23128 13268 23180
rect 13320 23168 13326 23180
rect 16408 23177 16436 23208
rect 19426 23196 19432 23208
rect 19484 23196 19490 23248
rect 19794 23236 19800 23248
rect 19755 23208 19800 23236
rect 19794 23196 19800 23208
rect 19852 23196 19858 23248
rect 20254 23196 20260 23248
rect 20312 23236 20318 23248
rect 20533 23239 20591 23245
rect 20533 23236 20545 23239
rect 20312 23208 20545 23236
rect 20312 23196 20318 23208
rect 20533 23205 20545 23208
rect 20579 23205 20591 23239
rect 20533 23199 20591 23205
rect 22833 23239 22891 23245
rect 22833 23205 22845 23239
rect 22879 23236 22891 23239
rect 23661 23239 23719 23245
rect 23661 23236 23673 23239
rect 22879 23208 23673 23236
rect 22879 23205 22891 23208
rect 22833 23199 22891 23205
rect 23661 23205 23673 23208
rect 23707 23236 23719 23239
rect 24762 23236 24768 23248
rect 23707 23208 24768 23236
rect 23707 23205 23719 23208
rect 23661 23199 23719 23205
rect 24762 23196 24768 23208
rect 24820 23196 24826 23248
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 13320 23140 13553 23168
rect 13320 23128 13326 23140
rect 13541 23137 13553 23140
rect 13587 23168 13599 23171
rect 16393 23171 16451 23177
rect 13587 23140 16252 23168
rect 13587 23137 13599 23140
rect 13541 23131 13599 23137
rect 14550 23100 14556 23112
rect 11164 23072 11376 23100
rect 12926 23072 14556 23100
rect 11348 23032 11376 23072
rect 14550 23060 14556 23072
rect 14608 23060 14614 23112
rect 14737 23103 14795 23109
rect 14737 23069 14749 23103
rect 14783 23069 14795 23103
rect 14737 23063 14795 23069
rect 11790 23032 11796 23044
rect 5474 23004 11284 23032
rect 11348 23004 11796 23032
rect 1762 22964 1768 22976
rect 1723 22936 1768 22964
rect 1762 22924 1768 22936
rect 1820 22924 1826 22976
rect 11256 22964 11284 23004
rect 11790 22992 11796 23004
rect 11848 22992 11854 23044
rect 13814 22992 13820 23044
rect 13872 23032 13878 23044
rect 14752 23032 14780 23063
rect 15286 23060 15292 23112
rect 15344 23100 15350 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 15344 23072 15393 23100
rect 15344 23060 15350 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 15381 23063 15439 23069
rect 13872 23004 14780 23032
rect 13872 22992 13878 23004
rect 14829 22967 14887 22973
rect 14829 22964 14841 22967
rect 11256 22936 14841 22964
rect 14829 22933 14841 22936
rect 14875 22933 14887 22967
rect 14829 22927 14887 22933
rect 15473 22967 15531 22973
rect 15473 22933 15485 22967
rect 15519 22964 15531 22967
rect 15654 22964 15660 22976
rect 15519 22936 15660 22964
rect 15519 22933 15531 22936
rect 15473 22927 15531 22933
rect 15654 22924 15660 22936
rect 15712 22924 15718 22976
rect 16224 22964 16252 23140
rect 16393 23137 16405 23171
rect 16439 23137 16451 23171
rect 16758 23168 16764 23180
rect 16719 23140 16764 23168
rect 16393 23131 16451 23137
rect 16758 23128 16764 23140
rect 16816 23128 16822 23180
rect 17052 23140 19656 23168
rect 16482 22992 16488 23044
rect 16540 23032 16546 23044
rect 16540 23004 16585 23032
rect 16540 22992 16546 23004
rect 17052 22964 17080 23140
rect 17126 23060 17132 23112
rect 17184 23100 17190 23112
rect 17497 23103 17555 23109
rect 17497 23100 17509 23103
rect 17184 23072 17509 23100
rect 17184 23060 17190 23072
rect 17497 23069 17509 23072
rect 17543 23069 17555 23103
rect 17497 23063 17555 23069
rect 17954 23060 17960 23112
rect 18012 23100 18018 23112
rect 18141 23103 18199 23109
rect 18141 23100 18153 23103
rect 18012 23072 18153 23100
rect 18012 23060 18018 23072
rect 18141 23069 18153 23072
rect 18187 23100 18199 23103
rect 18690 23100 18696 23112
rect 18187 23072 18696 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 18690 23060 18696 23072
rect 18748 23060 18754 23112
rect 19521 23103 19579 23109
rect 19521 23069 19533 23103
rect 19567 23069 19579 23103
rect 19521 23063 19579 23069
rect 18230 22992 18236 23044
rect 18288 23032 18294 23044
rect 19536 23032 19564 23063
rect 18288 23004 19564 23032
rect 19628 23032 19656 23140
rect 19702 23128 19708 23180
rect 19760 23168 19766 23180
rect 20349 23171 20407 23177
rect 20349 23168 20361 23171
rect 19760 23140 20361 23168
rect 19760 23128 19766 23140
rect 20349 23137 20361 23140
rect 20395 23137 20407 23171
rect 22186 23168 22192 23180
rect 22147 23140 22192 23168
rect 20349 23131 20407 23137
rect 22186 23128 22192 23140
rect 22244 23128 22250 23180
rect 23290 23168 23296 23180
rect 23251 23140 23296 23168
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 23477 23171 23535 23177
rect 23477 23137 23489 23171
rect 23523 23168 23535 23171
rect 24946 23168 24952 23180
rect 23523 23140 24952 23168
rect 23523 23137 23535 23140
rect 23477 23131 23535 23137
rect 24946 23128 24952 23140
rect 25004 23128 25010 23180
rect 27341 23171 27399 23177
rect 27341 23137 27353 23171
rect 27387 23168 27399 23171
rect 28445 23171 28503 23177
rect 28445 23168 28457 23171
rect 27387 23140 28457 23168
rect 27387 23137 27399 23140
rect 27341 23131 27399 23137
rect 28445 23137 28457 23140
rect 28491 23137 28503 23171
rect 28445 23131 28503 23137
rect 19794 23060 19800 23112
rect 19852 23100 19858 23112
rect 20165 23103 20223 23109
rect 20165 23100 20177 23103
rect 19852 23072 20177 23100
rect 19852 23060 19858 23072
rect 20165 23069 20177 23072
rect 20211 23069 20223 23103
rect 20165 23063 20223 23069
rect 21358 23060 21364 23112
rect 21416 23100 21422 23112
rect 22373 23103 22431 23109
rect 22373 23100 22385 23103
rect 21416 23072 22385 23100
rect 21416 23060 21422 23072
rect 22373 23069 22385 23072
rect 22419 23069 22431 23103
rect 22373 23063 22431 23069
rect 25593 23103 25651 23109
rect 25593 23069 25605 23103
rect 25639 23069 25651 23103
rect 26789 23103 26847 23109
rect 26789 23100 26801 23103
rect 25593 23063 25651 23069
rect 26206 23072 26801 23100
rect 20622 23032 20628 23044
rect 19628 23004 20628 23032
rect 18288 22992 18294 23004
rect 20622 22992 20628 23004
rect 20680 22992 20686 23044
rect 20806 22992 20812 23044
rect 20864 23032 20870 23044
rect 22002 23032 22008 23044
rect 20864 23004 22008 23032
rect 20864 22992 20870 23004
rect 22002 22992 22008 23004
rect 22060 23032 22066 23044
rect 25608 23032 25636 23063
rect 22060 23004 25636 23032
rect 22060 22992 22066 23004
rect 16224 22936 17080 22964
rect 17589 22967 17647 22973
rect 17589 22933 17601 22967
rect 17635 22964 17647 22967
rect 18690 22964 18696 22976
rect 17635 22936 18696 22964
rect 17635 22933 17647 22936
rect 17589 22927 17647 22933
rect 18690 22924 18696 22936
rect 18748 22924 18754 22976
rect 19334 22964 19340 22976
rect 19295 22936 19340 22964
rect 19334 22924 19340 22936
rect 19392 22924 19398 22976
rect 25409 22967 25467 22973
rect 25409 22933 25421 22967
rect 25455 22964 25467 22967
rect 26206 22964 26234 23072
rect 26789 23069 26801 23072
rect 26835 23069 26847 23103
rect 26789 23063 26847 23069
rect 27525 23103 27583 23109
rect 27525 23069 27537 23103
rect 27571 23100 27583 23103
rect 28258 23100 28264 23112
rect 27571 23072 28264 23100
rect 27571 23069 27583 23072
rect 27525 23063 27583 23069
rect 28258 23060 28264 23072
rect 28316 23060 28322 23112
rect 25455 22936 26234 22964
rect 25455 22933 25467 22936
rect 25409 22927 25467 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 6454 22720 6460 22772
rect 6512 22760 6518 22772
rect 16209 22763 16267 22769
rect 6512 22732 15608 22760
rect 6512 22720 6518 22732
rect 2041 22695 2099 22701
rect 2041 22661 2053 22695
rect 2087 22692 2099 22695
rect 2682 22692 2688 22704
rect 2087 22664 2688 22692
rect 2087 22661 2099 22664
rect 2041 22655 2099 22661
rect 2682 22652 2688 22664
rect 2740 22652 2746 22704
rect 9122 22692 9128 22704
rect 8864 22664 9128 22692
rect 2593 22627 2651 22633
rect 2593 22593 2605 22627
rect 2639 22624 2651 22627
rect 7374 22624 7380 22636
rect 2639 22596 7380 22624
rect 2639 22593 2651 22596
rect 2593 22587 2651 22593
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22624 7619 22627
rect 7742 22624 7748 22636
rect 7607 22596 7748 22624
rect 7607 22593 7619 22596
rect 7561 22587 7619 22593
rect 7742 22584 7748 22596
rect 7800 22584 7806 22636
rect 8202 22624 8208 22636
rect 8163 22596 8208 22624
rect 8202 22584 8208 22596
rect 8260 22584 8266 22636
rect 8864 22633 8892 22664
rect 9122 22652 9128 22664
rect 9180 22652 9186 22704
rect 15473 22695 15531 22701
rect 15473 22692 15485 22695
rect 10350 22664 15485 22692
rect 15473 22661 15485 22664
rect 15519 22661 15531 22695
rect 15580 22692 15608 22732
rect 16209 22729 16221 22763
rect 16255 22760 16267 22763
rect 16482 22760 16488 22772
rect 16255 22732 16488 22760
rect 16255 22729 16267 22732
rect 16209 22723 16267 22729
rect 16482 22720 16488 22732
rect 16540 22720 16546 22772
rect 19613 22763 19671 22769
rect 16592 22732 18092 22760
rect 16592 22692 16620 22732
rect 17494 22692 17500 22704
rect 15580 22664 16620 22692
rect 17455 22664 17500 22692
rect 15473 22655 15531 22661
rect 17494 22652 17500 22664
rect 17552 22652 17558 22704
rect 18064 22701 18092 22732
rect 19613 22729 19625 22763
rect 19659 22760 19671 22763
rect 19978 22760 19984 22772
rect 19659 22732 19984 22760
rect 19659 22729 19671 22732
rect 19613 22723 19671 22729
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 21358 22760 21364 22772
rect 21319 22732 21364 22760
rect 21358 22720 21364 22732
rect 21416 22720 21422 22772
rect 25869 22763 25927 22769
rect 25869 22760 25881 22763
rect 24872 22732 25881 22760
rect 18049 22695 18107 22701
rect 18049 22661 18061 22695
rect 18095 22661 18107 22695
rect 20346 22692 20352 22704
rect 18049 22655 18107 22661
rect 18524 22664 20352 22692
rect 8849 22627 8907 22633
rect 8849 22593 8861 22627
rect 8895 22593 8907 22627
rect 8849 22587 8907 22593
rect 10594 22584 10600 22636
rect 10652 22624 10658 22636
rect 10873 22627 10931 22633
rect 10873 22624 10885 22627
rect 10652 22596 10885 22624
rect 10652 22584 10658 22596
rect 10873 22593 10885 22596
rect 10919 22593 10931 22627
rect 10873 22587 10931 22593
rect 15286 22584 15292 22636
rect 15344 22624 15350 22636
rect 15381 22627 15439 22633
rect 15381 22624 15393 22627
rect 15344 22596 15393 22624
rect 15344 22584 15350 22596
rect 15381 22593 15393 22596
rect 15427 22593 15439 22627
rect 15381 22587 15439 22593
rect 15562 22584 15568 22636
rect 15620 22624 15626 22636
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 15620 22596 16129 22624
rect 15620 22584 15626 22596
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 18524 22624 18552 22664
rect 20346 22652 20352 22664
rect 20404 22652 20410 22704
rect 24762 22692 24768 22704
rect 24723 22664 24768 22692
rect 24762 22652 24768 22664
rect 24820 22652 24826 22704
rect 24872 22701 24900 22732
rect 25869 22729 25881 22732
rect 25915 22729 25927 22763
rect 25869 22723 25927 22729
rect 24857 22695 24915 22701
rect 24857 22661 24869 22695
rect 24903 22661 24915 22695
rect 27338 22692 27344 22704
rect 27299 22664 27344 22692
rect 24857 22655 24915 22661
rect 27338 22652 27344 22664
rect 27396 22652 27402 22704
rect 18690 22624 18696 22636
rect 16117 22587 16175 22593
rect 18064 22596 18552 22624
rect 18651 22596 18696 22624
rect 1949 22559 2007 22565
rect 1949 22525 1961 22559
rect 1995 22556 2007 22559
rect 2130 22556 2136 22568
rect 1995 22528 2136 22556
rect 1995 22525 2007 22528
rect 1949 22519 2007 22525
rect 2130 22516 2136 22528
rect 2188 22516 2194 22568
rect 9125 22559 9183 22565
rect 9125 22525 9137 22559
rect 9171 22556 9183 22559
rect 17405 22559 17463 22565
rect 9171 22528 10824 22556
rect 9171 22525 9183 22528
rect 9125 22519 9183 22525
rect 4614 22448 4620 22500
rect 4672 22488 4678 22500
rect 8297 22491 8355 22497
rect 8297 22488 8309 22491
rect 4672 22460 8309 22488
rect 4672 22448 4678 22460
rect 8297 22457 8309 22460
rect 8343 22457 8355 22491
rect 10796 22488 10824 22528
rect 17405 22525 17417 22559
rect 17451 22556 17463 22559
rect 18064 22556 18092 22596
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 19797 22627 19855 22633
rect 19797 22593 19809 22627
rect 19843 22624 19855 22627
rect 20070 22624 20076 22636
rect 19843 22596 20076 22624
rect 19843 22593 19855 22596
rect 19797 22587 19855 22593
rect 20070 22584 20076 22596
rect 20128 22584 20134 22636
rect 20622 22584 20628 22636
rect 20680 22624 20686 22636
rect 21269 22627 21327 22633
rect 21269 22624 21281 22627
rect 20680 22596 21281 22624
rect 20680 22584 20686 22596
rect 21269 22593 21281 22596
rect 21315 22593 21327 22627
rect 26050 22624 26056 22636
rect 26011 22596 26056 22624
rect 21269 22587 21327 22593
rect 17451 22528 18092 22556
rect 17451 22525 17463 22528
rect 17405 22519 17463 22525
rect 18138 22516 18144 22568
rect 18196 22556 18202 22568
rect 18509 22559 18567 22565
rect 18509 22556 18521 22559
rect 18196 22528 18521 22556
rect 18196 22516 18202 22528
rect 18509 22525 18521 22528
rect 18555 22525 18567 22559
rect 21284 22556 21312 22587
rect 26050 22584 26056 22596
rect 26108 22584 26114 22636
rect 25406 22556 25412 22568
rect 21284 22528 25412 22556
rect 18509 22519 18567 22525
rect 25406 22516 25412 22528
rect 25464 22516 25470 22568
rect 27249 22559 27307 22565
rect 27249 22525 27261 22559
rect 27295 22556 27307 22559
rect 27614 22556 27620 22568
rect 27295 22528 27620 22556
rect 27295 22525 27307 22528
rect 27249 22519 27307 22525
rect 27614 22516 27620 22528
rect 27672 22516 27678 22568
rect 27706 22516 27712 22568
rect 27764 22556 27770 22568
rect 28350 22556 28356 22568
rect 27764 22528 27809 22556
rect 28311 22528 28356 22556
rect 27764 22516 27770 22528
rect 28350 22516 28356 22528
rect 28408 22516 28414 22568
rect 12158 22488 12164 22500
rect 10796 22460 12164 22488
rect 8297 22451 8355 22457
rect 12158 22448 12164 22460
rect 12216 22488 12222 22500
rect 17770 22488 17776 22500
rect 12216 22460 17776 22488
rect 12216 22448 12222 22460
rect 17770 22448 17776 22460
rect 17828 22448 17834 22500
rect 25317 22491 25375 22497
rect 18064 22460 22094 22488
rect 7558 22380 7564 22432
rect 7616 22420 7622 22432
rect 7653 22423 7711 22429
rect 7653 22420 7665 22423
rect 7616 22392 7665 22420
rect 7616 22380 7622 22392
rect 7653 22389 7665 22392
rect 7699 22389 7711 22423
rect 7653 22383 7711 22389
rect 7742 22380 7748 22432
rect 7800 22420 7806 22432
rect 9490 22420 9496 22432
rect 7800 22392 9496 22420
rect 7800 22380 7806 22392
rect 9490 22380 9496 22392
rect 9548 22380 9554 22432
rect 11790 22380 11796 22432
rect 11848 22420 11854 22432
rect 18064 22420 18092 22460
rect 18874 22420 18880 22432
rect 11848 22392 18092 22420
rect 18835 22392 18880 22420
rect 11848 22380 11854 22392
rect 18874 22380 18880 22392
rect 18932 22380 18938 22432
rect 22066 22420 22094 22460
rect 25317 22457 25329 22491
rect 25363 22488 25375 22491
rect 27724 22488 27752 22516
rect 25363 22460 27752 22488
rect 25363 22457 25375 22460
rect 25317 22451 25375 22457
rect 28534 22420 28540 22432
rect 22066 22392 28540 22420
rect 28534 22380 28540 22392
rect 28592 22380 28598 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 1844 22219 1902 22225
rect 1844 22185 1856 22219
rect 1890 22216 1902 22219
rect 3694 22216 3700 22228
rect 1890 22188 3700 22216
rect 1890 22185 1902 22188
rect 1844 22179 1902 22185
rect 3694 22176 3700 22188
rect 3752 22176 3758 22228
rect 8294 22216 8300 22228
rect 7852 22188 8300 22216
rect 1581 22083 1639 22089
rect 1581 22049 1593 22083
rect 1627 22080 1639 22083
rect 2222 22080 2228 22092
rect 1627 22052 2228 22080
rect 1627 22049 1639 22052
rect 1581 22043 1639 22049
rect 2222 22040 2228 22052
rect 2280 22040 2286 22092
rect 6825 22083 6883 22089
rect 6825 22049 6837 22083
rect 6871 22080 6883 22083
rect 7852 22080 7880 22188
rect 8294 22176 8300 22188
rect 8352 22216 8358 22228
rect 9582 22216 9588 22228
rect 8352 22188 9588 22216
rect 8352 22176 8358 22188
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 17770 22176 17776 22228
rect 17828 22216 17834 22228
rect 18230 22216 18236 22228
rect 17828 22188 18236 22216
rect 17828 22176 17834 22188
rect 18230 22176 18236 22188
rect 18288 22176 18294 22228
rect 20073 22219 20131 22225
rect 20073 22185 20085 22219
rect 20119 22216 20131 22219
rect 20254 22216 20260 22228
rect 20119 22188 20260 22216
rect 20119 22185 20131 22188
rect 20073 22179 20131 22185
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 26050 22216 26056 22228
rect 26011 22188 26056 22216
rect 26050 22176 26056 22188
rect 26108 22176 26114 22228
rect 27249 22219 27307 22225
rect 27249 22185 27261 22219
rect 27295 22216 27307 22219
rect 27338 22216 27344 22228
rect 27295 22188 27344 22216
rect 27295 22185 27307 22188
rect 27249 22179 27307 22185
rect 27338 22176 27344 22188
rect 27396 22176 27402 22228
rect 11808 22120 13216 22148
rect 8570 22080 8576 22092
rect 6871 22052 7880 22080
rect 8531 22052 8576 22080
rect 6871 22049 6883 22052
rect 6825 22043 6883 22049
rect 8570 22040 8576 22052
rect 8628 22040 8634 22092
rect 11808 22080 11836 22120
rect 13188 22092 13216 22120
rect 16022 22108 16028 22160
rect 16080 22148 16086 22160
rect 20806 22148 20812 22160
rect 16080 22120 20812 22148
rect 16080 22108 16086 22120
rect 20806 22108 20812 22120
rect 20864 22108 20870 22160
rect 24581 22151 24639 22157
rect 24581 22148 24593 22151
rect 23124 22120 23336 22148
rect 10520 22052 11836 22080
rect 6546 22012 6552 22024
rect 6507 21984 6552 22012
rect 6546 21972 6552 21984
rect 6604 21972 6610 22024
rect 9582 22012 9588 22024
rect 9543 21984 9588 22012
rect 9582 21972 9588 21984
rect 9640 21972 9646 22024
rect 10520 22021 10548 22052
rect 12894 22040 12900 22092
rect 12952 22080 12958 22092
rect 13170 22080 13176 22092
rect 12952 22052 13176 22080
rect 12952 22040 12958 22052
rect 13170 22040 13176 22052
rect 13228 22080 13234 22092
rect 14277 22083 14335 22089
rect 14277 22080 14289 22083
rect 13228 22052 14289 22080
rect 13228 22040 13234 22052
rect 14277 22049 14289 22052
rect 14323 22049 14335 22083
rect 14277 22043 14335 22049
rect 14553 22083 14611 22089
rect 14553 22049 14565 22083
rect 14599 22080 14611 22083
rect 15930 22080 15936 22092
rect 14599 22052 15936 22080
rect 14599 22049 14611 22052
rect 14553 22043 14611 22049
rect 15930 22040 15936 22052
rect 15988 22040 15994 22092
rect 17862 22040 17868 22092
rect 17920 22080 17926 22092
rect 18141 22083 18199 22089
rect 18141 22080 18153 22083
rect 17920 22052 18153 22080
rect 17920 22040 17926 22052
rect 18141 22049 18153 22052
rect 18187 22049 18199 22083
rect 18141 22043 18199 22049
rect 21177 22083 21235 22089
rect 21177 22049 21189 22083
rect 21223 22080 21235 22083
rect 21266 22080 21272 22092
rect 21223 22052 21272 22080
rect 21223 22049 21235 22052
rect 21177 22043 21235 22049
rect 21266 22040 21272 22052
rect 21324 22040 21330 22092
rect 23124 22080 23152 22120
rect 22204 22052 23152 22080
rect 23308 22080 23336 22120
rect 23952 22120 24593 22148
rect 23952 22080 23980 22120
rect 24581 22117 24593 22120
rect 24627 22117 24639 22151
rect 28902 22148 28908 22160
rect 28863 22120 28908 22148
rect 24581 22111 24639 22117
rect 28902 22108 28908 22120
rect 28960 22108 28966 22160
rect 23308 22052 23980 22080
rect 24029 22083 24087 22089
rect 10505 22015 10563 22021
rect 10505 21981 10517 22015
rect 10551 21981 10563 22015
rect 13541 22015 13599 22021
rect 11914 21984 13492 22012
rect 10505 21975 10563 21981
rect 4614 21944 4620 21956
rect 3082 21916 4620 21944
rect 4614 21904 4620 21916
rect 4672 21904 4678 21956
rect 7834 21904 7840 21956
rect 7892 21904 7898 21956
rect 9490 21904 9496 21956
rect 9548 21944 9554 21956
rect 10520 21944 10548 21975
rect 9548 21916 10548 21944
rect 10781 21947 10839 21953
rect 9548 21904 9554 21916
rect 10781 21913 10793 21947
rect 10827 21944 10839 21947
rect 11054 21944 11060 21956
rect 10827 21916 11060 21944
rect 10827 21913 10839 21916
rect 10781 21907 10839 21913
rect 11054 21904 11060 21916
rect 11112 21904 11118 21956
rect 12526 21944 12532 21956
rect 12487 21916 12532 21944
rect 12526 21904 12532 21916
rect 12584 21904 12590 21956
rect 13464 21944 13492 21984
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 17313 22015 17371 22021
rect 13587 21984 14320 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 14292 21944 14320 21984
rect 17313 21981 17325 22015
rect 17359 21981 17371 22015
rect 17313 21975 17371 21981
rect 17957 22015 18015 22021
rect 17957 21981 17969 22015
rect 18003 22012 18015 22015
rect 19150 22012 19156 22024
rect 18003 21984 19156 22012
rect 18003 21981 18015 21984
rect 17957 21975 18015 21981
rect 14458 21944 14464 21956
rect 13464 21916 13768 21944
rect 14292 21916 14464 21944
rect 3329 21879 3387 21885
rect 3329 21845 3341 21879
rect 3375 21876 3387 21879
rect 9398 21876 9404 21888
rect 3375 21848 9404 21876
rect 3375 21845 3387 21848
rect 3329 21839 3387 21845
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 9674 21876 9680 21888
rect 9635 21848 9680 21876
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 11146 21836 11152 21888
rect 11204 21876 11210 21888
rect 13633 21879 13691 21885
rect 13633 21876 13645 21879
rect 11204 21848 13645 21876
rect 11204 21836 11210 21848
rect 13633 21845 13645 21848
rect 13679 21845 13691 21879
rect 13740 21876 13768 21916
rect 14458 21904 14464 21916
rect 14516 21904 14522 21956
rect 14550 21904 14556 21956
rect 14608 21944 14614 21956
rect 16301 21947 16359 21953
rect 14608 21916 15042 21944
rect 14608 21904 14614 21916
rect 16301 21913 16313 21947
rect 16347 21944 16359 21947
rect 16390 21944 16396 21956
rect 16347 21916 16396 21944
rect 16347 21913 16359 21916
rect 16301 21907 16359 21913
rect 16390 21904 16396 21916
rect 16448 21904 16454 21956
rect 17328 21944 17356 21975
rect 19150 21972 19156 21984
rect 19208 21972 19214 22024
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 22012 19671 22015
rect 20162 22012 20168 22024
rect 19659 21984 20168 22012
rect 19659 21981 19671 21984
rect 19613 21975 19671 21981
rect 19444 21944 19472 21975
rect 20162 21972 20168 21984
rect 20220 21972 20226 22024
rect 20530 22012 20536 22024
rect 20491 21984 20536 22012
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 20717 22015 20775 22021
rect 20717 21981 20729 22015
rect 20763 22012 20775 22015
rect 22204 22012 22232 22052
rect 24029 22049 24041 22083
rect 24075 22080 24087 22083
rect 24118 22080 24124 22092
rect 24075 22052 24124 22080
rect 24075 22049 24087 22052
rect 24029 22043 24087 22049
rect 24118 22040 24124 22052
rect 24176 22040 24182 22092
rect 28350 22080 28356 22092
rect 28311 22052 28356 22080
rect 28350 22040 28356 22052
rect 28408 22040 28414 22092
rect 37274 22080 37280 22092
rect 30116 22052 37280 22080
rect 20763 21984 22232 22012
rect 22281 22015 22339 22021
rect 20763 21981 20775 21984
rect 20717 21975 20775 21981
rect 22281 21981 22293 22015
rect 22327 22012 22339 22015
rect 22370 22012 22376 22024
rect 22327 21984 22376 22012
rect 22327 21981 22339 21984
rect 22281 21975 22339 21981
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 24210 21972 24216 22024
rect 24268 22012 24274 22024
rect 30116 22021 30144 22052
rect 37274 22040 37280 22052
rect 37332 22040 37338 22092
rect 24765 22015 24823 22021
rect 24765 22012 24777 22015
rect 24268 21984 24777 22012
rect 24268 21972 24274 21984
rect 24765 21981 24777 21984
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 26237 22015 26295 22021
rect 26237 21981 26249 22015
rect 26283 22012 26295 22015
rect 27157 22015 27215 22021
rect 26283 21984 26317 22012
rect 26283 21981 26295 21984
rect 26237 21975 26295 21981
rect 27157 21981 27169 22015
rect 27203 21981 27215 22015
rect 27157 21975 27215 21981
rect 30101 22015 30159 22021
rect 30101 21981 30113 22015
rect 30147 21981 30159 22015
rect 30101 21975 30159 21981
rect 23106 21944 23112 21956
rect 17328 21916 19380 21944
rect 19444 21916 23112 21944
rect 15194 21876 15200 21888
rect 13740 21848 15200 21876
rect 13633 21839 13691 21845
rect 15194 21836 15200 21848
rect 15252 21836 15258 21888
rect 16666 21836 16672 21888
rect 16724 21876 16730 21888
rect 17126 21876 17132 21888
rect 16724 21848 17132 21876
rect 16724 21836 16730 21848
rect 17126 21836 17132 21848
rect 17184 21836 17190 21888
rect 17402 21876 17408 21888
rect 17363 21848 17408 21876
rect 17402 21836 17408 21848
rect 17460 21836 17466 21888
rect 18414 21836 18420 21888
rect 18472 21876 18478 21888
rect 18598 21876 18604 21888
rect 18472 21848 18604 21876
rect 18472 21836 18478 21848
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 19352 21876 19380 21916
rect 23106 21904 23112 21916
rect 23164 21904 23170 21956
rect 23198 21904 23204 21956
rect 23256 21944 23262 21956
rect 23385 21947 23443 21953
rect 23385 21944 23397 21947
rect 23256 21916 23397 21944
rect 23256 21904 23262 21916
rect 23385 21913 23397 21916
rect 23431 21913 23443 21947
rect 23385 21907 23443 21913
rect 23477 21947 23535 21953
rect 23477 21913 23489 21947
rect 23523 21913 23535 21947
rect 23477 21907 23535 21913
rect 20806 21876 20812 21888
rect 19352 21848 20812 21876
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 22373 21879 22431 21885
rect 22373 21845 22385 21879
rect 22419 21876 22431 21879
rect 23492 21876 23520 21907
rect 23566 21904 23572 21956
rect 23624 21944 23630 21956
rect 26252 21944 26280 21975
rect 27172 21944 27200 21975
rect 30926 21972 30932 22024
rect 30984 22012 30990 22024
rect 38013 22015 38071 22021
rect 38013 22012 38025 22015
rect 30984 21984 38025 22012
rect 30984 21972 30990 21984
rect 38013 21981 38025 21984
rect 38059 21981 38071 22015
rect 38013 21975 38071 21981
rect 28442 21944 28448 21956
rect 23624 21916 27200 21944
rect 28403 21916 28448 21944
rect 23624 21904 23630 21916
rect 28442 21904 28448 21916
rect 28500 21904 28506 21956
rect 30190 21876 30196 21888
rect 22419 21848 23520 21876
rect 30151 21848 30196 21876
rect 22419 21845 22431 21848
rect 22373 21839 22431 21845
rect 30190 21836 30196 21848
rect 30248 21836 30254 21888
rect 38194 21876 38200 21888
rect 38155 21848 38200 21876
rect 38194 21836 38200 21848
rect 38252 21836 38258 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 6178 21632 6184 21684
rect 6236 21672 6242 21684
rect 14550 21672 14556 21684
rect 6236 21644 12434 21672
rect 14511 21644 14556 21672
rect 6236 21632 6242 21644
rect 4798 21564 4804 21616
rect 4856 21604 4862 21616
rect 4856 21576 7314 21604
rect 4856 21564 4862 21576
rect 9398 21564 9404 21616
rect 9456 21604 9462 21616
rect 12250 21604 12256 21616
rect 9456 21576 12256 21604
rect 9456 21564 9462 21576
rect 12250 21564 12256 21576
rect 12308 21564 12314 21616
rect 12406 21604 12434 21644
rect 14550 21632 14556 21644
rect 14608 21632 14614 21684
rect 16945 21675 17003 21681
rect 16945 21641 16957 21675
rect 16991 21672 17003 21675
rect 17494 21672 17500 21684
rect 16991 21644 17500 21672
rect 16991 21641 17003 21644
rect 16945 21635 17003 21641
rect 17494 21632 17500 21644
rect 17552 21632 17558 21684
rect 20162 21672 20168 21684
rect 20123 21644 20168 21672
rect 20162 21632 20168 21644
rect 20220 21632 20226 21684
rect 23566 21672 23572 21684
rect 22066 21644 23572 21672
rect 12526 21604 12532 21616
rect 12406 21576 12532 21604
rect 12526 21564 12532 21576
rect 12584 21604 12590 21616
rect 17954 21604 17960 21616
rect 12584 21576 17960 21604
rect 12584 21564 12590 21576
rect 17954 21564 17960 21576
rect 18012 21564 18018 21616
rect 21910 21604 21916 21616
rect 18064 21576 21916 21604
rect 1762 21536 1768 21548
rect 1723 21508 1768 21536
rect 1762 21496 1768 21508
rect 1820 21496 1826 21548
rect 12268 21536 12296 21564
rect 13538 21536 13544 21548
rect 12268 21508 13544 21536
rect 13538 21496 13544 21508
rect 13596 21496 13602 21548
rect 13814 21536 13820 21548
rect 13775 21508 13820 21536
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 14458 21536 14464 21548
rect 14419 21508 14464 21536
rect 14458 21496 14464 21508
rect 14516 21536 14522 21548
rect 14826 21536 14832 21548
rect 14516 21508 14832 21536
rect 14516 21496 14522 21508
rect 14826 21496 14832 21508
rect 14884 21496 14890 21548
rect 16853 21539 16911 21545
rect 16853 21505 16865 21539
rect 16899 21536 16911 21539
rect 17310 21536 17316 21548
rect 16899 21508 17316 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 17310 21496 17316 21508
rect 17368 21496 17374 21548
rect 18064 21536 18092 21576
rect 21910 21564 21916 21576
rect 21968 21564 21974 21616
rect 22066 21604 22094 21644
rect 23566 21632 23572 21644
rect 23624 21632 23630 21684
rect 24210 21672 24216 21684
rect 24171 21644 24216 21672
rect 24210 21632 24216 21644
rect 24268 21632 24274 21684
rect 29546 21672 29552 21684
rect 29507 21644 29552 21672
rect 29546 21632 29552 21644
rect 29604 21632 29610 21684
rect 22186 21604 22192 21616
rect 22020 21576 22094 21604
rect 22147 21576 22192 21604
rect 20070 21536 20076 21548
rect 17420 21508 18092 21536
rect 20031 21508 20076 21536
rect 4614 21428 4620 21480
rect 4672 21468 4678 21480
rect 6546 21468 6552 21480
rect 4672 21440 6552 21468
rect 4672 21428 4678 21440
rect 6546 21428 6552 21440
rect 6604 21428 6610 21480
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6656 21440 6837 21468
rect 6270 21360 6276 21412
rect 6328 21400 6334 21412
rect 6656 21400 6684 21440
rect 6825 21437 6837 21440
rect 6871 21468 6883 21471
rect 8297 21471 8355 21477
rect 6871 21440 8064 21468
rect 6871 21437 6883 21440
rect 6825 21431 6883 21437
rect 6328 21372 6684 21400
rect 8036 21400 8064 21440
rect 8297 21437 8309 21471
rect 8343 21468 8355 21471
rect 9398 21468 9404 21480
rect 8343 21440 9404 21468
rect 8343 21437 8355 21440
rect 8297 21431 8355 21437
rect 9398 21428 9404 21440
rect 9456 21468 9462 21480
rect 17420 21468 17448 21508
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 9456 21440 17448 21468
rect 9456 21428 9462 21440
rect 17862 21428 17868 21480
rect 17920 21468 17926 21480
rect 18233 21471 18291 21477
rect 18233 21468 18245 21471
rect 17920 21440 18245 21468
rect 17920 21428 17926 21440
rect 18233 21437 18245 21440
rect 18279 21437 18291 21471
rect 18233 21431 18291 21437
rect 18417 21471 18475 21477
rect 18417 21437 18429 21471
rect 18463 21468 18475 21471
rect 20438 21468 20444 21480
rect 18463 21440 20444 21468
rect 18463 21437 18475 21440
rect 18417 21431 18475 21437
rect 20438 21428 20444 21440
rect 20496 21428 20502 21480
rect 22020 21468 22048 21576
rect 22186 21564 22192 21576
rect 22244 21564 22250 21616
rect 22281 21607 22339 21613
rect 22281 21573 22293 21607
rect 22327 21604 22339 21607
rect 22830 21604 22836 21616
rect 22327 21576 22836 21604
rect 22327 21573 22339 21576
rect 22281 21567 22339 21573
rect 22830 21564 22836 21576
rect 22888 21564 22894 21616
rect 24397 21539 24455 21545
rect 24397 21505 24409 21539
rect 24443 21505 24455 21539
rect 24397 21499 24455 21505
rect 20548 21440 22048 21468
rect 8665 21403 8723 21409
rect 8665 21400 8677 21403
rect 8036 21372 8677 21400
rect 6328 21360 6334 21372
rect 8665 21369 8677 21372
rect 8711 21400 8723 21403
rect 17126 21400 17132 21412
rect 8711 21372 17132 21400
rect 8711 21369 8723 21372
rect 8665 21363 8723 21369
rect 17126 21360 17132 21372
rect 17184 21360 17190 21412
rect 20548 21400 20576 21440
rect 22370 21428 22376 21480
rect 22428 21468 22434 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22428 21440 22477 21468
rect 22428 21428 22434 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 17236 21372 20576 21400
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 2406 21332 2412 21344
rect 1627 21304 2412 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 2406 21292 2412 21304
rect 2464 21292 2470 21344
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 7466 21332 7472 21344
rect 2832 21304 7472 21332
rect 2832 21292 2838 21304
rect 7466 21292 7472 21304
rect 7524 21292 7530 21344
rect 13906 21332 13912 21344
rect 13867 21304 13912 21332
rect 13906 21292 13912 21304
rect 13964 21292 13970 21344
rect 14642 21292 14648 21344
rect 14700 21332 14706 21344
rect 17236 21332 17264 21372
rect 21082 21360 21088 21412
rect 21140 21400 21146 21412
rect 24412 21400 24440 21499
rect 27522 21496 27528 21548
rect 27580 21536 27586 21548
rect 28261 21539 28319 21545
rect 28261 21536 28273 21539
rect 27580 21508 28273 21536
rect 27580 21496 27586 21508
rect 28261 21505 28273 21508
rect 28307 21505 28319 21539
rect 28261 21499 28319 21505
rect 28353 21539 28411 21545
rect 28353 21505 28365 21539
rect 28399 21536 28411 21539
rect 29089 21539 29147 21545
rect 29089 21536 29101 21539
rect 28399 21508 29101 21536
rect 28399 21505 28411 21508
rect 28353 21499 28411 21505
rect 29089 21505 29101 21508
rect 29135 21505 29147 21539
rect 29089 21499 29147 21505
rect 31205 21539 31263 21545
rect 31205 21505 31217 21539
rect 31251 21536 31263 21539
rect 33042 21536 33048 21548
rect 31251 21508 33048 21536
rect 31251 21505 31263 21508
rect 31205 21499 31263 21505
rect 33042 21496 33048 21508
rect 33100 21496 33106 21548
rect 28905 21471 28963 21477
rect 28905 21437 28917 21471
rect 28951 21468 28963 21471
rect 31297 21471 31355 21477
rect 31297 21468 31309 21471
rect 28951 21440 31309 21468
rect 28951 21437 28963 21440
rect 28905 21431 28963 21437
rect 31297 21437 31309 21440
rect 31343 21437 31355 21471
rect 31297 21431 31355 21437
rect 21140 21372 24440 21400
rect 21140 21360 21146 21372
rect 14700 21304 17264 21332
rect 18877 21335 18935 21341
rect 14700 21292 14706 21304
rect 18877 21301 18889 21335
rect 18923 21332 18935 21335
rect 19242 21332 19248 21344
rect 18923 21304 19248 21332
rect 18923 21301 18935 21304
rect 18877 21295 18935 21301
rect 19242 21292 19248 21304
rect 19300 21292 19306 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 4236 21131 4294 21137
rect 4236 21097 4248 21131
rect 4282 21128 4294 21131
rect 6086 21128 6092 21140
rect 4282 21100 6092 21128
rect 4282 21097 4294 21100
rect 4236 21091 4294 21097
rect 6086 21088 6092 21100
rect 6144 21088 6150 21140
rect 12069 21131 12127 21137
rect 12069 21097 12081 21131
rect 12115 21128 12127 21131
rect 12158 21128 12164 21140
rect 12115 21100 12164 21128
rect 12115 21097 12127 21100
rect 12069 21091 12127 21097
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 14918 21088 14924 21140
rect 14976 21128 14982 21140
rect 16390 21128 16396 21140
rect 14976 21100 16396 21128
rect 14976 21088 14982 21100
rect 16390 21088 16396 21100
rect 16448 21128 16454 21140
rect 21542 21128 21548 21140
rect 16448 21100 21548 21128
rect 16448 21088 16454 21100
rect 21542 21088 21548 21100
rect 21600 21088 21606 21140
rect 22830 21128 22836 21140
rect 22791 21100 22836 21128
rect 22830 21088 22836 21100
rect 22888 21088 22894 21140
rect 28442 21088 28448 21140
rect 28500 21128 28506 21140
rect 29733 21131 29791 21137
rect 29733 21128 29745 21131
rect 28500 21100 29745 21128
rect 28500 21088 28506 21100
rect 29733 21097 29745 21100
rect 29779 21097 29791 21131
rect 30926 21128 30932 21140
rect 30887 21100 30932 21128
rect 29733 21091 29791 21097
rect 30926 21088 30932 21100
rect 30984 21088 30990 21140
rect 16761 21063 16819 21069
rect 16761 21029 16773 21063
rect 16807 21029 16819 21063
rect 16761 21023 16819 21029
rect 2774 20952 2780 21004
rect 2832 20992 2838 21004
rect 3970 20992 3976 21004
rect 2832 20964 2877 20992
rect 3883 20964 3976 20992
rect 2832 20952 2838 20964
rect 3970 20952 3976 20964
rect 4028 20992 4034 21004
rect 4614 20992 4620 21004
rect 4028 20964 4620 20992
rect 4028 20952 4034 20964
rect 4614 20952 4620 20964
rect 4672 20952 4678 21004
rect 10597 20995 10655 21001
rect 10597 20961 10609 20995
rect 10643 20992 10655 20995
rect 14090 20992 14096 21004
rect 10643 20964 14096 20992
rect 10643 20961 10655 20964
rect 10597 20955 10655 20961
rect 14090 20952 14096 20964
rect 14148 20952 14154 21004
rect 16776 20992 16804 21023
rect 17126 21020 17132 21072
rect 17184 21060 17190 21072
rect 23014 21060 23020 21072
rect 17184 21032 23020 21060
rect 17184 21020 17190 21032
rect 23014 21020 23020 21032
rect 23072 21020 23078 21072
rect 28537 21063 28595 21069
rect 28537 21029 28549 21063
rect 28583 21060 28595 21063
rect 29546 21060 29552 21072
rect 28583 21032 29552 21060
rect 28583 21029 28595 21032
rect 28537 21023 28595 21029
rect 29546 21020 29552 21032
rect 29604 21020 29610 21072
rect 15672 20964 16804 20992
rect 17865 20995 17923 21001
rect 9490 20884 9496 20936
rect 9548 20924 9554 20936
rect 10321 20927 10379 20933
rect 10321 20924 10333 20927
rect 9548 20896 10333 20924
rect 9548 20884 9554 20896
rect 10321 20893 10333 20896
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20924 14887 20927
rect 15286 20924 15292 20936
rect 14875 20896 15292 20924
rect 14875 20893 14887 20896
rect 14829 20887 14887 20893
rect 15286 20884 15292 20896
rect 15344 20924 15350 20936
rect 15470 20924 15476 20936
rect 15344 20896 15476 20924
rect 15344 20884 15350 20896
rect 15470 20884 15476 20896
rect 15528 20884 15534 20936
rect 15672 20933 15700 20964
rect 17865 20961 17877 20995
rect 17911 20992 17923 20995
rect 18414 20992 18420 21004
rect 17911 20964 18420 20992
rect 17911 20961 17923 20964
rect 17865 20955 17923 20961
rect 18414 20952 18420 20964
rect 18472 20952 18478 21004
rect 20714 20952 20720 21004
rect 20772 20992 20778 21004
rect 21269 20995 21327 21001
rect 21269 20992 21281 20995
rect 20772 20964 21281 20992
rect 20772 20952 20778 20964
rect 21269 20961 21281 20964
rect 21315 20961 21327 20995
rect 27893 20995 27951 21001
rect 27893 20992 27905 20995
rect 21269 20955 21327 20961
rect 22066 20964 27905 20992
rect 15657 20927 15715 20933
rect 15657 20893 15669 20927
rect 15703 20893 15715 20927
rect 16114 20924 16120 20936
rect 16075 20896 16120 20924
rect 15657 20887 15715 20893
rect 16114 20884 16120 20896
rect 16172 20884 16178 20936
rect 16945 20927 17003 20933
rect 16945 20893 16957 20927
rect 16991 20924 17003 20927
rect 17678 20924 17684 20936
rect 16991 20896 17684 20924
rect 16991 20893 17003 20896
rect 16945 20887 17003 20893
rect 17678 20884 17684 20896
rect 17736 20884 17742 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19392 20896 19809 20924
rect 19392 20884 19398 20896
rect 19797 20893 19809 20896
rect 19843 20893 19855 20927
rect 21450 20924 21456 20936
rect 21411 20896 21456 20924
rect 19797 20887 19855 20893
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 2869 20859 2927 20865
rect 2869 20825 2881 20859
rect 2915 20825 2927 20859
rect 3418 20856 3424 20868
rect 3379 20828 3424 20856
rect 2869 20819 2927 20825
rect 2884 20788 2912 20819
rect 3418 20816 3424 20828
rect 3476 20816 3482 20868
rect 4706 20816 4712 20868
rect 4764 20816 4770 20868
rect 9674 20816 9680 20868
rect 9732 20856 9738 20868
rect 16209 20859 16267 20865
rect 9732 20828 11086 20856
rect 9732 20816 9738 20828
rect 16209 20825 16221 20859
rect 16255 20856 16267 20859
rect 17957 20859 18015 20865
rect 16255 20828 17816 20856
rect 16255 20825 16267 20828
rect 16209 20819 16267 20825
rect 5626 20788 5632 20800
rect 2884 20760 5632 20788
rect 5626 20748 5632 20760
rect 5684 20748 5690 20800
rect 5721 20791 5779 20797
rect 5721 20757 5733 20791
rect 5767 20788 5779 20791
rect 7926 20788 7932 20800
rect 5767 20760 7932 20788
rect 5767 20757 5779 20760
rect 5721 20751 5779 20757
rect 7926 20748 7932 20760
rect 7984 20748 7990 20800
rect 13446 20748 13452 20800
rect 13504 20788 13510 20800
rect 14921 20791 14979 20797
rect 14921 20788 14933 20791
rect 13504 20760 14933 20788
rect 13504 20748 13510 20760
rect 14921 20757 14933 20760
rect 14967 20757 14979 20791
rect 14921 20751 14979 20757
rect 15473 20791 15531 20797
rect 15473 20757 15485 20791
rect 15519 20788 15531 20791
rect 16482 20788 16488 20800
rect 15519 20760 16488 20788
rect 15519 20757 15531 20760
rect 15473 20751 15531 20757
rect 16482 20748 16488 20760
rect 16540 20748 16546 20800
rect 17788 20788 17816 20828
rect 17957 20825 17969 20859
rect 18003 20825 18015 20859
rect 17957 20819 18015 20825
rect 17972 20788 18000 20819
rect 18506 20816 18512 20868
rect 18564 20856 18570 20868
rect 18782 20856 18788 20868
rect 18564 20828 18788 20856
rect 18564 20816 18570 20828
rect 18782 20816 18788 20828
rect 18840 20856 18846 20868
rect 18877 20859 18935 20865
rect 18877 20856 18889 20859
rect 18840 20828 18889 20856
rect 18840 20816 18846 20828
rect 18877 20825 18889 20828
rect 18923 20825 18935 20859
rect 22066 20856 22094 20964
rect 27893 20961 27905 20964
rect 27939 20992 27951 20995
rect 27982 20992 27988 21004
rect 27939 20964 27988 20992
rect 27939 20961 27951 20964
rect 27893 20955 27951 20961
rect 27982 20952 27988 20964
rect 28040 20952 28046 21004
rect 23014 20924 23020 20936
rect 22975 20896 23020 20924
rect 23014 20884 23020 20896
rect 23072 20884 23078 20936
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20924 23535 20927
rect 24762 20924 24768 20936
rect 23523 20896 24768 20924
rect 23523 20893 23535 20896
rect 23477 20887 23535 20893
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 27433 20927 27491 20933
rect 27433 20893 27445 20927
rect 27479 20924 27491 20927
rect 27522 20924 27528 20936
rect 27479 20896 27528 20924
rect 27479 20893 27491 20896
rect 27433 20887 27491 20893
rect 27522 20884 27528 20896
rect 27580 20884 27586 20936
rect 28074 20924 28080 20936
rect 28035 20896 28080 20924
rect 28074 20884 28080 20896
rect 28132 20884 28138 20936
rect 29914 20924 29920 20936
rect 29875 20896 29920 20924
rect 29914 20884 29920 20896
rect 29972 20884 29978 20936
rect 31110 20924 31116 20936
rect 31071 20896 31116 20924
rect 31110 20884 31116 20896
rect 31168 20884 31174 20936
rect 18877 20819 18935 20825
rect 19260 20828 22094 20856
rect 17788 20760 18000 20788
rect 18046 20748 18052 20800
rect 18104 20788 18110 20800
rect 19260 20788 19288 20828
rect 18104 20760 19288 20788
rect 18104 20748 18110 20760
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 19392 20760 19625 20788
rect 19392 20748 19398 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 19613 20751 19671 20757
rect 21913 20791 21971 20797
rect 21913 20757 21925 20791
rect 21959 20788 21971 20791
rect 23198 20788 23204 20800
rect 21959 20760 23204 20788
rect 21959 20757 21971 20760
rect 21913 20751 21971 20757
rect 23198 20748 23204 20760
rect 23256 20748 23262 20800
rect 23566 20788 23572 20800
rect 23527 20760 23572 20788
rect 23566 20748 23572 20760
rect 23624 20748 23630 20800
rect 27249 20791 27307 20797
rect 27249 20757 27261 20791
rect 27295 20788 27307 20791
rect 27890 20788 27896 20800
rect 27295 20760 27896 20788
rect 27295 20757 27307 20760
rect 27249 20751 27307 20757
rect 27890 20748 27896 20760
rect 27948 20748 27954 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1578 20544 1584 20596
rect 1636 20584 1642 20596
rect 1765 20587 1823 20593
rect 1765 20584 1777 20587
rect 1636 20556 1777 20584
rect 1636 20544 1642 20556
rect 1765 20553 1777 20556
rect 1811 20553 1823 20587
rect 1765 20547 1823 20553
rect 14645 20587 14703 20593
rect 14645 20553 14657 20587
rect 14691 20584 14703 20587
rect 14734 20584 14740 20596
rect 14691 20556 14740 20584
rect 14691 20553 14703 20556
rect 14645 20547 14703 20553
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 16022 20584 16028 20596
rect 15488 20556 16028 20584
rect 7561 20519 7619 20525
rect 7561 20485 7573 20519
rect 7607 20516 7619 20519
rect 7834 20516 7840 20528
rect 7607 20488 7840 20516
rect 7607 20485 7619 20488
rect 7561 20479 7619 20485
rect 7834 20476 7840 20488
rect 7892 20476 7898 20528
rect 13446 20516 13452 20528
rect 8786 20488 13452 20516
rect 13446 20476 13452 20488
rect 13504 20476 13510 20528
rect 1946 20448 1952 20460
rect 1907 20420 1952 20448
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 4614 20408 4620 20460
rect 4672 20448 4678 20460
rect 7285 20451 7343 20457
rect 7285 20448 7297 20451
rect 4672 20420 7297 20448
rect 4672 20408 4678 20420
rect 7285 20417 7297 20420
rect 7331 20417 7343 20451
rect 7285 20411 7343 20417
rect 14182 20408 14188 20460
rect 14240 20408 14246 20460
rect 15194 20448 15200 20460
rect 14306 20420 15200 20448
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15488 20457 15516 20556
rect 16022 20544 16028 20556
rect 16080 20584 16086 20596
rect 16298 20584 16304 20596
rect 16080 20556 16304 20584
rect 16080 20544 16086 20556
rect 16298 20544 16304 20556
rect 16356 20544 16362 20596
rect 20438 20584 20444 20596
rect 20399 20556 20444 20584
rect 20438 20544 20444 20556
rect 20496 20544 20502 20596
rect 21450 20544 21456 20596
rect 21508 20584 21514 20596
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 21508 20556 22017 20584
rect 21508 20544 21514 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 22005 20547 22063 20553
rect 27709 20587 27767 20593
rect 27709 20553 27721 20587
rect 27755 20584 27767 20587
rect 28074 20584 28080 20596
rect 27755 20556 28080 20584
rect 27755 20553 27767 20556
rect 27709 20547 27767 20553
rect 28074 20544 28080 20556
rect 28132 20544 28138 20596
rect 29273 20587 29331 20593
rect 29273 20553 29285 20587
rect 29319 20584 29331 20587
rect 29914 20584 29920 20596
rect 29319 20556 29920 20584
rect 29319 20553 29331 20556
rect 29273 20547 29331 20553
rect 29914 20544 29920 20556
rect 29972 20544 29978 20596
rect 31110 20584 31116 20596
rect 31071 20556 31116 20584
rect 31110 20544 31116 20556
rect 31168 20544 31174 20596
rect 16209 20519 16267 20525
rect 16209 20485 16221 20519
rect 16255 20516 16267 20519
rect 17037 20519 17095 20525
rect 17037 20516 17049 20519
rect 16255 20488 17049 20516
rect 16255 20485 16267 20488
rect 16209 20479 16267 20485
rect 17037 20485 17049 20488
rect 17083 20485 17095 20519
rect 19334 20516 19340 20528
rect 19295 20488 19340 20516
rect 17037 20479 17095 20485
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20417 15531 20451
rect 16114 20448 16120 20460
rect 16075 20420 16120 20448
rect 15473 20411 15531 20417
rect 16114 20408 16120 20420
rect 16172 20408 16178 20460
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20448 18107 20451
rect 18230 20448 18236 20460
rect 18095 20420 18236 20448
rect 18095 20417 18107 20420
rect 18049 20411 18107 20417
rect 18230 20408 18236 20420
rect 18288 20408 18294 20460
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 9306 20380 9312 20392
rect 9267 20352 9312 20380
rect 9306 20340 9312 20352
rect 9364 20340 9370 20392
rect 12894 20380 12900 20392
rect 12855 20352 12900 20380
rect 12894 20340 12900 20352
rect 12952 20340 12958 20392
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 14200 20380 14228 20408
rect 15562 20380 15568 20392
rect 13219 20352 14228 20380
rect 14660 20352 15568 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 3970 20204 3976 20256
rect 4028 20244 4034 20256
rect 14660 20244 14688 20352
rect 15562 20340 15568 20352
rect 15620 20380 15626 20392
rect 15930 20380 15936 20392
rect 15620 20352 15936 20380
rect 15620 20340 15626 20352
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 16942 20380 16948 20392
rect 16903 20352 16948 20380
rect 16942 20340 16948 20352
rect 17000 20340 17006 20392
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 17052 20352 17233 20380
rect 15562 20244 15568 20256
rect 4028 20216 14688 20244
rect 15523 20216 15568 20244
rect 4028 20204 4034 20216
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 16942 20204 16948 20256
rect 17000 20244 17006 20256
rect 17052 20244 17080 20352
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 19242 20380 19248 20392
rect 19203 20352 19248 20380
rect 17221 20343 17279 20349
rect 19242 20340 19248 20352
rect 19300 20340 19306 20392
rect 19889 20383 19947 20389
rect 19889 20349 19901 20383
rect 19935 20380 19947 20383
rect 19978 20380 19984 20392
rect 19935 20352 19984 20380
rect 19935 20349 19947 20352
rect 19889 20343 19947 20349
rect 19978 20340 19984 20352
rect 20036 20340 20042 20392
rect 20364 20380 20392 20411
rect 21910 20408 21916 20460
rect 21968 20448 21974 20460
rect 22189 20451 22247 20457
rect 22189 20448 22201 20451
rect 21968 20420 22201 20448
rect 21968 20408 21974 20420
rect 22189 20417 22201 20420
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 23293 20451 23351 20457
rect 23293 20417 23305 20451
rect 23339 20448 23351 20451
rect 23566 20448 23572 20460
rect 23339 20420 23572 20448
rect 23339 20417 23351 20420
rect 23293 20411 23351 20417
rect 23566 20408 23572 20420
rect 23624 20408 23630 20460
rect 27890 20448 27896 20460
rect 27851 20420 27896 20448
rect 27890 20408 27896 20420
rect 27948 20408 27954 20460
rect 29454 20448 29460 20460
rect 29415 20420 29460 20448
rect 29454 20408 29460 20420
rect 29512 20408 29518 20460
rect 29917 20451 29975 20457
rect 29917 20417 29929 20451
rect 29963 20448 29975 20451
rect 30190 20448 30196 20460
rect 29963 20420 30196 20448
rect 29963 20417 29975 20420
rect 29917 20411 29975 20417
rect 30190 20408 30196 20420
rect 30248 20408 30254 20460
rect 31018 20448 31024 20460
rect 30979 20420 31024 20448
rect 31018 20408 31024 20420
rect 31076 20408 31082 20460
rect 32953 20451 33011 20457
rect 32953 20417 32965 20451
rect 32999 20448 33011 20451
rect 36446 20448 36452 20460
rect 32999 20420 36452 20448
rect 32999 20417 33011 20420
rect 32953 20411 33011 20417
rect 36446 20408 36452 20420
rect 36504 20408 36510 20460
rect 22738 20380 22744 20392
rect 20364 20352 22744 20380
rect 17402 20272 17408 20324
rect 17460 20312 17466 20324
rect 20364 20312 20392 20352
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 23106 20380 23112 20392
rect 23067 20352 23112 20380
rect 23106 20340 23112 20352
rect 23164 20340 23170 20392
rect 30101 20383 30159 20389
rect 30101 20349 30113 20383
rect 30147 20380 30159 20383
rect 30374 20380 30380 20392
rect 30147 20352 30380 20380
rect 30147 20349 30159 20352
rect 30101 20343 30159 20349
rect 30374 20340 30380 20352
rect 30432 20340 30438 20392
rect 17460 20284 20392 20312
rect 17460 20272 17466 20284
rect 17000 20216 17080 20244
rect 17000 20204 17006 20216
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 18141 20247 18199 20253
rect 18141 20244 18153 20247
rect 18012 20216 18153 20244
rect 18012 20204 18018 20216
rect 18141 20213 18153 20216
rect 18187 20213 18199 20247
rect 18141 20207 18199 20213
rect 22830 20204 22836 20256
rect 22888 20244 22894 20256
rect 23477 20247 23535 20253
rect 23477 20244 23489 20247
rect 22888 20216 23489 20244
rect 22888 20204 22894 20216
rect 23477 20213 23489 20216
rect 23523 20213 23535 20247
rect 30466 20244 30472 20256
rect 30427 20216 30472 20244
rect 23477 20207 23535 20213
rect 30466 20204 30472 20216
rect 30524 20204 30530 20256
rect 31754 20204 31760 20256
rect 31812 20244 31818 20256
rect 32769 20247 32827 20253
rect 32769 20244 32781 20247
rect 31812 20216 32781 20244
rect 31812 20204 31818 20216
rect 32769 20213 32781 20216
rect 32815 20213 32827 20247
rect 32769 20207 32827 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 2866 20040 2872 20052
rect 1627 20012 2872 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 5828 20012 10811 20040
rect 1762 19836 1768 19848
rect 1723 19808 1768 19836
rect 1762 19796 1768 19808
rect 1820 19796 1826 19848
rect 2222 19796 2228 19848
rect 2280 19836 2286 19848
rect 4433 19839 4491 19845
rect 4433 19836 4445 19839
rect 2280 19808 4445 19836
rect 2280 19796 2286 19808
rect 4433 19805 4445 19808
rect 4479 19805 4491 19839
rect 5828 19822 5856 20012
rect 10783 19972 10811 20012
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11241 20043 11299 20049
rect 11241 20040 11253 20043
rect 11112 20012 11253 20040
rect 11112 20000 11118 20012
rect 11241 20009 11253 20012
rect 11287 20009 11299 20043
rect 13906 20040 13912 20052
rect 11241 20003 11299 20009
rect 11348 20012 13912 20040
rect 11348 19972 11376 20012
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 15194 20040 15200 20052
rect 15155 20012 15200 20040
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 17218 20000 17224 20052
rect 17276 20040 17282 20052
rect 17773 20043 17831 20049
rect 17773 20040 17785 20043
rect 17276 20012 17785 20040
rect 17276 20000 17282 20012
rect 17773 20009 17785 20012
rect 17819 20009 17831 20043
rect 21910 20040 21916 20052
rect 21871 20012 21916 20040
rect 17773 20003 17831 20009
rect 21910 20000 21916 20012
rect 21968 20000 21974 20052
rect 23014 20000 23020 20052
rect 23072 20040 23078 20052
rect 23201 20043 23259 20049
rect 23201 20040 23213 20043
rect 23072 20012 23213 20040
rect 23072 20000 23078 20012
rect 23201 20009 23213 20012
rect 23247 20009 23259 20043
rect 28166 20040 28172 20052
rect 23201 20003 23259 20009
rect 24596 20012 28172 20040
rect 10783 19944 11376 19972
rect 11422 19932 11428 19984
rect 11480 19972 11486 19984
rect 15654 19972 15660 19984
rect 11480 19944 15660 19972
rect 11480 19932 11486 19944
rect 15654 19932 15660 19944
rect 15712 19932 15718 19984
rect 9490 19904 9496 19916
rect 9451 19876 9496 19904
rect 9490 19864 9496 19876
rect 9548 19864 9554 19916
rect 9769 19907 9827 19913
rect 9769 19873 9781 19907
rect 9815 19904 9827 19907
rect 14918 19904 14924 19916
rect 9815 19876 14924 19904
rect 9815 19873 9827 19876
rect 9769 19867 9827 19873
rect 14918 19864 14924 19876
rect 14976 19864 14982 19916
rect 23106 19904 23112 19916
rect 15028 19876 23112 19904
rect 7653 19839 7711 19845
rect 4433 19799 4491 19805
rect 7653 19805 7665 19839
rect 7699 19836 7711 19839
rect 7926 19836 7932 19848
rect 7699 19808 7932 19836
rect 7699 19805 7711 19808
rect 7653 19799 7711 19805
rect 4448 19768 4476 19799
rect 7926 19796 7932 19808
rect 7984 19796 7990 19848
rect 11514 19796 11520 19848
rect 11572 19836 11578 19848
rect 15028 19836 15056 19876
rect 23106 19864 23112 19876
rect 23164 19864 23170 19916
rect 24596 19913 24624 20012
rect 28166 20000 28172 20012
rect 28224 20000 28230 20052
rect 30374 20040 30380 20052
rect 30335 20012 30380 20040
rect 30374 20000 30380 20012
rect 30432 20000 30438 20052
rect 33042 20000 33048 20052
rect 33100 20040 33106 20052
rect 38105 20043 38163 20049
rect 38105 20040 38117 20043
rect 33100 20012 38117 20040
rect 33100 20000 33106 20012
rect 38105 20009 38117 20012
rect 38151 20009 38163 20043
rect 38105 20003 38163 20009
rect 25685 19975 25743 19981
rect 25685 19941 25697 19975
rect 25731 19972 25743 19975
rect 25731 19944 26234 19972
rect 25731 19941 25743 19944
rect 25685 19935 25743 19941
rect 24581 19907 24639 19913
rect 24581 19873 24593 19907
rect 24627 19873 24639 19907
rect 24581 19867 24639 19873
rect 11572 19808 15056 19836
rect 15105 19839 15163 19845
rect 11572 19796 11578 19808
rect 15105 19805 15117 19839
rect 15151 19805 15163 19839
rect 15105 19799 15163 19805
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19836 17739 19839
rect 17770 19836 17776 19848
rect 17727 19808 17776 19836
rect 17727 19805 17739 19808
rect 17681 19799 17739 19805
rect 4614 19768 4620 19780
rect 4448 19740 4620 19768
rect 4614 19728 4620 19740
rect 4672 19728 4678 19780
rect 4709 19771 4767 19777
rect 4709 19737 4721 19771
rect 4755 19737 4767 19771
rect 6454 19768 6460 19780
rect 6415 19740 6460 19768
rect 4709 19731 4767 19737
rect 4724 19700 4752 19731
rect 6454 19728 6460 19740
rect 6512 19728 6518 19780
rect 11146 19768 11152 19780
rect 10994 19740 11152 19768
rect 11146 19728 11152 19740
rect 11204 19728 11210 19780
rect 14366 19728 14372 19780
rect 14424 19768 14430 19780
rect 15010 19768 15016 19780
rect 14424 19740 15016 19768
rect 14424 19728 14430 19740
rect 15010 19728 15016 19740
rect 15068 19768 15074 19780
rect 15120 19768 15148 19799
rect 17770 19796 17776 19808
rect 17828 19796 17834 19848
rect 22097 19839 22155 19845
rect 22097 19805 22109 19839
rect 22143 19836 22155 19839
rect 22554 19836 22560 19848
rect 22143 19808 22560 19836
rect 22143 19805 22155 19808
rect 22097 19799 22155 19805
rect 22554 19796 22560 19808
rect 22612 19796 22618 19848
rect 22738 19836 22744 19848
rect 22699 19808 22744 19836
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 23290 19796 23296 19848
rect 23348 19836 23354 19848
rect 23385 19839 23443 19845
rect 23385 19836 23397 19839
rect 23348 19808 23397 19836
rect 23348 19796 23354 19808
rect 23385 19805 23397 19808
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19836 24823 19839
rect 25314 19836 25320 19848
rect 24811 19808 25320 19836
rect 24811 19805 24823 19808
rect 24765 19799 24823 19805
rect 25314 19796 25320 19808
rect 25372 19796 25378 19848
rect 25866 19836 25872 19848
rect 25827 19808 25872 19836
rect 25866 19796 25872 19808
rect 25924 19796 25930 19848
rect 26206 19836 26234 19944
rect 28261 19907 28319 19913
rect 28261 19873 28273 19907
rect 28307 19904 28319 19907
rect 28626 19904 28632 19916
rect 28307 19876 28632 19904
rect 28307 19873 28319 19876
rect 28261 19867 28319 19873
rect 28626 19864 28632 19876
rect 28684 19864 28690 19916
rect 28902 19904 28908 19916
rect 28863 19876 28908 19904
rect 28902 19864 28908 19876
rect 28960 19864 28966 19916
rect 26513 19839 26571 19845
rect 26513 19836 26525 19839
rect 26206 19808 26525 19836
rect 26513 19805 26525 19808
rect 26559 19805 26571 19839
rect 30282 19836 30288 19848
rect 30243 19808 30288 19836
rect 26513 19799 26571 19805
rect 30282 19796 30288 19808
rect 30340 19796 30346 19848
rect 38286 19836 38292 19848
rect 38247 19808 38292 19836
rect 38286 19796 38292 19808
rect 38344 19796 38350 19848
rect 15068 19740 15148 19768
rect 15068 19728 15074 19740
rect 28350 19728 28356 19780
rect 28408 19768 28414 19780
rect 28408 19740 28453 19768
rect 28408 19728 28414 19740
rect 5534 19700 5540 19712
rect 4724 19672 5540 19700
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 5626 19660 5632 19712
rect 5684 19700 5690 19712
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 5684 19672 7757 19700
rect 5684 19660 5690 19672
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 11701 19703 11759 19709
rect 11701 19669 11713 19703
rect 11747 19700 11759 19703
rect 11790 19700 11796 19712
rect 11747 19672 11796 19700
rect 11747 19669 11759 19672
rect 11701 19663 11759 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 22554 19700 22560 19712
rect 22515 19672 22560 19700
rect 22554 19660 22560 19672
rect 22612 19660 22618 19712
rect 25225 19703 25283 19709
rect 25225 19669 25237 19703
rect 25271 19700 25283 19703
rect 25406 19700 25412 19712
rect 25271 19672 25412 19700
rect 25271 19669 25283 19672
rect 25225 19663 25283 19669
rect 25406 19660 25412 19672
rect 25464 19660 25470 19712
rect 26326 19700 26332 19712
rect 26287 19672 26332 19700
rect 26326 19660 26332 19672
rect 26384 19660 26390 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 3970 19496 3976 19508
rect 3931 19468 3976 19496
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 10778 19456 10784 19508
rect 10836 19496 10842 19508
rect 10836 19468 13492 19496
rect 10836 19456 10842 19468
rect 11422 19428 11428 19440
rect 3726 19400 11428 19428
rect 11422 19388 11428 19400
rect 11480 19388 11486 19440
rect 11790 19428 11796 19440
rect 11751 19400 11796 19428
rect 11790 19388 11796 19400
rect 11848 19388 11854 19440
rect 11885 19431 11943 19437
rect 11885 19397 11897 19431
rect 11931 19428 11943 19431
rect 13354 19428 13360 19440
rect 11931 19400 13360 19428
rect 11931 19397 11943 19400
rect 11885 19391 11943 19397
rect 13354 19388 13360 19400
rect 13412 19388 13418 19440
rect 13464 19428 13492 19468
rect 14090 19456 14096 19508
rect 14148 19496 14154 19508
rect 14148 19468 15240 19496
rect 14148 19456 14154 19468
rect 15212 19437 15240 19468
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 21269 19499 21327 19505
rect 21269 19496 21281 19499
rect 19300 19468 21281 19496
rect 19300 19456 19306 19468
rect 21269 19465 21281 19468
rect 21315 19465 21327 19499
rect 25314 19496 25320 19508
rect 25275 19468 25320 19496
rect 21269 19459 21327 19465
rect 25314 19456 25320 19468
rect 25372 19456 25378 19508
rect 15197 19431 15255 19437
rect 13464 19400 13938 19428
rect 15197 19397 15209 19431
rect 15243 19428 15255 19431
rect 17402 19428 17408 19440
rect 15243 19400 17408 19428
rect 15243 19397 15255 19400
rect 15197 19391 15255 19397
rect 17402 19388 17408 19400
rect 17460 19388 17466 19440
rect 19334 19428 19340 19440
rect 19295 19400 19340 19428
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 27338 19428 27344 19440
rect 27299 19400 27344 19428
rect 27338 19388 27344 19400
rect 27396 19388 27402 19440
rect 22554 19360 22560 19372
rect 22515 19332 22560 19360
rect 22554 19320 22560 19332
rect 22612 19320 22618 19372
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19360 25283 19363
rect 25866 19360 25872 19372
rect 25271 19332 25872 19360
rect 25271 19329 25283 19332
rect 25225 19323 25283 19329
rect 25866 19320 25872 19332
rect 25924 19320 25930 19372
rect 28353 19363 28411 19369
rect 28353 19329 28365 19363
rect 28399 19360 28411 19363
rect 28442 19360 28448 19372
rect 28399 19332 28448 19360
rect 28399 19329 28411 19332
rect 28353 19323 28411 19329
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 28626 19320 28632 19372
rect 28684 19360 28690 19372
rect 28997 19363 29055 19369
rect 28997 19360 29009 19363
rect 28684 19332 29009 19360
rect 28684 19320 28690 19332
rect 28997 19329 29009 19332
rect 29043 19329 29055 19363
rect 28997 19323 29055 19329
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 2498 19292 2504 19304
rect 2459 19264 2504 19292
rect 2498 19252 2504 19264
rect 2556 19292 2562 19304
rect 9306 19292 9312 19304
rect 2556 19264 9312 19292
rect 2556 19252 2562 19264
rect 9306 19252 9312 19264
rect 9364 19252 9370 19304
rect 12250 19292 12256 19304
rect 12211 19264 12256 19292
rect 12250 19252 12256 19264
rect 12308 19252 12314 19304
rect 12406 19264 12848 19292
rect 6730 19184 6736 19236
rect 6788 19224 6794 19236
rect 12406 19224 12434 19264
rect 6788 19196 12434 19224
rect 12820 19224 12848 19264
rect 12894 19252 12900 19304
rect 12952 19292 12958 19304
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 12952 19264 13185 19292
rect 12952 19252 12958 19264
rect 13173 19261 13185 19264
rect 13219 19261 13231 19295
rect 13449 19295 13507 19301
rect 13449 19292 13461 19295
rect 13173 19255 13231 19261
rect 13280 19264 13461 19292
rect 13280 19224 13308 19264
rect 13449 19261 13461 19264
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 13906 19252 13912 19304
rect 13964 19292 13970 19304
rect 16850 19292 16856 19304
rect 13964 19264 14504 19292
rect 16811 19264 16856 19292
rect 13964 19252 13970 19264
rect 12820 19196 13308 19224
rect 14476 19224 14504 19264
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 19245 19295 19303 19301
rect 19245 19261 19257 19295
rect 19291 19292 19303 19295
rect 19426 19292 19432 19304
rect 19291 19264 19432 19292
rect 19291 19261 19303 19264
rect 19245 19255 19303 19261
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 19521 19295 19579 19301
rect 19521 19261 19533 19295
rect 19567 19261 19579 19295
rect 20622 19292 20628 19304
rect 20583 19264 20628 19292
rect 19521 19255 19579 19261
rect 18138 19224 18144 19236
rect 14476 19196 18144 19224
rect 6788 19184 6794 19196
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 16666 19156 16672 19168
rect 8444 19128 16672 19156
rect 8444 19116 8450 19128
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 19536 19156 19564 19255
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 27246 19292 27252 19304
rect 20855 19264 22416 19292
rect 27207 19264 27252 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 22388 19233 22416 19264
rect 27246 19252 27252 19264
rect 27304 19252 27310 19304
rect 28537 19295 28595 19301
rect 28537 19261 28549 19295
rect 28583 19261 28595 19295
rect 28537 19255 28595 19261
rect 22373 19227 22431 19233
rect 22373 19193 22385 19227
rect 22419 19193 22431 19227
rect 27798 19224 27804 19236
rect 27759 19196 27804 19224
rect 22373 19187 22431 19193
rect 27798 19184 27804 19196
rect 27856 19184 27862 19236
rect 27890 19184 27896 19236
rect 27948 19224 27954 19236
rect 28552 19224 28580 19255
rect 27948 19196 28580 19224
rect 27948 19184 27954 19196
rect 19300 19128 19564 19156
rect 19300 19116 19306 19128
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 8294 18952 8300 18964
rect 2746 18924 6684 18952
rect 8255 18924 8300 18952
rect 2406 18748 2412 18760
rect 2367 18720 2412 18748
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 2501 18615 2559 18621
rect 2501 18581 2513 18615
rect 2547 18612 2559 18615
rect 2746 18612 2774 18924
rect 6086 18884 6092 18896
rect 6047 18856 6092 18884
rect 6086 18844 6092 18856
rect 6144 18844 6150 18896
rect 4341 18819 4399 18825
rect 4341 18785 4353 18819
rect 4387 18816 4399 18819
rect 4614 18816 4620 18828
rect 4387 18788 4620 18816
rect 4387 18785 4399 18788
rect 4341 18779 4399 18785
rect 4614 18776 4620 18788
rect 4672 18816 4678 18828
rect 6549 18819 6607 18825
rect 6549 18816 6561 18819
rect 4672 18788 6561 18816
rect 4672 18776 4678 18788
rect 6549 18785 6561 18788
rect 6595 18785 6607 18819
rect 6656 18816 6684 18924
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 9030 18912 9036 18964
rect 9088 18952 9094 18964
rect 9088 18924 15792 18952
rect 9088 18912 9094 18924
rect 13354 18844 13360 18896
rect 13412 18884 13418 18896
rect 15013 18887 15071 18893
rect 15013 18884 15025 18887
rect 13412 18856 15025 18884
rect 13412 18844 13418 18856
rect 15013 18853 15025 18856
rect 15059 18853 15071 18887
rect 15013 18847 15071 18853
rect 15657 18887 15715 18893
rect 15657 18853 15669 18887
rect 15703 18853 15715 18887
rect 15657 18847 15715 18853
rect 13906 18816 13912 18828
rect 6656 18788 13912 18816
rect 6549 18779 6607 18785
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 15672 18816 15700 18847
rect 15212 18788 15700 18816
rect 15764 18816 15792 18924
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19705 18955 19763 18961
rect 19705 18952 19717 18955
rect 19392 18924 19717 18952
rect 19392 18912 19398 18924
rect 19705 18921 19717 18924
rect 19751 18921 19763 18955
rect 26789 18955 26847 18961
rect 19705 18915 19763 18921
rect 19996 18924 26234 18952
rect 16224 18856 18276 18884
rect 15764 18788 15884 18816
rect 10318 18748 10324 18760
rect 10279 18720 10324 18748
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 15212 18757 15240 18788
rect 15856 18757 15884 18788
rect 15197 18751 15255 18757
rect 11730 18720 13860 18748
rect 4617 18683 4675 18689
rect 4617 18649 4629 18683
rect 4663 18680 4675 18683
rect 4663 18652 4752 18680
rect 4663 18649 4675 18652
rect 4617 18643 4675 18649
rect 2547 18584 2774 18612
rect 4724 18612 4752 18652
rect 4890 18640 4896 18692
rect 4948 18680 4954 18692
rect 6822 18680 6828 18692
rect 4948 18652 5106 18680
rect 6783 18652 6828 18680
rect 4948 18640 4954 18652
rect 6822 18640 6828 18652
rect 6880 18640 6886 18692
rect 7558 18640 7564 18692
rect 7616 18640 7622 18692
rect 10597 18683 10655 18689
rect 10597 18649 10609 18683
rect 10643 18680 10655 18683
rect 10870 18680 10876 18692
rect 10643 18652 10876 18680
rect 10643 18649 10655 18652
rect 10597 18643 10655 18649
rect 10870 18640 10876 18652
rect 10928 18640 10934 18692
rect 12342 18680 12348 18692
rect 12303 18652 12348 18680
rect 12342 18640 12348 18652
rect 12400 18640 12406 18692
rect 13832 18680 13860 18720
rect 15197 18717 15209 18751
rect 15243 18717 15255 18751
rect 15197 18711 15255 18717
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 15562 18680 15568 18692
rect 13832 18652 15568 18680
rect 15562 18640 15568 18652
rect 15620 18640 15626 18692
rect 16224 18680 16252 18856
rect 16393 18819 16451 18825
rect 16393 18785 16405 18819
rect 16439 18816 16451 18819
rect 16850 18816 16856 18828
rect 16439 18788 16856 18816
rect 16439 18785 16451 18788
rect 16393 18779 16451 18785
rect 16850 18776 16856 18788
rect 16908 18776 16914 18828
rect 18248 18748 18276 18856
rect 19150 18776 19156 18828
rect 19208 18816 19214 18828
rect 19996 18816 20024 18924
rect 20162 18844 20168 18896
rect 20220 18884 20226 18896
rect 24762 18884 24768 18896
rect 20220 18856 24768 18884
rect 20220 18844 20226 18856
rect 24762 18844 24768 18856
rect 24820 18844 24826 18896
rect 26053 18887 26111 18893
rect 26053 18853 26065 18887
rect 26099 18853 26111 18887
rect 26053 18847 26111 18853
rect 20622 18816 20628 18828
rect 19208 18788 20024 18816
rect 20583 18788 20628 18816
rect 19208 18776 19214 18788
rect 20622 18776 20628 18788
rect 20680 18776 20686 18828
rect 19334 18748 19340 18760
rect 18248 18720 19340 18748
rect 19334 18708 19340 18720
rect 19392 18748 19398 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19392 18720 19625 18748
rect 19392 18708 19398 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 25593 18751 25651 18757
rect 25593 18717 25605 18751
rect 25639 18748 25651 18751
rect 26068 18748 26096 18847
rect 26206 18816 26234 18924
rect 26789 18921 26801 18955
rect 26835 18952 26847 18955
rect 27338 18952 27344 18964
rect 26835 18924 27344 18952
rect 26835 18921 26847 18924
rect 26789 18915 26847 18921
rect 27338 18912 27344 18924
rect 27396 18912 27402 18964
rect 27801 18955 27859 18961
rect 27801 18921 27813 18955
rect 27847 18952 27859 18955
rect 27890 18952 27896 18964
rect 27847 18924 27896 18952
rect 27847 18921 27859 18924
rect 27801 18915 27859 18921
rect 27890 18912 27896 18924
rect 27948 18912 27954 18964
rect 28350 18912 28356 18964
rect 28408 18952 28414 18964
rect 28445 18955 28503 18961
rect 28445 18952 28457 18955
rect 28408 18924 28457 18952
rect 28408 18912 28414 18924
rect 28445 18921 28457 18924
rect 28491 18921 28503 18955
rect 28445 18915 28503 18921
rect 30377 18955 30435 18961
rect 30377 18921 30389 18955
rect 30423 18952 30435 18955
rect 30466 18952 30472 18964
rect 30423 18924 30472 18952
rect 30423 18921 30435 18924
rect 30377 18915 30435 18921
rect 30466 18912 30472 18924
rect 30524 18912 30530 18964
rect 28442 18816 28448 18828
rect 26206 18788 28448 18816
rect 28442 18776 28448 18788
rect 28500 18816 28506 18828
rect 33505 18819 33563 18825
rect 33505 18816 33517 18819
rect 28500 18788 33517 18816
rect 28500 18776 28506 18788
rect 33505 18785 33517 18788
rect 33551 18785 33563 18819
rect 33505 18779 33563 18785
rect 25639 18720 26096 18748
rect 26237 18751 26295 18757
rect 25639 18717 25651 18720
rect 25593 18711 25651 18717
rect 26237 18717 26249 18751
rect 26283 18717 26295 18751
rect 26237 18711 26295 18717
rect 26697 18751 26755 18757
rect 26697 18717 26709 18751
rect 26743 18717 26755 18751
rect 27706 18748 27712 18760
rect 27667 18720 27712 18748
rect 26697 18711 26755 18717
rect 16482 18680 16488 18692
rect 15672 18652 16252 18680
rect 16443 18652 16488 18680
rect 11514 18612 11520 18624
rect 4724 18584 11520 18612
rect 2547 18581 2559 18584
rect 2501 18575 2559 18581
rect 11514 18572 11520 18584
rect 11572 18612 11578 18624
rect 15672 18612 15700 18652
rect 16482 18640 16488 18652
rect 16540 18640 16546 18692
rect 17034 18680 17040 18692
rect 16995 18652 17040 18680
rect 17034 18640 17040 18652
rect 17092 18640 17098 18692
rect 17589 18683 17647 18689
rect 17589 18649 17601 18683
rect 17635 18649 17647 18683
rect 17589 18643 17647 18649
rect 17681 18683 17739 18689
rect 17681 18649 17693 18683
rect 17727 18680 17739 18683
rect 17954 18680 17960 18692
rect 17727 18652 17960 18680
rect 17727 18649 17739 18652
rect 17681 18643 17739 18649
rect 11572 18584 15700 18612
rect 11572 18572 11578 18584
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 17604 18612 17632 18643
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 18233 18683 18291 18689
rect 18233 18649 18245 18683
rect 18279 18680 18291 18683
rect 19426 18680 19432 18692
rect 18279 18652 19432 18680
rect 18279 18649 18291 18652
rect 18233 18643 18291 18649
rect 19426 18640 19432 18652
rect 19484 18680 19490 18692
rect 19978 18680 19984 18692
rect 19484 18652 19984 18680
rect 19484 18640 19490 18652
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 25038 18640 25044 18692
rect 25096 18680 25102 18692
rect 26252 18680 26280 18711
rect 25096 18652 26280 18680
rect 25096 18640 25102 18652
rect 22646 18612 22652 18624
rect 15804 18584 17632 18612
rect 22607 18584 22652 18612
rect 15804 18572 15810 18584
rect 22646 18572 22652 18584
rect 22704 18572 22710 18624
rect 24302 18572 24308 18624
rect 24360 18612 24366 18624
rect 25409 18615 25467 18621
rect 25409 18612 25421 18615
rect 24360 18584 25421 18612
rect 24360 18572 24366 18584
rect 25409 18581 25421 18584
rect 25455 18581 25467 18615
rect 25409 18575 25467 18581
rect 26050 18572 26056 18624
rect 26108 18612 26114 18624
rect 26712 18612 26740 18711
rect 27706 18708 27712 18720
rect 27764 18708 27770 18760
rect 28350 18748 28356 18760
rect 28263 18720 28356 18748
rect 28350 18708 28356 18720
rect 28408 18748 28414 18760
rect 29454 18748 29460 18760
rect 28408 18720 29460 18748
rect 28408 18708 28414 18720
rect 29454 18708 29460 18720
rect 29512 18708 29518 18760
rect 29638 18708 29644 18760
rect 29696 18748 29702 18760
rect 29733 18751 29791 18757
rect 29733 18748 29745 18751
rect 29696 18720 29745 18748
rect 29696 18708 29702 18720
rect 29733 18717 29745 18720
rect 29779 18717 29791 18751
rect 29733 18711 29791 18717
rect 29822 18708 29828 18760
rect 29880 18748 29886 18760
rect 29917 18751 29975 18757
rect 29917 18748 29929 18751
rect 29880 18720 29929 18748
rect 29880 18708 29886 18720
rect 29917 18717 29929 18720
rect 29963 18717 29975 18751
rect 29917 18711 29975 18717
rect 33413 18751 33471 18757
rect 33413 18717 33425 18751
rect 33459 18748 33471 18751
rect 38286 18748 38292 18760
rect 33459 18720 35894 18748
rect 38247 18720 38292 18748
rect 33459 18717 33471 18720
rect 33413 18711 33471 18717
rect 26108 18584 26740 18612
rect 35866 18612 35894 18720
rect 38286 18708 38292 18720
rect 38344 18708 38350 18760
rect 38105 18615 38163 18621
rect 38105 18612 38117 18615
rect 35866 18584 38117 18612
rect 26108 18572 26114 18584
rect 38105 18581 38117 18584
rect 38151 18581 38163 18615
rect 38105 18575 38163 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 3326 18368 3332 18420
rect 3384 18408 3390 18420
rect 3878 18408 3884 18420
rect 3384 18380 3884 18408
rect 3384 18368 3390 18380
rect 3878 18368 3884 18380
rect 3936 18408 3942 18420
rect 6822 18408 6828 18420
rect 3936 18380 6828 18408
rect 3936 18368 3942 18380
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 12342 18368 12348 18420
rect 12400 18408 12406 18420
rect 20162 18408 20168 18420
rect 12400 18380 20168 18408
rect 12400 18368 12406 18380
rect 20162 18368 20168 18380
rect 20220 18368 20226 18420
rect 26234 18408 26240 18420
rect 24044 18380 26240 18408
rect 4062 18300 4068 18352
rect 4120 18340 4126 18352
rect 4890 18340 4896 18352
rect 4120 18312 4896 18340
rect 4120 18300 4126 18312
rect 4890 18300 4896 18312
rect 4948 18300 4954 18352
rect 14918 18340 14924 18352
rect 14398 18312 14924 18340
rect 14918 18300 14924 18312
rect 14976 18300 14982 18352
rect 23842 18340 23848 18352
rect 15856 18312 23848 18340
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 1578 18164 1584 18216
rect 1636 18204 1642 18216
rect 2222 18204 2228 18216
rect 1636 18176 2228 18204
rect 1636 18164 1642 18176
rect 2222 18164 2228 18176
rect 2280 18204 2286 18216
rect 2317 18207 2375 18213
rect 2317 18204 2329 18207
rect 2280 18176 2329 18204
rect 2280 18164 2286 18176
rect 2317 18173 2329 18176
rect 2363 18173 2375 18207
rect 2317 18167 2375 18173
rect 2593 18207 2651 18213
rect 2593 18173 2605 18207
rect 2639 18204 2651 18207
rect 3712 18204 3740 18258
rect 3786 18204 3792 18216
rect 2639 18176 3648 18204
rect 3712 18176 3792 18204
rect 2639 18173 2651 18176
rect 2593 18167 2651 18173
rect 3620 18136 3648 18176
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 12894 18204 12900 18216
rect 12855 18176 12900 18204
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13170 18204 13176 18216
rect 13083 18176 13176 18204
rect 13170 18164 13176 18176
rect 13228 18204 13234 18216
rect 15856 18204 15884 18312
rect 23842 18300 23848 18312
rect 23900 18300 23906 18352
rect 16301 18275 16359 18281
rect 16301 18241 16313 18275
rect 16347 18272 16359 18275
rect 16666 18272 16672 18284
rect 16347 18244 16672 18272
rect 16347 18241 16359 18244
rect 16301 18235 16359 18241
rect 16666 18232 16672 18244
rect 16724 18232 16730 18284
rect 17405 18275 17463 18281
rect 17405 18272 17417 18275
rect 16776 18244 17417 18272
rect 13228 18176 15884 18204
rect 13228 18164 13234 18176
rect 9214 18136 9220 18148
rect 3620 18108 9220 18136
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 14645 18139 14703 18145
rect 14645 18105 14657 18139
rect 14691 18105 14703 18139
rect 14645 18099 14703 18105
rect 16117 18139 16175 18145
rect 16117 18105 16129 18139
rect 16163 18136 16175 18139
rect 16776 18136 16804 18244
rect 17405 18241 17417 18244
rect 17451 18241 17463 18275
rect 17405 18235 17463 18241
rect 19150 18232 19156 18284
rect 19208 18272 19214 18284
rect 19797 18275 19855 18281
rect 19797 18272 19809 18275
rect 19208 18244 19809 18272
rect 19208 18232 19214 18244
rect 19797 18241 19809 18244
rect 19843 18241 19855 18275
rect 20898 18272 20904 18284
rect 20859 18244 20904 18272
rect 19797 18235 19855 18241
rect 20898 18232 20904 18244
rect 20956 18232 20962 18284
rect 22465 18275 22523 18281
rect 22465 18241 22477 18275
rect 22511 18272 22523 18275
rect 24044 18272 24072 18380
rect 26234 18368 26240 18380
rect 26292 18408 26298 18420
rect 26602 18408 26608 18420
rect 26292 18380 26608 18408
rect 26292 18368 26298 18380
rect 26602 18368 26608 18380
rect 26660 18368 26666 18420
rect 29638 18408 29644 18420
rect 29599 18380 29644 18408
rect 29638 18368 29644 18380
rect 29696 18368 29702 18420
rect 24302 18340 24308 18352
rect 24263 18312 24308 18340
rect 24302 18300 24308 18312
rect 24360 18300 24366 18352
rect 25498 18340 25504 18352
rect 25459 18312 25504 18340
rect 25498 18300 25504 18312
rect 25556 18300 25562 18352
rect 22511 18244 24072 18272
rect 22511 18241 22523 18244
rect 22465 18235 22523 18241
rect 26786 18232 26792 18284
rect 26844 18272 26850 18284
rect 30282 18272 30288 18284
rect 26844 18244 30288 18272
rect 26844 18232 26850 18244
rect 30282 18232 30288 18244
rect 30340 18272 30346 18284
rect 30469 18275 30527 18281
rect 30469 18272 30481 18275
rect 30340 18244 30481 18272
rect 30340 18232 30346 18244
rect 30469 18241 30481 18244
rect 30515 18241 30527 18275
rect 30469 18235 30527 18241
rect 19981 18207 20039 18213
rect 16163 18108 16804 18136
rect 16868 18176 17448 18204
rect 16163 18105 16175 18108
rect 16117 18099 16175 18105
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18068 1639 18071
rect 2314 18068 2320 18080
rect 1627 18040 2320 18068
rect 1627 18037 1639 18040
rect 1581 18031 1639 18037
rect 2314 18028 2320 18040
rect 2372 18028 2378 18080
rect 4065 18071 4123 18077
rect 4065 18037 4077 18071
rect 4111 18068 4123 18071
rect 7282 18068 7288 18080
rect 4111 18040 7288 18068
rect 4111 18037 4123 18040
rect 4065 18031 4123 18037
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 14550 18028 14556 18080
rect 14608 18068 14614 18080
rect 14660 18068 14688 18099
rect 16868 18068 16896 18176
rect 14608 18040 16896 18068
rect 14608 18028 14614 18040
rect 17218 18028 17224 18080
rect 17276 18068 17282 18080
rect 17420 18068 17448 18176
rect 19981 18173 19993 18207
rect 20027 18204 20039 18207
rect 20993 18207 21051 18213
rect 20993 18204 21005 18207
rect 20027 18176 21005 18204
rect 20027 18173 20039 18176
rect 19981 18167 20039 18173
rect 20993 18173 21005 18176
rect 21039 18173 21051 18207
rect 20993 18167 21051 18173
rect 22554 18164 22560 18216
rect 22612 18204 22618 18216
rect 22649 18207 22707 18213
rect 22649 18204 22661 18207
rect 22612 18176 22661 18204
rect 22612 18164 22618 18176
rect 22649 18173 22661 18176
rect 22695 18173 22707 18207
rect 24210 18204 24216 18216
rect 24171 18176 24216 18204
rect 22649 18167 22707 18173
rect 24210 18164 24216 18176
rect 24268 18164 24274 18216
rect 25406 18204 25412 18216
rect 25367 18176 25412 18204
rect 25406 18164 25412 18176
rect 25464 18164 25470 18216
rect 25685 18207 25743 18213
rect 25685 18173 25697 18207
rect 25731 18173 25743 18207
rect 30926 18204 30932 18216
rect 30887 18176 30932 18204
rect 25685 18167 25743 18173
rect 19334 18096 19340 18148
rect 19392 18136 19398 18148
rect 20070 18136 20076 18148
rect 19392 18108 20076 18136
rect 19392 18096 19398 18108
rect 20070 18096 20076 18108
rect 20128 18096 20134 18148
rect 24765 18139 24823 18145
rect 20180 18108 24716 18136
rect 20180 18068 20208 18108
rect 17276 18040 17321 18068
rect 17420 18040 20208 18068
rect 20441 18071 20499 18077
rect 17276 18028 17282 18040
rect 20441 18037 20453 18071
rect 20487 18068 20499 18071
rect 20622 18068 20628 18080
rect 20487 18040 20628 18068
rect 20487 18037 20499 18040
rect 20441 18031 20499 18037
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 22462 18028 22468 18080
rect 22520 18068 22526 18080
rect 22833 18071 22891 18077
rect 22833 18068 22845 18071
rect 22520 18040 22845 18068
rect 22520 18028 22526 18040
rect 22833 18037 22845 18040
rect 22879 18037 22891 18071
rect 24688 18068 24716 18108
rect 24765 18105 24777 18139
rect 24811 18136 24823 18139
rect 25700 18136 25728 18167
rect 30926 18164 30932 18176
rect 30984 18164 30990 18216
rect 31018 18136 31024 18148
rect 24811 18108 31024 18136
rect 24811 18105 24823 18108
rect 24765 18099 24823 18105
rect 31018 18096 31024 18108
rect 31076 18096 31082 18148
rect 25038 18068 25044 18080
rect 24688 18040 25044 18068
rect 22833 18031 22891 18037
rect 25038 18028 25044 18040
rect 25096 18028 25102 18080
rect 29914 18028 29920 18080
rect 29972 18068 29978 18080
rect 30285 18071 30343 18077
rect 30285 18068 30297 18071
rect 29972 18040 30297 18068
rect 29972 18028 29978 18040
rect 30285 18037 30297 18040
rect 30331 18037 30343 18071
rect 30285 18031 30343 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 4604 17867 4662 17873
rect 4604 17833 4616 17867
rect 4650 17864 4662 17867
rect 5074 17864 5080 17876
rect 4650 17836 5080 17864
rect 4650 17833 4662 17836
rect 4604 17827 4662 17833
rect 5074 17824 5080 17836
rect 5132 17864 5138 17876
rect 10778 17864 10784 17876
rect 5132 17836 10784 17864
rect 5132 17824 5138 17836
rect 10778 17824 10784 17836
rect 10836 17824 10842 17876
rect 14918 17864 14924 17876
rect 14879 17836 14924 17864
rect 14918 17824 14924 17836
rect 14976 17824 14982 17876
rect 17681 17867 17739 17873
rect 17681 17833 17693 17867
rect 17727 17864 17739 17867
rect 18230 17864 18236 17876
rect 17727 17836 18236 17864
rect 17727 17833 17739 17836
rect 17681 17827 17739 17833
rect 18230 17824 18236 17836
rect 18288 17864 18294 17876
rect 18874 17864 18880 17876
rect 18288 17836 18880 17864
rect 18288 17824 18294 17836
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 22097 17867 22155 17873
rect 22097 17833 22109 17867
rect 22143 17864 22155 17867
rect 22554 17864 22560 17876
rect 22143 17836 22560 17864
rect 22143 17833 22155 17836
rect 22097 17827 22155 17833
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 25133 17867 25191 17873
rect 25133 17833 25145 17867
rect 25179 17864 25191 17867
rect 25498 17864 25504 17876
rect 25179 17836 25504 17864
rect 25179 17833 25191 17836
rect 25133 17827 25191 17833
rect 25498 17824 25504 17836
rect 25556 17824 25562 17876
rect 29733 17867 29791 17873
rect 29733 17833 29745 17867
rect 29779 17864 29791 17867
rect 29822 17864 29828 17876
rect 29779 17836 29828 17864
rect 29779 17833 29791 17836
rect 29733 17827 29791 17833
rect 29822 17824 29828 17836
rect 29880 17824 29886 17876
rect 12434 17756 12440 17808
rect 12492 17796 12498 17808
rect 12492 17768 18276 17796
rect 12492 17756 12498 17768
rect 4338 17728 4344 17740
rect 4299 17700 4344 17728
rect 4338 17688 4344 17700
rect 4396 17728 4402 17740
rect 4614 17728 4620 17740
rect 4396 17700 4620 17728
rect 4396 17688 4402 17700
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 5074 17688 5080 17740
rect 5132 17728 5138 17740
rect 5132 17700 10548 17728
rect 5132 17688 5138 17700
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 8996 17632 9137 17660
rect 8996 17620 9002 17632
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 10520 17646 10548 17700
rect 14918 17688 14924 17740
rect 14976 17728 14982 17740
rect 17218 17728 17224 17740
rect 14976 17700 15792 17728
rect 17179 17700 17224 17728
rect 14976 17688 14982 17700
rect 14829 17663 14887 17669
rect 9125 17623 9183 17629
rect 14829 17629 14841 17663
rect 14875 17660 14887 17663
rect 15470 17660 15476 17672
rect 14875 17632 15476 17660
rect 14875 17629 14887 17632
rect 14829 17623 14887 17629
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 15764 17669 15792 17700
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 18248 17737 18276 17768
rect 20806 17756 20812 17808
rect 20864 17796 20870 17808
rect 20901 17799 20959 17805
rect 20901 17796 20913 17799
rect 20864 17768 20913 17796
rect 20864 17756 20870 17768
rect 20901 17765 20913 17768
rect 20947 17765 20959 17799
rect 26326 17796 26332 17808
rect 20901 17759 20959 17765
rect 22848 17768 26332 17796
rect 18233 17731 18291 17737
rect 18233 17697 18245 17731
rect 18279 17697 18291 17731
rect 18233 17691 18291 17697
rect 20349 17731 20407 17737
rect 20349 17697 20361 17731
rect 20395 17728 20407 17731
rect 22462 17728 22468 17740
rect 20395 17700 22468 17728
rect 20395 17697 20407 17700
rect 20349 17691 20407 17697
rect 22462 17688 22468 17700
rect 22520 17688 22526 17740
rect 22646 17728 22652 17740
rect 22607 17700 22652 17728
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 22848 17737 22876 17768
rect 26326 17756 26332 17768
rect 26384 17756 26390 17808
rect 26418 17756 26424 17808
rect 26476 17796 26482 17808
rect 26789 17799 26847 17805
rect 26789 17796 26801 17799
rect 26476 17768 26801 17796
rect 26476 17756 26482 17768
rect 26789 17765 26801 17768
rect 26835 17796 26847 17799
rect 28077 17799 28135 17805
rect 28077 17796 28089 17799
rect 26835 17768 28089 17796
rect 26835 17765 26847 17768
rect 26789 17759 26847 17765
rect 28077 17765 28089 17768
rect 28123 17765 28135 17799
rect 28077 17759 28135 17765
rect 22833 17731 22891 17737
rect 22833 17697 22845 17731
rect 22879 17697 22891 17731
rect 22833 17691 22891 17697
rect 26602 17688 26608 17740
rect 26660 17728 26666 17740
rect 27709 17731 27767 17737
rect 27709 17728 27721 17731
rect 26660 17700 27721 17728
rect 26660 17688 26666 17700
rect 27709 17697 27721 17700
rect 27755 17697 27767 17731
rect 27709 17691 27767 17697
rect 30377 17731 30435 17737
rect 30377 17697 30389 17731
rect 30423 17728 30435 17731
rect 30926 17728 30932 17740
rect 30423 17700 30932 17728
rect 30423 17697 30435 17700
rect 30377 17691 30435 17697
rect 30926 17688 30932 17700
rect 30984 17688 30990 17740
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17660 15807 17663
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 15795 17632 16405 17660
rect 15795 17629 15807 17632
rect 15749 17623 15807 17629
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 17037 17663 17095 17669
rect 17037 17629 17049 17663
rect 17083 17660 17095 17663
rect 17862 17660 17868 17672
rect 17083 17632 17868 17660
rect 17083 17629 17095 17632
rect 17037 17623 17095 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 22002 17660 22008 17672
rect 21963 17632 22008 17660
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 25038 17660 25044 17672
rect 24999 17632 25044 17660
rect 25038 17620 25044 17632
rect 25096 17620 25102 17672
rect 26145 17663 26203 17669
rect 26145 17629 26157 17663
rect 26191 17629 26203 17663
rect 26326 17660 26332 17672
rect 26287 17632 26332 17660
rect 26145 17623 26203 17629
rect 6362 17592 6368 17604
rect 5842 17564 6224 17592
rect 6323 17564 6368 17592
rect 6196 17524 6224 17564
rect 6362 17552 6368 17564
rect 6420 17552 6426 17604
rect 9398 17592 9404 17604
rect 9359 17564 9404 17592
rect 9398 17552 9404 17564
rect 9456 17552 9462 17604
rect 16485 17595 16543 17601
rect 16485 17592 16497 17595
rect 10704 17564 16497 17592
rect 10704 17524 10732 17564
rect 16485 17561 16497 17564
rect 16531 17561 16543 17595
rect 16485 17555 16543 17561
rect 18322 17552 18328 17604
rect 18380 17592 18386 17604
rect 18877 17595 18935 17601
rect 18380 17564 18425 17592
rect 18380 17552 18386 17564
rect 18877 17561 18889 17595
rect 18923 17592 18935 17595
rect 19334 17592 19340 17604
rect 18923 17564 19340 17592
rect 18923 17561 18935 17564
rect 18877 17555 18935 17561
rect 19334 17552 19340 17564
rect 19392 17552 19398 17604
rect 20438 17592 20444 17604
rect 20399 17564 20444 17592
rect 20438 17552 20444 17564
rect 20496 17552 20502 17604
rect 26160 17592 26188 17623
rect 26326 17620 26332 17632
rect 26384 17620 26390 17672
rect 27890 17660 27896 17672
rect 27851 17632 27896 17660
rect 27890 17620 27896 17632
rect 27948 17620 27954 17672
rect 29181 17663 29239 17669
rect 29181 17629 29193 17663
rect 29227 17629 29239 17663
rect 29914 17660 29920 17672
rect 29875 17632 29920 17660
rect 29181 17623 29239 17629
rect 26234 17592 26240 17604
rect 26160 17564 26240 17592
rect 26234 17552 26240 17564
rect 26292 17552 26298 17604
rect 27338 17552 27344 17604
rect 27396 17592 27402 17604
rect 29196 17592 29224 17623
rect 29914 17620 29920 17632
rect 29972 17620 29978 17672
rect 30558 17660 30564 17672
rect 30519 17632 30564 17660
rect 30558 17620 30564 17632
rect 30616 17620 30622 17672
rect 30374 17592 30380 17604
rect 27396 17564 30380 17592
rect 27396 17552 27402 17564
rect 30374 17552 30380 17564
rect 30432 17552 30438 17604
rect 6196 17496 10732 17524
rect 10873 17527 10931 17533
rect 10873 17493 10885 17527
rect 10919 17524 10931 17527
rect 13630 17524 13636 17536
rect 10919 17496 13636 17524
rect 10919 17493 10931 17496
rect 10873 17487 10931 17493
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 15838 17524 15844 17536
rect 15799 17496 15844 17524
rect 15838 17484 15844 17496
rect 15896 17484 15902 17536
rect 17954 17484 17960 17536
rect 18012 17524 18018 17536
rect 20530 17524 20536 17536
rect 18012 17496 20536 17524
rect 18012 17484 18018 17496
rect 20530 17484 20536 17496
rect 20588 17484 20594 17536
rect 23293 17527 23351 17533
rect 23293 17493 23305 17527
rect 23339 17524 23351 17527
rect 24210 17524 24216 17536
rect 23339 17496 24216 17524
rect 23339 17493 23351 17496
rect 23293 17487 23351 17493
rect 24210 17484 24216 17496
rect 24268 17484 24274 17536
rect 28994 17524 29000 17536
rect 28955 17496 29000 17524
rect 28994 17484 29000 17496
rect 29052 17484 29058 17536
rect 31018 17524 31024 17536
rect 30979 17496 31024 17524
rect 31018 17484 31024 17496
rect 31076 17484 31082 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 9125 17323 9183 17329
rect 9125 17289 9137 17323
rect 9171 17320 9183 17323
rect 9214 17320 9220 17332
rect 9171 17292 9220 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 18233 17323 18291 17329
rect 9364 17292 16160 17320
rect 9364 17280 9370 17292
rect 7653 17255 7711 17261
rect 7653 17221 7665 17255
rect 7699 17252 7711 17255
rect 7926 17252 7932 17264
rect 7699 17224 7932 17252
rect 7699 17221 7711 17224
rect 7653 17215 7711 17221
rect 7926 17212 7932 17224
rect 7984 17212 7990 17264
rect 8662 17212 8668 17264
rect 8720 17212 8726 17264
rect 13538 17252 13544 17264
rect 13499 17224 13544 17252
rect 13538 17212 13544 17224
rect 13596 17212 13602 17264
rect 15838 17252 15844 17264
rect 14766 17224 15844 17252
rect 15838 17212 15844 17224
rect 15896 17212 15902 17264
rect 16132 17252 16160 17292
rect 18233 17289 18245 17323
rect 18279 17320 18291 17323
rect 18322 17320 18328 17332
rect 18279 17292 18328 17320
rect 18279 17289 18291 17292
rect 18233 17283 18291 17289
rect 18322 17280 18328 17292
rect 18380 17280 18386 17332
rect 20438 17280 20444 17332
rect 20496 17320 20502 17332
rect 21177 17323 21235 17329
rect 21177 17320 21189 17323
rect 20496 17292 21189 17320
rect 20496 17280 20502 17292
rect 21177 17289 21189 17292
rect 21223 17289 21235 17323
rect 27249 17323 27307 17329
rect 21177 17283 21235 17289
rect 23124 17292 27200 17320
rect 17954 17252 17960 17264
rect 16132 17224 17960 17252
rect 16132 17193 16160 17224
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 18966 17252 18972 17264
rect 18927 17224 18972 17252
rect 18966 17212 18972 17224
rect 19024 17212 19030 17264
rect 23124 17252 23152 17292
rect 25958 17252 25964 17264
rect 19996 17224 23152 17252
rect 25919 17224 25964 17252
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17184 16267 17187
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16255 17156 17049 17184
rect 16255 17153 16267 17156
rect 16209 17147 16267 17153
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 18141 17187 18199 17193
rect 18141 17153 18153 17187
rect 18187 17184 18199 17187
rect 18414 17184 18420 17196
rect 18187 17156 18420 17184
rect 18187 17153 18199 17156
rect 18141 17147 18199 17153
rect 18414 17144 18420 17156
rect 18472 17144 18478 17196
rect 19996 17193 20024 17224
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 26053 17255 26111 17261
rect 26053 17221 26065 17255
rect 26099 17252 26111 17255
rect 26602 17252 26608 17264
rect 26099 17224 26608 17252
rect 26099 17221 26111 17224
rect 26053 17215 26111 17221
rect 26602 17212 26608 17224
rect 26660 17212 26666 17264
rect 27172 17252 27200 17292
rect 27249 17289 27261 17323
rect 27295 17320 27307 17323
rect 27890 17320 27896 17332
rect 27295 17292 27896 17320
rect 27295 17289 27307 17292
rect 27249 17283 27307 17289
rect 27890 17280 27896 17292
rect 27948 17280 27954 17332
rect 29825 17323 29883 17329
rect 29825 17289 29837 17323
rect 29871 17320 29883 17323
rect 30558 17320 30564 17332
rect 29871 17292 30564 17320
rect 29871 17289 29883 17292
rect 29825 17283 29883 17289
rect 30558 17280 30564 17292
rect 30616 17280 30622 17332
rect 31018 17280 31024 17332
rect 31076 17320 31082 17332
rect 32953 17323 33011 17329
rect 32953 17320 32965 17323
rect 31076 17292 32965 17320
rect 31076 17280 31082 17292
rect 32953 17289 32965 17292
rect 32999 17289 33011 17323
rect 32953 17283 33011 17289
rect 31754 17252 31760 17264
rect 27172 17224 31760 17252
rect 31754 17212 31760 17224
rect 31812 17212 31818 17264
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17153 20039 17187
rect 20622 17184 20628 17196
rect 19981 17147 20039 17153
rect 20088 17156 20628 17184
rect 4338 17076 4344 17128
rect 4396 17116 4402 17128
rect 5166 17116 5172 17128
rect 4396 17088 5172 17116
rect 4396 17076 4402 17088
rect 5166 17076 5172 17088
rect 5224 17116 5230 17128
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 5224 17088 7389 17116
rect 5224 17076 5230 17088
rect 7377 17085 7389 17088
rect 7423 17116 7435 17119
rect 8938 17116 8944 17128
rect 7423 17088 8944 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 8938 17076 8944 17088
rect 8996 17076 9002 17128
rect 12894 17076 12900 17128
rect 12952 17116 12958 17128
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 12952 17088 13277 17116
rect 12952 17076 12958 17088
rect 13265 17085 13277 17088
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 13630 17076 13636 17128
rect 13688 17116 13694 17128
rect 16853 17119 16911 17125
rect 13688 17088 14583 17116
rect 13688 17076 13694 17088
rect 14555 17048 14583 17088
rect 16853 17085 16865 17119
rect 16899 17116 16911 17119
rect 17586 17116 17592 17128
rect 16899 17088 17592 17116
rect 16899 17085 16911 17088
rect 16853 17079 16911 17085
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 18877 17119 18935 17125
rect 18877 17085 18889 17119
rect 18923 17116 18935 17119
rect 20088 17116 20116 17156
rect 20622 17144 20628 17156
rect 20680 17144 20686 17196
rect 21082 17184 21088 17196
rect 21043 17156 21088 17184
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 22557 17187 22615 17193
rect 22557 17153 22569 17187
rect 22603 17184 22615 17187
rect 27157 17187 27215 17193
rect 22603 17156 24440 17184
rect 22603 17153 22615 17156
rect 22557 17147 22615 17153
rect 18923 17088 20116 17116
rect 20165 17119 20223 17125
rect 18923 17085 18935 17088
rect 18877 17079 18935 17085
rect 20165 17085 20177 17119
rect 20211 17116 20223 17119
rect 20990 17116 20996 17128
rect 20211 17088 20996 17116
rect 20211 17085 20223 17088
rect 20165 17079 20223 17085
rect 20990 17076 20996 17088
rect 21048 17076 21054 17128
rect 22741 17119 22799 17125
rect 22741 17085 22753 17119
rect 22787 17085 22799 17119
rect 24412 17116 24440 17156
rect 27157 17153 27169 17187
rect 27203 17184 27215 17187
rect 27338 17184 27344 17196
rect 27203 17156 27344 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 27338 17144 27344 17156
rect 27396 17144 27402 17196
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 30009 17187 30067 17193
rect 30009 17184 30021 17187
rect 29052 17156 30021 17184
rect 29052 17144 29058 17156
rect 30009 17153 30021 17156
rect 30055 17153 30067 17187
rect 30009 17147 30067 17153
rect 30374 17144 30380 17196
rect 30432 17184 30438 17196
rect 30469 17187 30527 17193
rect 30469 17184 30481 17187
rect 30432 17156 30481 17184
rect 30432 17144 30438 17156
rect 30469 17153 30481 17156
rect 30515 17153 30527 17187
rect 30469 17147 30527 17153
rect 30561 17187 30619 17193
rect 30561 17153 30573 17187
rect 30607 17184 30619 17187
rect 32493 17187 32551 17193
rect 32493 17184 32505 17187
rect 30607 17156 32505 17184
rect 30607 17153 30619 17156
rect 30561 17147 30619 17153
rect 32493 17153 32505 17156
rect 32539 17153 32551 17187
rect 38286 17184 38292 17196
rect 38247 17156 38292 17184
rect 32493 17147 32551 17153
rect 38286 17144 38292 17156
rect 38344 17144 38350 17196
rect 26234 17116 26240 17128
rect 24412 17088 26240 17116
rect 22741 17079 22799 17085
rect 14555 17020 17632 17048
rect 14642 16940 14648 16992
rect 14700 16980 14706 16992
rect 15013 16983 15071 16989
rect 15013 16980 15025 16983
rect 14700 16952 15025 16980
rect 14700 16940 14706 16952
rect 15013 16949 15025 16952
rect 15059 16949 15071 16983
rect 17494 16980 17500 16992
rect 17455 16952 17500 16980
rect 15013 16943 15071 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 17604 16980 17632 17020
rect 18506 17008 18512 17060
rect 18564 17048 18570 17060
rect 19429 17051 19487 17057
rect 19429 17048 19441 17051
rect 18564 17020 19441 17048
rect 18564 17008 18570 17020
rect 19429 17017 19441 17020
rect 19475 17017 19487 17051
rect 22756 17048 22784 17079
rect 26234 17076 26240 17088
rect 26292 17076 26298 17128
rect 32309 17119 32367 17125
rect 32309 17085 32321 17119
rect 32355 17116 32367 17119
rect 32398 17116 32404 17128
rect 32355 17088 32404 17116
rect 32355 17085 32367 17088
rect 32309 17079 32367 17085
rect 32398 17076 32404 17088
rect 32456 17076 32462 17128
rect 24762 17048 24768 17060
rect 22756 17020 24768 17048
rect 19429 17011 19487 17017
rect 24762 17008 24768 17020
rect 24820 17008 24826 17060
rect 26510 17048 26516 17060
rect 26471 17020 26516 17048
rect 26510 17008 26516 17020
rect 26568 17008 26574 17060
rect 22278 16980 22284 16992
rect 17604 16952 22284 16980
rect 22278 16940 22284 16952
rect 22336 16940 22342 16992
rect 22462 16940 22468 16992
rect 22520 16980 22526 16992
rect 22925 16983 22983 16989
rect 22925 16980 22937 16983
rect 22520 16952 22937 16980
rect 22520 16940 22526 16952
rect 22925 16949 22937 16952
rect 22971 16949 22983 16983
rect 22925 16943 22983 16949
rect 35894 16940 35900 16992
rect 35952 16980 35958 16992
rect 38105 16983 38163 16989
rect 38105 16980 38117 16983
rect 35952 16952 38117 16980
rect 35952 16940 35958 16952
rect 38105 16949 38117 16952
rect 38151 16949 38163 16983
rect 38105 16943 38163 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 6168 16779 6226 16785
rect 6168 16745 6180 16779
rect 6214 16776 6226 16779
rect 8386 16776 8392 16788
rect 6214 16748 8392 16776
rect 6214 16745 6226 16748
rect 6168 16739 6226 16745
rect 8386 16736 8392 16748
rect 8444 16776 8450 16788
rect 8754 16776 8760 16788
rect 8444 16748 8760 16776
rect 8444 16736 8450 16748
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 18417 16779 18475 16785
rect 12406 16748 18368 16776
rect 5166 16600 5172 16652
rect 5224 16640 5230 16652
rect 5905 16643 5963 16649
rect 5905 16640 5917 16643
rect 5224 16612 5917 16640
rect 5224 16600 5230 16612
rect 5905 16609 5917 16612
rect 5951 16609 5963 16643
rect 5905 16603 5963 16609
rect 10597 16643 10655 16649
rect 10597 16609 10609 16643
rect 10643 16640 10655 16643
rect 11146 16640 11152 16652
rect 10643 16612 11152 16640
rect 10643 16609 10655 16612
rect 10597 16603 10655 16609
rect 11146 16600 11152 16612
rect 11204 16640 11210 16652
rect 12406 16640 12434 16748
rect 16482 16668 16488 16720
rect 16540 16708 16546 16720
rect 16577 16711 16635 16717
rect 16577 16708 16589 16711
rect 16540 16680 16589 16708
rect 16540 16668 16546 16680
rect 16577 16677 16589 16680
rect 16623 16708 16635 16711
rect 16758 16708 16764 16720
rect 16623 16680 16764 16708
rect 16623 16677 16635 16680
rect 16577 16671 16635 16677
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 18340 16708 18368 16748
rect 18417 16745 18429 16779
rect 18463 16776 18475 16779
rect 18966 16776 18972 16788
rect 18463 16748 18972 16776
rect 18463 16745 18475 16748
rect 18417 16739 18475 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 20990 16776 20996 16788
rect 20951 16748 20996 16776
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 23198 16776 23204 16788
rect 22336 16748 23204 16776
rect 22336 16736 22342 16748
rect 23198 16736 23204 16748
rect 23256 16736 23262 16788
rect 32398 16776 32404 16788
rect 32359 16748 32404 16776
rect 32398 16736 32404 16748
rect 32456 16736 32462 16788
rect 21082 16708 21088 16720
rect 18340 16680 21088 16708
rect 21082 16668 21088 16680
rect 21140 16668 21146 16720
rect 15470 16640 15476 16652
rect 11204 16612 12434 16640
rect 15304 16612 15476 16640
rect 11204 16600 11210 16612
rect 1762 16572 1768 16584
rect 1723 16544 1768 16572
rect 1762 16532 1768 16544
rect 1820 16532 1826 16584
rect 8938 16532 8944 16584
rect 8996 16572 9002 16584
rect 10318 16572 10324 16584
rect 8996 16544 10324 16572
rect 8996 16532 9002 16544
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 12805 16575 12863 16581
rect 12805 16541 12817 16575
rect 12851 16572 12863 16575
rect 14826 16572 14832 16584
rect 12851 16544 14832 16572
rect 12851 16541 12863 16544
rect 12805 16535 12863 16541
rect 14826 16532 14832 16544
rect 14884 16532 14890 16584
rect 15304 16581 15332 16612
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 16025 16643 16083 16649
rect 16025 16609 16037 16643
rect 16071 16640 16083 16643
rect 17494 16640 17500 16652
rect 16071 16612 17500 16640
rect 16071 16609 16083 16612
rect 16025 16603 16083 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 27890 16640 27896 16652
rect 26528 16612 27896 16640
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 18104 16544 18337 16572
rect 18104 16532 18110 16544
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 20990 16532 20996 16584
rect 21048 16572 21054 16584
rect 21177 16575 21235 16581
rect 21177 16572 21189 16575
rect 21048 16544 21189 16572
rect 21048 16532 21054 16544
rect 21177 16541 21189 16544
rect 21223 16541 21235 16575
rect 21177 16535 21235 16541
rect 25133 16575 25191 16581
rect 25133 16541 25145 16575
rect 25179 16572 25191 16575
rect 25498 16572 25504 16584
rect 25179 16544 25504 16572
rect 25179 16541 25191 16544
rect 25133 16535 25191 16541
rect 25498 16532 25504 16544
rect 25556 16532 25562 16584
rect 25866 16532 25872 16584
rect 25924 16532 25930 16584
rect 26528 16581 26556 16612
rect 27890 16600 27896 16612
rect 27948 16600 27954 16652
rect 30469 16643 30527 16649
rect 30469 16609 30481 16643
rect 30515 16640 30527 16643
rect 31018 16640 31024 16652
rect 30515 16612 31024 16640
rect 30515 16609 30527 16612
rect 30469 16603 30527 16609
rect 31018 16600 31024 16612
rect 31076 16600 31082 16652
rect 37090 16640 37096 16652
rect 33520 16612 37096 16640
rect 26053 16575 26111 16581
rect 26053 16541 26065 16575
rect 26099 16572 26111 16575
rect 26513 16575 26571 16581
rect 26099 16544 26234 16572
rect 26099 16541 26111 16544
rect 26053 16535 26111 16541
rect 12897 16507 12955 16513
rect 12897 16504 12909 16507
rect 6288 16476 6670 16504
rect 11822 16476 12909 16504
rect 1486 16396 1492 16448
rect 1544 16436 1550 16448
rect 1581 16439 1639 16445
rect 1581 16436 1593 16439
rect 1544 16408 1593 16436
rect 1544 16396 1550 16408
rect 1581 16405 1593 16408
rect 1627 16405 1639 16439
rect 1581 16399 1639 16405
rect 5442 16396 5448 16448
rect 5500 16436 5506 16448
rect 6288 16436 6316 16476
rect 12897 16473 12909 16476
rect 12943 16473 12955 16507
rect 12897 16467 12955 16473
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 16117 16507 16175 16513
rect 13320 16476 15516 16504
rect 13320 16464 13326 16476
rect 5500 16408 6316 16436
rect 5500 16396 5506 16408
rect 7558 16396 7564 16448
rect 7616 16436 7622 16448
rect 7653 16439 7711 16445
rect 7653 16436 7665 16439
rect 7616 16408 7665 16436
rect 7616 16396 7622 16408
rect 7653 16405 7665 16408
rect 7699 16405 7711 16439
rect 7653 16399 7711 16405
rect 12069 16439 12127 16445
rect 12069 16405 12081 16439
rect 12115 16436 12127 16439
rect 13280 16436 13308 16464
rect 15378 16436 15384 16448
rect 12115 16408 13308 16436
rect 15339 16408 15384 16436
rect 12115 16405 12127 16408
rect 12069 16399 12127 16405
rect 15378 16396 15384 16408
rect 15436 16396 15442 16448
rect 15488 16436 15516 16476
rect 16117 16473 16129 16507
rect 16163 16504 16175 16507
rect 16390 16504 16396 16516
rect 16163 16476 16396 16504
rect 16163 16473 16175 16476
rect 16117 16467 16175 16473
rect 16390 16464 16396 16476
rect 16448 16464 16454 16516
rect 23842 16464 23848 16516
rect 23900 16504 23906 16516
rect 25884 16504 25912 16532
rect 23900 16476 25912 16504
rect 26206 16504 26234 16544
rect 26513 16541 26525 16575
rect 26559 16574 26571 16575
rect 26559 16546 26593 16574
rect 27338 16572 27344 16584
rect 26559 16541 26571 16546
rect 27299 16544 27344 16572
rect 26513 16535 26571 16541
rect 27338 16532 27344 16544
rect 27396 16532 27402 16584
rect 30650 16572 30656 16584
rect 30611 16544 30656 16572
rect 30650 16532 30656 16544
rect 30708 16532 30714 16584
rect 33520 16581 33548 16612
rect 37090 16600 37096 16612
rect 37148 16600 37154 16652
rect 32401 16575 32459 16581
rect 32401 16541 32413 16575
rect 32447 16541 32459 16575
rect 32401 16535 32459 16541
rect 33505 16575 33563 16581
rect 33505 16541 33517 16575
rect 33551 16574 33563 16575
rect 33551 16546 33585 16574
rect 33551 16541 33563 16546
rect 33505 16535 33563 16541
rect 32416 16504 32444 16535
rect 26206 16476 27200 16504
rect 32416 16476 35894 16504
rect 23900 16464 23906 16476
rect 19978 16436 19984 16448
rect 15488 16408 19984 16436
rect 19978 16396 19984 16408
rect 20036 16396 20042 16448
rect 24762 16396 24768 16448
rect 24820 16436 24826 16448
rect 24949 16439 25007 16445
rect 24949 16436 24961 16439
rect 24820 16408 24961 16436
rect 24820 16396 24826 16408
rect 24949 16405 24961 16408
rect 24995 16405 25007 16439
rect 24949 16399 25007 16405
rect 25869 16439 25927 16445
rect 25869 16405 25881 16439
rect 25915 16436 25927 16439
rect 26326 16436 26332 16448
rect 25915 16408 26332 16436
rect 25915 16405 25927 16408
rect 25869 16399 25927 16405
rect 26326 16396 26332 16408
rect 26384 16396 26390 16448
rect 26602 16436 26608 16448
rect 26563 16408 26608 16436
rect 26602 16396 26608 16408
rect 26660 16396 26666 16448
rect 27172 16445 27200 16476
rect 35866 16448 35894 16476
rect 27157 16439 27215 16445
rect 27157 16405 27169 16439
rect 27203 16405 27215 16439
rect 31110 16436 31116 16448
rect 31071 16408 31116 16436
rect 27157 16399 27215 16405
rect 31110 16396 31116 16408
rect 31168 16396 31174 16448
rect 33594 16436 33600 16448
rect 33555 16408 33600 16436
rect 33594 16396 33600 16408
rect 33652 16396 33658 16448
rect 35866 16408 35900 16448
rect 35894 16396 35900 16408
rect 35952 16396 35958 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 3970 16232 3976 16244
rect 1872 16204 3976 16232
rect 1872 16173 1900 16204
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 15378 16232 15384 16244
rect 8772 16204 15384 16232
rect 1857 16167 1915 16173
rect 1857 16133 1869 16167
rect 1903 16133 1915 16167
rect 8772 16164 8800 16204
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 19981 16235 20039 16241
rect 19981 16201 19993 16235
rect 20027 16201 20039 16235
rect 20990 16232 20996 16244
rect 20951 16204 20996 16232
rect 19981 16195 20039 16201
rect 11330 16164 11336 16176
rect 3082 16136 8800 16164
rect 10442 16136 11336 16164
rect 1857 16127 1915 16133
rect 11330 16124 11336 16136
rect 11388 16124 11394 16176
rect 13173 16167 13231 16173
rect 13173 16133 13185 16167
rect 13219 16164 13231 16167
rect 13262 16164 13268 16176
rect 13219 16136 13268 16164
rect 13219 16133 13231 16136
rect 13173 16127 13231 16133
rect 13262 16124 13268 16136
rect 13320 16124 13326 16176
rect 17218 16124 17224 16176
rect 17276 16164 17282 16176
rect 17497 16167 17555 16173
rect 17497 16164 17509 16167
rect 17276 16136 17509 16164
rect 17276 16124 17282 16136
rect 17497 16133 17509 16136
rect 17543 16133 17555 16167
rect 17497 16127 17555 16133
rect 18693 16167 18751 16173
rect 18693 16133 18705 16167
rect 18739 16164 18751 16167
rect 19996 16164 20024 16195
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 23106 16192 23112 16244
rect 23164 16232 23170 16244
rect 23201 16235 23259 16241
rect 23201 16232 23213 16235
rect 23164 16204 23213 16232
rect 23164 16192 23170 16204
rect 23201 16201 23213 16204
rect 23247 16201 23259 16235
rect 23201 16195 23259 16201
rect 24210 16192 24216 16244
rect 24268 16232 24274 16244
rect 24397 16235 24455 16241
rect 24397 16232 24409 16235
rect 24268 16204 24409 16232
rect 24268 16192 24274 16204
rect 24397 16201 24409 16204
rect 24443 16201 24455 16235
rect 25498 16232 25504 16244
rect 25459 16204 25504 16232
rect 24397 16195 24455 16201
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 18739 16136 20024 16164
rect 18739 16133 18751 16136
rect 18693 16127 18751 16133
rect 1578 16096 1584 16108
rect 1539 16068 1584 16096
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 8938 16096 8944 16108
rect 8899 16068 8944 16096
rect 8938 16056 8944 16068
rect 8996 16056 9002 16108
rect 14274 16056 14280 16108
rect 14332 16056 14338 16108
rect 19242 16056 19248 16108
rect 19300 16096 19306 16108
rect 20162 16096 20168 16108
rect 19300 16068 19345 16096
rect 20123 16068 20168 16096
rect 19300 16056 19306 16068
rect 20162 16056 20168 16068
rect 20220 16056 20226 16108
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21177 16099 21235 16105
rect 21177 16096 21189 16099
rect 20956 16068 21189 16096
rect 20956 16056 20962 16068
rect 21177 16065 21189 16068
rect 21223 16065 21235 16099
rect 21177 16059 21235 16065
rect 24762 16056 24768 16108
rect 24820 16096 24826 16108
rect 25685 16099 25743 16105
rect 25685 16096 25697 16099
rect 24820 16068 25697 16096
rect 24820 16056 24826 16068
rect 25685 16065 25697 16068
rect 25731 16065 25743 16099
rect 25685 16059 25743 16065
rect 3602 16028 3608 16040
rect 3563 16000 3608 16028
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 9214 16028 9220 16040
rect 9175 16000 9220 16028
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 12894 16028 12900 16040
rect 11020 16000 12900 16028
rect 11020 15988 11026 16000
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 14182 15988 14188 16040
rect 14240 16028 14246 16040
rect 14645 16031 14703 16037
rect 14645 16028 14657 16031
rect 14240 16000 14657 16028
rect 14240 15988 14246 16000
rect 14645 15997 14657 16000
rect 14691 16028 14703 16031
rect 15102 16028 15108 16040
rect 14691 16000 15108 16028
rect 14691 15997 14703 16000
rect 14645 15991 14703 15997
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 17402 16028 17408 16040
rect 17363 16000 17408 16028
rect 17402 15988 17408 16000
rect 17460 15988 17466 16040
rect 18601 16031 18659 16037
rect 18601 15997 18613 16031
rect 18647 16028 18659 16031
rect 18690 16028 18696 16040
rect 18647 16000 18696 16028
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 22186 15988 22192 16040
rect 22244 16028 22250 16040
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 22244 16000 22569 16028
rect 22244 15988 22250 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22738 16028 22744 16040
rect 22699 16000 22744 16028
rect 22557 15991 22615 15997
rect 22738 15988 22744 16000
rect 22796 15988 22802 16040
rect 23753 16031 23811 16037
rect 23753 15997 23765 16031
rect 23799 15997 23811 16031
rect 23934 16028 23940 16040
rect 23895 16000 23940 16028
rect 23753 15991 23811 15997
rect 17957 15963 18015 15969
rect 14568 15932 14780 15960
rect 10594 15852 10600 15904
rect 10652 15892 10658 15904
rect 10689 15895 10747 15901
rect 10689 15892 10701 15895
rect 10652 15864 10701 15892
rect 10652 15852 10658 15864
rect 10689 15861 10701 15864
rect 10735 15892 10747 15895
rect 14568 15892 14596 15932
rect 10735 15864 14596 15892
rect 14752 15892 14780 15932
rect 17957 15929 17969 15963
rect 18003 15960 18015 15963
rect 18506 15960 18512 15972
rect 18003 15932 18512 15960
rect 18003 15929 18015 15932
rect 17957 15923 18015 15929
rect 18506 15920 18512 15932
rect 18564 15920 18570 15972
rect 20438 15920 20444 15972
rect 20496 15960 20502 15972
rect 23768 15960 23796 15991
rect 23934 15988 23940 16000
rect 23992 15988 23998 16040
rect 24578 15988 24584 16040
rect 24636 16028 24642 16040
rect 24857 16031 24915 16037
rect 24857 16028 24869 16031
rect 24636 16000 24869 16028
rect 24636 15988 24642 16000
rect 24857 15997 24869 16000
rect 24903 15997 24915 16031
rect 28442 16028 28448 16040
rect 28403 16000 28448 16028
rect 24857 15991 24915 15997
rect 28442 15988 28448 16000
rect 28500 15988 28506 16040
rect 28534 15988 28540 16040
rect 28592 16028 28598 16040
rect 28629 16031 28687 16037
rect 28629 16028 28641 16031
rect 28592 16000 28641 16028
rect 28592 15988 28598 16000
rect 28629 15997 28641 16000
rect 28675 15997 28687 16031
rect 29546 16028 29552 16040
rect 29507 16000 29552 16028
rect 28629 15991 28687 15997
rect 29546 15988 29552 16000
rect 29604 15988 29610 16040
rect 29733 16031 29791 16037
rect 29733 15997 29745 16031
rect 29779 16028 29791 16031
rect 29822 16028 29828 16040
rect 29779 16000 29828 16028
rect 29779 15997 29791 16000
rect 29733 15991 29791 15997
rect 29822 15988 29828 16000
rect 29880 15988 29886 16040
rect 20496 15932 23796 15960
rect 29089 15963 29147 15969
rect 20496 15920 20502 15932
rect 29089 15929 29101 15963
rect 29135 15960 29147 15963
rect 29917 15963 29975 15969
rect 29917 15960 29929 15963
rect 29135 15932 29929 15960
rect 29135 15929 29147 15932
rect 29089 15923 29147 15929
rect 29917 15929 29929 15932
rect 29963 15960 29975 15963
rect 30098 15960 30104 15972
rect 29963 15932 30104 15960
rect 29963 15929 29975 15932
rect 29917 15923 29975 15929
rect 30098 15920 30104 15932
rect 30156 15920 30162 15972
rect 28350 15892 28356 15904
rect 14752 15864 28356 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 3602 15648 3608 15700
rect 3660 15688 3666 15700
rect 13170 15688 13176 15700
rect 3660 15660 13176 15688
rect 3660 15648 3666 15660
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 14274 15648 14280 15700
rect 14332 15688 14338 15700
rect 14369 15691 14427 15697
rect 14369 15688 14381 15691
rect 14332 15660 14381 15688
rect 14332 15648 14338 15660
rect 14369 15657 14381 15660
rect 14415 15657 14427 15691
rect 16390 15688 16396 15700
rect 16351 15660 16396 15688
rect 14369 15651 14427 15657
rect 16390 15648 16396 15660
rect 16448 15648 16454 15700
rect 17218 15688 17224 15700
rect 17179 15660 17224 15688
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 17586 15648 17592 15700
rect 17644 15688 17650 15700
rect 22738 15688 22744 15700
rect 17644 15660 20944 15688
rect 22699 15660 22744 15688
rect 17644 15648 17650 15660
rect 4062 15620 4068 15632
rect 4023 15592 4068 15620
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 15749 15623 15807 15629
rect 15749 15589 15761 15623
rect 15795 15589 15807 15623
rect 15749 15583 15807 15589
rect 17865 15623 17923 15629
rect 17865 15589 17877 15623
rect 17911 15589 17923 15623
rect 17865 15583 17923 15589
rect 18156 15592 20484 15620
rect 10318 15512 10324 15564
rect 10376 15552 10382 15564
rect 10962 15552 10968 15564
rect 10376 15524 10968 15552
rect 10376 15512 10382 15524
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 15764 15552 15792 15583
rect 15764 15524 16620 15552
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15484 4031 15487
rect 4062 15484 4068 15496
rect 4019 15456 4068 15484
rect 4019 15453 4031 15456
rect 3973 15447 4031 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15484 14335 15487
rect 14826 15484 14832 15496
rect 14323 15456 14832 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 15930 15484 15936 15496
rect 15891 15456 15936 15484
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 16592 15493 16620 15524
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15453 16635 15487
rect 16577 15447 16635 15453
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15484 17463 15487
rect 17880 15484 17908 15583
rect 18046 15484 18052 15496
rect 17451 15456 17908 15484
rect 18007 15456 18052 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 11241 15419 11299 15425
rect 11241 15385 11253 15419
rect 11287 15385 11299 15419
rect 12802 15416 12808 15428
rect 12466 15388 12808 15416
rect 11241 15379 11299 15385
rect 11256 15348 11284 15379
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 12986 15376 12992 15428
rect 13044 15416 13050 15428
rect 18156 15416 18184 15592
rect 18690 15552 18696 15564
rect 18651 15524 18696 15552
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 19797 15555 19855 15561
rect 19797 15521 19809 15555
rect 19843 15552 19855 15555
rect 20254 15552 20260 15564
rect 19843 15524 20260 15552
rect 19843 15521 19855 15524
rect 19797 15515 19855 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 20456 15484 20484 15592
rect 20916 15561 20944 15660
rect 22738 15648 22744 15660
rect 22796 15648 22802 15700
rect 23934 15688 23940 15700
rect 23895 15660 23940 15688
rect 23934 15648 23940 15660
rect 23992 15648 23998 15700
rect 25222 15688 25228 15700
rect 25183 15660 25228 15688
rect 25222 15648 25228 15660
rect 25280 15648 25286 15700
rect 27801 15691 27859 15697
rect 27801 15657 27813 15691
rect 27847 15688 27859 15691
rect 28534 15688 28540 15700
rect 27847 15660 28540 15688
rect 27847 15657 27859 15660
rect 27801 15651 27859 15657
rect 28534 15648 28540 15660
rect 28592 15648 28598 15700
rect 29822 15688 29828 15700
rect 29783 15660 29828 15688
rect 29822 15648 29828 15660
rect 29880 15648 29886 15700
rect 30377 15691 30435 15697
rect 30377 15657 30389 15691
rect 30423 15688 30435 15691
rect 30650 15688 30656 15700
rect 30423 15660 30656 15688
rect 30423 15657 30435 15660
rect 30377 15651 30435 15657
rect 30650 15648 30656 15660
rect 30708 15648 30714 15700
rect 21545 15623 21603 15629
rect 21545 15589 21557 15623
rect 21591 15620 21603 15623
rect 25406 15620 25412 15632
rect 21591 15592 25412 15620
rect 21591 15589 21603 15592
rect 21545 15583 21603 15589
rect 25406 15580 25412 15592
rect 25464 15580 25470 15632
rect 27065 15623 27123 15629
rect 27065 15589 27077 15623
rect 27111 15620 27123 15623
rect 31110 15620 31116 15632
rect 27111 15592 31116 15620
rect 27111 15589 27123 15592
rect 27065 15583 27123 15589
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15521 20959 15555
rect 24578 15552 24584 15564
rect 20901 15515 20959 15521
rect 21008 15524 22094 15552
rect 24539 15524 24584 15552
rect 21008 15484 21036 15524
rect 20456 15456 21036 15484
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15484 21143 15487
rect 21358 15484 21364 15496
rect 21131 15456 21364 15484
rect 21131 15453 21143 15456
rect 21085 15447 21143 15453
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 22066 15484 22094 15524
rect 24578 15512 24584 15524
rect 24636 15512 24642 15564
rect 26418 15552 26424 15564
rect 26379 15524 26424 15552
rect 26418 15512 26424 15524
rect 26476 15512 26482 15564
rect 28442 15552 28448 15564
rect 28403 15524 28448 15552
rect 28442 15512 28448 15524
rect 28500 15512 28506 15564
rect 22646 15484 22652 15496
rect 22066 15456 22652 15484
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 23842 15484 23848 15496
rect 23803 15456 23848 15484
rect 23842 15444 23848 15456
rect 23900 15444 23906 15496
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15484 24823 15487
rect 25866 15484 25872 15496
rect 24811 15456 25872 15484
rect 24811 15453 24823 15456
rect 24765 15447 24823 15453
rect 25866 15444 25872 15456
rect 25924 15444 25930 15496
rect 26602 15484 26608 15496
rect 26563 15456 26608 15484
rect 26602 15444 26608 15456
rect 26660 15444 26666 15496
rect 27982 15484 27988 15496
rect 27943 15456 27988 15484
rect 27982 15444 27988 15456
rect 28040 15444 28046 15496
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 28552 15456 29745 15484
rect 28552 15428 28580 15456
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 30558 15484 30564 15496
rect 30519 15456 30564 15484
rect 29733 15447 29791 15453
rect 30558 15444 30564 15456
rect 30616 15444 30622 15496
rect 31036 15493 31064 15592
rect 31110 15580 31116 15592
rect 31168 15580 31174 15632
rect 32309 15623 32367 15629
rect 32309 15589 32321 15623
rect 32355 15620 32367 15623
rect 32355 15592 35894 15620
rect 32355 15589 32367 15592
rect 32309 15583 32367 15589
rect 31021 15487 31079 15493
rect 31021 15453 31033 15487
rect 31067 15453 31079 15487
rect 31021 15447 31079 15453
rect 31665 15487 31723 15493
rect 31665 15453 31677 15487
rect 31711 15484 31723 15487
rect 32398 15484 32404 15496
rect 31711 15456 32404 15484
rect 31711 15453 31723 15456
rect 31665 15447 31723 15453
rect 32398 15444 32404 15456
rect 32456 15444 32462 15496
rect 32493 15487 32551 15493
rect 32493 15453 32505 15487
rect 32539 15453 32551 15487
rect 35866 15484 35894 15592
rect 38013 15487 38071 15493
rect 38013 15484 38025 15487
rect 35866 15456 38025 15484
rect 32493 15447 32551 15453
rect 38013 15453 38025 15456
rect 38059 15453 38071 15487
rect 38013 15447 38071 15453
rect 13044 15388 18184 15416
rect 19889 15419 19947 15425
rect 13044 15376 13050 15388
rect 19889 15385 19901 15419
rect 19935 15385 19947 15419
rect 19889 15379 19947 15385
rect 20441 15419 20499 15425
rect 20441 15385 20453 15419
rect 20487 15416 20499 15419
rect 21266 15416 21272 15428
rect 20487 15388 21272 15416
rect 20487 15385 20499 15388
rect 20441 15379 20499 15385
rect 15378 15348 15384 15360
rect 11256 15320 15384 15348
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 19904 15348 19932 15379
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 22922 15376 22928 15428
rect 22980 15416 22986 15428
rect 28534 15416 28540 15428
rect 22980 15388 28540 15416
rect 22980 15376 22986 15388
rect 28534 15376 28540 15388
rect 28592 15376 28598 15428
rect 31113 15419 31171 15425
rect 31113 15385 31125 15419
rect 31159 15416 31171 15419
rect 32508 15416 32536 15447
rect 31159 15388 32536 15416
rect 31159 15385 31171 15388
rect 31113 15379 31171 15385
rect 20990 15348 20996 15360
rect 19904 15320 20996 15348
rect 20990 15308 20996 15320
rect 21048 15308 21054 15360
rect 28074 15308 28080 15360
rect 28132 15348 28138 15360
rect 31757 15351 31815 15357
rect 31757 15348 31769 15351
rect 28132 15320 31769 15348
rect 28132 15308 28138 15320
rect 31757 15317 31769 15320
rect 31803 15317 31815 15351
rect 38194 15348 38200 15360
rect 38155 15320 38200 15348
rect 31757 15311 31815 15317
rect 38194 15308 38200 15320
rect 38252 15308 38258 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 4433 15147 4491 15153
rect 4433 15113 4445 15147
rect 4479 15144 4491 15147
rect 10502 15144 10508 15156
rect 4479 15116 10508 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 12406 15116 17448 15144
rect 4890 15076 4896 15088
rect 3358 15048 4896 15076
rect 4890 15036 4896 15048
rect 4948 15036 4954 15088
rect 5074 15076 5080 15088
rect 5035 15048 5080 15076
rect 5074 15036 5080 15048
rect 5132 15036 5138 15088
rect 12158 15076 12164 15088
rect 8970 15048 12164 15076
rect 12158 15036 12164 15048
rect 12216 15036 12222 15088
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 1857 15011 1915 15017
rect 1857 15008 1869 15011
rect 1636 14980 1869 15008
rect 1636 14968 1642 14980
rect 1857 14977 1869 14980
rect 1903 14977 1915 15011
rect 3878 15008 3884 15020
rect 3839 14980 3884 15008
rect 1857 14971 1915 14977
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4341 15011 4399 15017
rect 4341 15008 4353 15011
rect 4120 14980 4353 15008
rect 4120 14968 4126 14980
rect 4341 14977 4353 14980
rect 4387 14977 4399 15011
rect 4341 14971 4399 14977
rect 4985 15011 5043 15017
rect 4985 14977 4997 15011
rect 5031 14977 5043 15011
rect 12406 15008 12434 15116
rect 16574 15076 16580 15088
rect 15226 15048 16580 15076
rect 16574 15036 16580 15048
rect 16632 15036 16638 15088
rect 17420 15076 17448 15116
rect 17494 15104 17500 15156
rect 17552 15144 17558 15156
rect 17589 15147 17647 15153
rect 17589 15144 17601 15147
rect 17552 15116 17601 15144
rect 17552 15104 17558 15116
rect 17589 15113 17601 15116
rect 17635 15113 17647 15147
rect 17589 15107 17647 15113
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15144 19947 15147
rect 20162 15144 20168 15156
rect 19935 15116 20168 15144
rect 19935 15113 19947 15116
rect 19889 15107 19947 15113
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20990 15144 20996 15156
rect 20951 15116 20996 15144
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 25222 15104 25228 15156
rect 25280 15144 25286 15156
rect 25409 15147 25467 15153
rect 25409 15144 25421 15147
rect 25280 15116 25421 15144
rect 25280 15104 25286 15116
rect 25409 15113 25421 15116
rect 25455 15113 25467 15147
rect 25866 15144 25872 15156
rect 25827 15116 25872 15144
rect 25409 15107 25467 15113
rect 25866 15104 25872 15116
rect 25924 15104 25930 15156
rect 26602 15104 26608 15156
rect 26660 15144 26666 15156
rect 27249 15147 27307 15153
rect 27249 15144 27261 15147
rect 26660 15116 27261 15144
rect 26660 15104 26666 15116
rect 27249 15113 27261 15116
rect 27295 15113 27307 15147
rect 27249 15107 27307 15113
rect 27982 15104 27988 15156
rect 28040 15144 28046 15156
rect 28353 15147 28411 15153
rect 28353 15144 28365 15147
rect 28040 15116 28365 15144
rect 28040 15104 28046 15116
rect 28353 15113 28365 15116
rect 28399 15113 28411 15147
rect 28353 15107 28411 15113
rect 28997 15147 29055 15153
rect 28997 15113 29009 15147
rect 29043 15144 29055 15147
rect 30558 15144 30564 15156
rect 29043 15116 30564 15144
rect 29043 15113 29055 15116
rect 28997 15107 29055 15113
rect 30558 15104 30564 15116
rect 30616 15104 30622 15156
rect 18046 15076 18052 15088
rect 17420 15048 18052 15076
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 22002 15076 22008 15088
rect 18156 15048 22008 15076
rect 18156 15008 18184 15048
rect 22002 15036 22008 15048
rect 22060 15076 22066 15088
rect 24394 15076 24400 15088
rect 22060 15048 24400 15076
rect 22060 15036 22066 15048
rect 24394 15036 24400 15048
rect 24452 15076 24458 15088
rect 24762 15076 24768 15088
rect 24452 15048 24768 15076
rect 24452 15036 24458 15048
rect 24762 15036 24768 15048
rect 24820 15036 24826 15088
rect 27172 15048 29224 15076
rect 20070 15008 20076 15020
rect 4985 14971 5043 14977
rect 8956 14980 12434 15008
rect 15764 14980 18184 15008
rect 20031 14980 20076 15008
rect 2130 14940 2136 14952
rect 2091 14912 2136 14940
rect 2130 14900 2136 14912
rect 2188 14900 2194 14952
rect 5000 14872 5028 14971
rect 5166 14900 5172 14952
rect 5224 14940 5230 14952
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 5224 14912 7481 14940
rect 5224 14900 5230 14912
rect 7469 14909 7481 14912
rect 7515 14909 7527 14943
rect 7742 14940 7748 14952
rect 7655 14912 7748 14940
rect 7469 14903 7527 14909
rect 7742 14900 7748 14912
rect 7800 14940 7806 14952
rect 8956 14940 8984 14980
rect 9490 14940 9496 14952
rect 7800 14912 8984 14940
rect 9451 14912 9496 14940
rect 7800 14900 7806 14912
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 12952 14912 13737 14940
rect 12952 14900 12958 14912
rect 13725 14909 13737 14912
rect 13771 14909 13783 14943
rect 13998 14940 14004 14952
rect 13959 14912 14004 14940
rect 13725 14903 13783 14909
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 15764 14949 15792 14980
rect 20070 14968 20076 14980
rect 20128 14968 20134 15020
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 15749 14943 15807 14949
rect 15749 14940 15761 14943
rect 15028 14912 15761 14940
rect 12618 14872 12624 14884
rect 5000 14844 7604 14872
rect 7576 14804 7604 14844
rect 8772 14844 12624 14872
rect 8772 14804 8800 14844
rect 12618 14832 12624 14844
rect 12676 14832 12682 14884
rect 7576 14776 8800 14804
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 15028 14804 15056 14912
rect 15749 14909 15761 14912
rect 15795 14909 15807 14943
rect 16942 14940 16948 14952
rect 16903 14912 16948 14940
rect 15749 14903 15807 14909
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 17954 14940 17960 14952
rect 17175 14912 17960 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 17954 14900 17960 14912
rect 18012 14900 18018 14952
rect 20916 14940 20944 14971
rect 21174 14968 21180 15020
rect 21232 15008 21238 15020
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 21232 14980 22201 15008
rect 21232 14968 21238 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 25590 14968 25596 15020
rect 25648 15008 25654 15020
rect 26053 15011 26111 15017
rect 26053 15008 26065 15011
rect 25648 14980 26065 15008
rect 25648 14968 25654 14980
rect 26053 14977 26065 14980
rect 26099 14977 26111 15011
rect 26053 14971 26111 14977
rect 27062 14968 27068 15020
rect 27120 15008 27126 15020
rect 27172 15017 27200 15048
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 27120 14980 27169 15008
rect 27120 14968 27126 14980
rect 27157 14977 27169 14980
rect 27203 14977 27215 15011
rect 28534 15008 28540 15020
rect 28495 14980 28540 15008
rect 27157 14971 27215 14977
rect 28534 14968 28540 14980
rect 28592 14968 28598 15020
rect 29196 15017 29224 15048
rect 29181 15011 29239 15017
rect 29181 14977 29193 15011
rect 29227 14977 29239 15011
rect 29181 14971 29239 14977
rect 24670 14940 24676 14952
rect 20916 14912 24676 14940
rect 15102 14832 15108 14884
rect 15160 14872 15166 14884
rect 20916 14872 20944 14912
rect 24670 14900 24676 14912
rect 24728 14900 24734 14952
rect 24765 14943 24823 14949
rect 24765 14909 24777 14943
rect 24811 14909 24823 14943
rect 24765 14903 24823 14909
rect 24949 14943 25007 14949
rect 24949 14909 24961 14943
rect 24995 14940 25007 14943
rect 26326 14940 26332 14952
rect 24995 14912 26332 14940
rect 24995 14909 25007 14912
rect 24949 14903 25007 14909
rect 15160 14844 20944 14872
rect 15160 14832 15166 14844
rect 21542 14832 21548 14884
rect 21600 14872 21606 14884
rect 24578 14872 24584 14884
rect 21600 14844 24584 14872
rect 21600 14832 21606 14844
rect 24578 14832 24584 14844
rect 24636 14832 24642 14884
rect 24780 14872 24808 14903
rect 26326 14900 26332 14912
rect 26384 14900 26390 14952
rect 27522 14872 27528 14884
rect 24780 14844 27528 14872
rect 27522 14832 27528 14844
rect 27580 14832 27586 14884
rect 9732 14776 15056 14804
rect 22005 14807 22063 14813
rect 9732 14764 9738 14776
rect 22005 14773 22017 14807
rect 22051 14804 22063 14807
rect 22830 14804 22836 14816
rect 22051 14776 22836 14804
rect 22051 14773 22063 14776
rect 22005 14767 22063 14773
rect 22830 14764 22836 14776
rect 22888 14764 22894 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 3329 14603 3387 14609
rect 3329 14569 3341 14603
rect 3375 14600 3387 14603
rect 4706 14600 4712 14612
rect 3375 14572 4712 14600
rect 3375 14569 3387 14572
rect 3329 14563 3387 14569
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 6641 14603 6699 14609
rect 6641 14569 6653 14603
rect 6687 14600 6699 14603
rect 7742 14600 7748 14612
rect 6687 14572 7748 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 11146 14600 11152 14612
rect 11107 14572 11152 14600
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 15473 14603 15531 14609
rect 15473 14600 15485 14603
rect 11388 14572 15485 14600
rect 11388 14560 11394 14572
rect 15473 14569 15485 14572
rect 15519 14569 15531 14603
rect 21358 14600 21364 14612
rect 21319 14572 21364 14600
rect 15473 14563 15531 14569
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 21468 14572 26234 14600
rect 4157 14535 4215 14541
rect 4157 14501 4169 14535
rect 4203 14532 4215 14535
rect 4798 14532 4804 14544
rect 4203 14504 4804 14532
rect 4203 14501 4215 14504
rect 4157 14495 4215 14501
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 6380 14504 9536 14532
rect 2498 14424 2504 14476
rect 2556 14464 2562 14476
rect 4893 14467 4951 14473
rect 4893 14464 4905 14467
rect 2556 14436 4905 14464
rect 2556 14424 2562 14436
rect 4893 14433 4905 14436
rect 4939 14464 4951 14467
rect 5166 14464 5172 14476
rect 4939 14436 5172 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 5166 14424 5172 14436
rect 5224 14424 5230 14476
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14396 3295 14399
rect 3326 14396 3332 14408
rect 3283 14368 3332 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 3326 14356 3332 14368
rect 3384 14396 3390 14408
rect 4062 14396 4068 14408
rect 3384 14368 4068 14396
rect 3384 14356 3390 14368
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 6380 14396 6408 14504
rect 8938 14424 8944 14476
rect 8996 14464 9002 14476
rect 9398 14464 9404 14476
rect 8996 14436 9404 14464
rect 8996 14424 9002 14436
rect 9398 14424 9404 14436
rect 9456 14424 9462 14476
rect 9508 14464 9536 14504
rect 10962 14492 10968 14544
rect 11020 14532 11026 14544
rect 11701 14535 11759 14541
rect 11701 14532 11713 14535
rect 11020 14504 11713 14532
rect 11020 14492 11026 14504
rect 11701 14501 11713 14504
rect 11747 14501 11759 14535
rect 11701 14495 11759 14501
rect 16758 14492 16764 14544
rect 16816 14532 16822 14544
rect 21468 14532 21496 14572
rect 16816 14504 21496 14532
rect 22005 14535 22063 14541
rect 16816 14492 16822 14504
rect 22005 14501 22017 14535
rect 22051 14501 22063 14535
rect 25590 14532 25596 14544
rect 25551 14504 25596 14532
rect 22005 14495 22063 14501
rect 14829 14467 14887 14473
rect 14829 14464 14841 14467
rect 9508 14436 14841 14464
rect 14829 14433 14841 14436
rect 14875 14433 14887 14467
rect 14829 14427 14887 14433
rect 15010 14424 15016 14476
rect 15068 14464 15074 14476
rect 15470 14464 15476 14476
rect 15068 14436 15476 14464
rect 15068 14424 15074 14436
rect 15470 14424 15476 14436
rect 15528 14464 15534 14476
rect 16577 14467 16635 14473
rect 16577 14464 16589 14467
rect 15528 14436 16589 14464
rect 15528 14424 15534 14436
rect 16577 14433 16589 14436
rect 16623 14433 16635 14467
rect 16577 14427 16635 14433
rect 16942 14424 16948 14476
rect 17000 14464 17006 14476
rect 17221 14467 17279 14473
rect 17221 14464 17233 14467
rect 17000 14436 17233 14464
rect 17000 14424 17006 14436
rect 17221 14433 17233 14436
rect 17267 14433 17279 14467
rect 17221 14427 17279 14433
rect 19797 14467 19855 14473
rect 19797 14433 19809 14467
rect 19843 14464 19855 14467
rect 20898 14464 20904 14476
rect 19843 14436 20904 14464
rect 19843 14433 19855 14436
rect 19797 14427 19855 14433
rect 20898 14424 20904 14436
rect 20956 14424 20962 14476
rect 11606 14396 11612 14408
rect 6302 14368 6408 14396
rect 11519 14368 11612 14396
rect 11606 14356 11612 14368
rect 11664 14396 11670 14408
rect 11664 14368 13768 14396
rect 11664 14356 11670 14368
rect 5169 14331 5227 14337
rect 2746 14300 4292 14328
rect 2130 14220 2136 14272
rect 2188 14260 2194 14272
rect 2746 14260 2774 14300
rect 2188 14232 2774 14260
rect 4264 14260 4292 14300
rect 5169 14297 5181 14331
rect 5215 14328 5227 14331
rect 5258 14328 5264 14340
rect 5215 14300 5264 14328
rect 5215 14297 5227 14300
rect 5169 14291 5227 14297
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 9674 14328 9680 14340
rect 9635 14300 9680 14328
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 11422 14328 11428 14340
rect 10902 14300 11428 14328
rect 11422 14288 11428 14300
rect 11480 14288 11486 14340
rect 5534 14260 5540 14272
rect 4264 14232 5540 14260
rect 2188 14220 2194 14232
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 10318 14260 10324 14272
rect 9272 14232 10324 14260
rect 9272 14220 9278 14232
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 13740 14260 13768 14368
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14734 14396 14740 14408
rect 14516 14368 14740 14396
rect 14516 14356 14522 14368
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14365 15439 14399
rect 16298 14396 16304 14408
rect 16259 14368 16304 14396
rect 15381 14359 15439 14365
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 15396 14328 15424 14359
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 18138 14356 18144 14408
rect 18196 14396 18202 14408
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 18196 14368 18245 14396
rect 18196 14356 18202 14368
rect 18233 14365 18245 14368
rect 18279 14365 18291 14399
rect 18233 14359 18291 14365
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 20806 14396 20812 14408
rect 20487 14368 20812 14396
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 21545 14399 21603 14405
rect 21545 14365 21557 14399
rect 21591 14396 21603 14399
rect 22020 14396 22048 14495
rect 25590 14492 25596 14504
rect 25648 14492 25654 14544
rect 26206 14532 26234 14572
rect 26326 14560 26332 14612
rect 26384 14600 26390 14612
rect 28626 14600 28632 14612
rect 26384 14572 26429 14600
rect 28587 14572 28632 14600
rect 26384 14560 26390 14572
rect 28626 14560 28632 14572
rect 28684 14560 28690 14612
rect 26206 14504 27568 14532
rect 23842 14464 23848 14476
rect 22204 14436 23848 14464
rect 22204 14405 22232 14436
rect 23842 14424 23848 14436
rect 23900 14424 23906 14476
rect 21591 14368 22048 14396
rect 22189 14399 22247 14405
rect 21591 14365 21603 14368
rect 21545 14359 21603 14365
rect 22189 14365 22201 14399
rect 22235 14365 22247 14399
rect 22830 14396 22836 14408
rect 22791 14368 22836 14396
rect 22189 14359 22247 14365
rect 22830 14356 22836 14368
rect 22888 14356 22894 14408
rect 24578 14356 24584 14408
rect 24636 14396 24642 14408
rect 27540 14405 27568 14504
rect 27985 14467 28043 14473
rect 27985 14433 27997 14467
rect 28031 14464 28043 14467
rect 29914 14464 29920 14476
rect 28031 14436 29920 14464
rect 28031 14433 28043 14436
rect 27985 14427 28043 14433
rect 29914 14424 29920 14436
rect 29972 14424 29978 14476
rect 25777 14399 25835 14405
rect 25777 14396 25789 14399
rect 24636 14368 25789 14396
rect 24636 14356 24642 14368
rect 25777 14365 25789 14368
rect 25823 14396 25835 14399
rect 26237 14399 26295 14405
rect 26237 14396 26249 14399
rect 25823 14368 26249 14396
rect 25823 14365 25835 14368
rect 25777 14359 25835 14365
rect 26237 14365 26249 14368
rect 26283 14365 26295 14399
rect 26237 14359 26295 14365
rect 27525 14399 27583 14405
rect 27525 14365 27537 14399
rect 27571 14396 27583 14399
rect 27706 14396 27712 14408
rect 27571 14368 27712 14396
rect 27571 14365 27583 14368
rect 27525 14359 27583 14365
rect 27706 14356 27712 14368
rect 27764 14356 27770 14408
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14396 28227 14399
rect 28258 14396 28264 14408
rect 28215 14368 28264 14396
rect 28215 14365 28227 14368
rect 28169 14359 28227 14365
rect 28258 14356 28264 14368
rect 28316 14356 28322 14408
rect 16666 14328 16672 14340
rect 13872 14300 16672 14328
rect 13872 14288 13878 14300
rect 16666 14288 16672 14300
rect 16724 14288 16730 14340
rect 19889 14331 19947 14337
rect 19889 14297 19901 14331
rect 19935 14297 19947 14331
rect 19889 14291 19947 14297
rect 14826 14260 14832 14272
rect 13740 14232 14832 14260
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 18049 14263 18107 14269
rect 18049 14229 18061 14263
rect 18095 14260 18107 14263
rect 18138 14260 18144 14272
rect 18095 14232 18144 14260
rect 18095 14229 18107 14232
rect 18049 14223 18107 14229
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 18693 14263 18751 14269
rect 18693 14229 18705 14263
rect 18739 14260 18751 14263
rect 18874 14260 18880 14272
rect 18739 14232 18880 14260
rect 18739 14229 18751 14232
rect 18693 14223 18751 14229
rect 18874 14220 18880 14232
rect 18932 14220 18938 14272
rect 19904 14260 19932 14291
rect 20530 14288 20536 14340
rect 20588 14328 20594 14340
rect 26326 14328 26332 14340
rect 20588 14300 26332 14328
rect 20588 14288 20594 14300
rect 26326 14288 26332 14300
rect 26384 14328 26390 14340
rect 26786 14328 26792 14340
rect 26384 14300 26792 14328
rect 26384 14288 26390 14300
rect 26786 14288 26792 14300
rect 26844 14288 26850 14340
rect 22649 14263 22707 14269
rect 22649 14260 22661 14263
rect 19904 14232 22661 14260
rect 22649 14229 22661 14232
rect 22695 14229 22707 14263
rect 22649 14223 22707 14229
rect 27341 14263 27399 14269
rect 27341 14229 27353 14263
rect 27387 14260 27399 14263
rect 28442 14260 28448 14272
rect 27387 14232 28448 14260
rect 27387 14229 27399 14232
rect 27341 14223 27399 14229
rect 28442 14220 28448 14232
rect 28500 14220 28506 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 20530 14056 20536 14068
rect 9548 14028 20536 14056
rect 9548 14016 9554 14028
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 22738 14016 22744 14068
rect 22796 14056 22802 14068
rect 22833 14059 22891 14065
rect 22833 14056 22845 14059
rect 22796 14028 22845 14056
rect 22796 14016 22802 14028
rect 22833 14025 22845 14028
rect 22879 14025 22891 14059
rect 24489 14059 24547 14065
rect 22833 14019 22891 14025
rect 23308 14028 24072 14056
rect 4890 13948 4896 14000
rect 4948 13988 4954 14000
rect 4948 13960 9628 13988
rect 4948 13948 4954 13960
rect 1578 13880 1584 13932
rect 1636 13920 1642 13932
rect 2498 13920 2504 13932
rect 1636 13892 2504 13920
rect 1636 13880 1642 13892
rect 2498 13880 2504 13892
rect 2556 13920 2562 13932
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 2556 13892 2605 13920
rect 2556 13880 2562 13892
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 9490 13920 9496 13932
rect 4002 13892 4108 13920
rect 2593 13883 2651 13889
rect 4080 13864 4108 13892
rect 4264 13892 9496 13920
rect 4062 13812 4068 13864
rect 4120 13812 4126 13864
rect 2856 13719 2914 13725
rect 2856 13685 2868 13719
rect 2902 13716 2914 13719
rect 4264 13716 4292 13892
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9600 13920 9628 13960
rect 10318 13948 10324 14000
rect 10376 13988 10382 14000
rect 16758 13988 16764 14000
rect 10376 13960 16764 13988
rect 10376 13948 10382 13960
rect 16758 13948 16764 13960
rect 16816 13948 16822 14000
rect 17218 13988 17224 14000
rect 17179 13960 17224 13988
rect 17218 13948 17224 13960
rect 17276 13948 17282 14000
rect 18874 13988 18880 14000
rect 18835 13960 18880 13988
rect 18874 13948 18880 13960
rect 18932 13948 18938 14000
rect 18966 13948 18972 14000
rect 19024 13988 19030 14000
rect 19024 13960 19069 13988
rect 19024 13948 19030 13960
rect 21266 13948 21272 14000
rect 21324 13988 21330 14000
rect 23308 13988 23336 14028
rect 23474 13988 23480 14000
rect 21324 13960 23336 13988
rect 23435 13960 23480 13988
rect 21324 13948 21330 13960
rect 23474 13948 23480 13960
rect 23532 13948 23538 14000
rect 24044 13997 24072 14028
rect 24489 14025 24501 14059
rect 24535 14056 24547 14059
rect 24946 14056 24952 14068
rect 24535 14028 24952 14056
rect 24535 14025 24547 14028
rect 24489 14019 24547 14025
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 26053 14059 26111 14065
rect 26053 14025 26065 14059
rect 26099 14056 26111 14059
rect 28258 14056 28264 14068
rect 26099 14028 27384 14056
rect 28219 14028 28264 14056
rect 26099 14025 26111 14028
rect 26053 14019 26111 14025
rect 24029 13991 24087 13997
rect 24029 13957 24041 13991
rect 24075 13957 24087 13991
rect 24029 13951 24087 13957
rect 15102 13920 15108 13932
rect 9600 13892 15108 13920
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15804 13892 15853 13920
rect 15804 13880 15810 13892
rect 15841 13889 15853 13892
rect 15887 13920 15899 13923
rect 16298 13920 16304 13932
rect 15887 13892 16304 13920
rect 15887 13889 15899 13892
rect 15841 13883 15899 13889
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 20898 13880 20904 13932
rect 20956 13920 20962 13932
rect 23014 13920 23020 13932
rect 20956 13892 23020 13920
rect 20956 13880 20962 13892
rect 23014 13880 23020 13892
rect 23072 13880 23078 13932
rect 4341 13855 4399 13861
rect 4341 13821 4353 13855
rect 4387 13852 4399 13855
rect 13998 13852 14004 13864
rect 4387 13824 14004 13852
rect 4387 13821 4399 13824
rect 4341 13815 4399 13821
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 14792 13824 16129 13852
rect 14792 13812 14798 13824
rect 16117 13821 16129 13824
rect 16163 13852 16175 13855
rect 16482 13852 16488 13864
rect 16163 13824 16488 13852
rect 16163 13821 16175 13824
rect 16117 13815 16175 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17586 13852 17592 13864
rect 17175 13824 17448 13852
rect 17547 13824 17592 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17420 13784 17448 13824
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 18230 13852 18236 13864
rect 17696 13824 18236 13852
rect 17696 13784 17724 13824
rect 18230 13812 18236 13824
rect 18288 13812 18294 13864
rect 19334 13852 19340 13864
rect 19295 13824 19340 13852
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19978 13852 19984 13864
rect 19939 13824 19984 13852
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 22186 13852 22192 13864
rect 22147 13824 22192 13852
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13852 22431 13855
rect 23382 13852 23388 13864
rect 22419 13824 23244 13852
rect 23343 13824 23388 13852
rect 22419 13821 22431 13824
rect 22373 13815 22431 13821
rect 17420 13756 17724 13784
rect 23216 13784 23244 13824
rect 23382 13812 23388 13824
rect 23440 13812 23446 13864
rect 24044 13852 24072 13951
rect 24670 13920 24676 13932
rect 24631 13892 24676 13920
rect 24670 13880 24676 13892
rect 24728 13880 24734 13932
rect 26237 13923 26295 13929
rect 26237 13889 26249 13923
rect 26283 13920 26295 13923
rect 26326 13920 26332 13932
rect 26283 13892 26332 13920
rect 26283 13889 26295 13892
rect 26237 13883 26295 13889
rect 26326 13880 26332 13892
rect 26384 13880 26390 13932
rect 27356 13929 27384 14028
rect 28258 14016 28264 14028
rect 28316 14016 28322 14068
rect 37090 14016 37096 14068
rect 37148 14056 37154 14068
rect 38105 14059 38163 14065
rect 38105 14056 38117 14059
rect 37148 14028 38117 14056
rect 37148 14016 37154 14028
rect 38105 14025 38117 14028
rect 38151 14025 38163 14059
rect 38105 14019 38163 14025
rect 27341 13923 27399 13929
rect 27341 13889 27353 13923
rect 27387 13889 27399 13923
rect 28442 13920 28448 13932
rect 28403 13892 28448 13920
rect 27341 13883 27399 13889
rect 28442 13880 28448 13892
rect 28500 13880 28506 13932
rect 38286 13920 38292 13932
rect 38247 13892 38292 13920
rect 38286 13880 38292 13892
rect 38344 13880 38350 13932
rect 26970 13852 26976 13864
rect 24044 13824 26976 13852
rect 26970 13812 26976 13824
rect 27028 13812 27034 13864
rect 23842 13784 23848 13796
rect 23216 13756 23848 13784
rect 23842 13744 23848 13756
rect 23900 13744 23906 13796
rect 27154 13716 27160 13728
rect 2902 13688 4292 13716
rect 27115 13688 27160 13716
rect 2902 13685 2914 13688
rect 2856 13679 2914 13685
rect 27154 13676 27160 13688
rect 27212 13676 27218 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 11514 13512 11520 13524
rect 11475 13484 11520 13512
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 12989 13515 13047 13521
rect 12989 13512 13001 13515
rect 12860 13484 13001 13512
rect 12860 13472 12866 13484
rect 12989 13481 13001 13484
rect 13035 13481 13047 13515
rect 12989 13475 13047 13481
rect 15841 13515 15899 13521
rect 15841 13481 15853 13515
rect 15887 13512 15899 13515
rect 17218 13512 17224 13524
rect 15887 13484 17224 13512
rect 15887 13481 15899 13484
rect 15841 13475 15899 13481
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 17954 13512 17960 13524
rect 17915 13484 17960 13512
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 23474 13472 23480 13524
rect 23532 13512 23538 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 23532 13484 24777 13512
rect 23532 13472 23538 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 29914 13512 29920 13524
rect 29875 13484 29920 13512
rect 24765 13475 24823 13481
rect 29914 13472 29920 13484
rect 29972 13472 29978 13524
rect 13998 13404 14004 13456
rect 14056 13444 14062 13456
rect 27798 13444 27804 13456
rect 14056 13416 27804 13444
rect 14056 13404 14062 13416
rect 27798 13404 27804 13416
rect 27856 13444 27862 13456
rect 30834 13444 30840 13456
rect 27856 13416 28396 13444
rect 30795 13416 30840 13444
rect 27856 13404 27862 13416
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 9766 13376 9772 13388
rect 9456 13348 9772 13376
rect 9456 13336 9462 13348
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 10042 13376 10048 13388
rect 9955 13348 10048 13376
rect 10042 13336 10048 13348
rect 10100 13376 10106 13388
rect 15562 13376 15568 13388
rect 10100 13348 15568 13376
rect 10100 13336 10106 13348
rect 15562 13336 15568 13348
rect 15620 13336 15626 13388
rect 19429 13379 19487 13385
rect 19429 13345 19441 13379
rect 19475 13376 19487 13379
rect 19978 13376 19984 13388
rect 19475 13348 19984 13376
rect 19475 13345 19487 13348
rect 19429 13339 19487 13345
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 23382 13376 23388 13388
rect 23343 13348 23388 13376
rect 23382 13336 23388 13348
rect 23440 13336 23446 13388
rect 26881 13379 26939 13385
rect 26881 13345 26893 13379
rect 26927 13376 26939 13379
rect 27154 13376 27160 13388
rect 26927 13348 27160 13376
rect 26927 13345 26939 13348
rect 26881 13339 26939 13345
rect 27154 13336 27160 13348
rect 27212 13336 27218 13388
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13308 1639 13311
rect 2682 13308 2688 13320
rect 1627 13280 2688 13308
rect 1627 13277 1639 13280
rect 1581 13271 1639 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 13446 13308 13452 13320
rect 12943 13280 13452 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 15010 13308 15016 13320
rect 14971 13280 15016 13308
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 15654 13268 15660 13320
rect 15712 13308 15718 13320
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 15712 13280 15761 13308
rect 15712 13268 15718 13280
rect 15749 13277 15761 13280
rect 15795 13277 15807 13311
rect 18138 13308 18144 13320
rect 18099 13280 18144 13308
rect 15749 13271 15807 13277
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13277 19671 13311
rect 21726 13308 21732 13320
rect 21687 13280 21732 13308
rect 19613 13271 19671 13277
rect 10502 13200 10508 13252
rect 10560 13200 10566 13252
rect 11422 13200 11428 13252
rect 11480 13240 11486 13252
rect 14458 13240 14464 13252
rect 11480 13212 14464 13240
rect 11480 13200 11486 13212
rect 14458 13200 14464 13212
rect 14516 13200 14522 13252
rect 19628 13240 19656 13271
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 24946 13308 24952 13320
rect 24907 13280 24952 13308
rect 24946 13268 24952 13280
rect 25004 13268 25010 13320
rect 26234 13268 26240 13320
rect 26292 13308 26298 13320
rect 26602 13308 26608 13320
rect 26292 13280 26608 13308
rect 26292 13268 26298 13280
rect 26602 13268 26608 13280
rect 26660 13308 26666 13320
rect 28368 13317 28396 13416
rect 30834 13404 30840 13416
rect 30892 13404 30898 13456
rect 30466 13376 30472 13388
rect 30427 13348 30472 13376
rect 30466 13336 30472 13348
rect 30524 13336 30530 13388
rect 36906 13376 36912 13388
rect 30576 13348 36912 13376
rect 26697 13311 26755 13317
rect 26697 13308 26709 13311
rect 26660 13280 26709 13308
rect 26660 13268 26666 13280
rect 26697 13277 26709 13280
rect 26743 13277 26755 13311
rect 26697 13271 26755 13277
rect 28353 13311 28411 13317
rect 28353 13277 28365 13311
rect 28399 13277 28411 13311
rect 28353 13271 28411 13277
rect 28997 13311 29055 13317
rect 28997 13277 29009 13311
rect 29043 13277 29055 13311
rect 28997 13271 29055 13277
rect 29825 13311 29883 13317
rect 29825 13277 29837 13311
rect 29871 13308 29883 13311
rect 30576 13308 30604 13348
rect 36906 13336 36912 13348
rect 36964 13336 36970 13388
rect 29871 13280 30604 13308
rect 30653 13311 30711 13317
rect 29871 13277 29883 13280
rect 29825 13271 29883 13277
rect 30653 13277 30665 13311
rect 30699 13277 30711 13311
rect 30653 13271 30711 13277
rect 23106 13240 23112 13252
rect 19628 13212 23112 13240
rect 23106 13200 23112 13212
rect 23164 13200 23170 13252
rect 29012 13240 29040 13271
rect 30668 13240 30696 13271
rect 28184 13212 29040 13240
rect 29840 13212 30696 13240
rect 1762 13172 1768 13184
rect 1723 13144 1768 13172
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 14550 13172 14556 13184
rect 13412 13144 14556 13172
rect 13412 13132 13418 13144
rect 14550 13132 14556 13144
rect 14608 13132 14614 13184
rect 15105 13175 15163 13181
rect 15105 13141 15117 13175
rect 15151 13172 15163 13175
rect 15194 13172 15200 13184
rect 15151 13144 15200 13172
rect 15151 13141 15163 13144
rect 15105 13135 15163 13141
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 20073 13175 20131 13181
rect 20073 13141 20085 13175
rect 20119 13172 20131 13175
rect 20806 13172 20812 13184
rect 20119 13144 20812 13172
rect 20119 13141 20131 13144
rect 20073 13135 20131 13141
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 20898 13132 20904 13184
rect 20956 13172 20962 13184
rect 21545 13175 21603 13181
rect 21545 13172 21557 13175
rect 20956 13144 21557 13172
rect 20956 13132 20962 13144
rect 21545 13141 21557 13144
rect 21591 13141 21603 13175
rect 21545 13135 21603 13141
rect 27341 13175 27399 13181
rect 27341 13141 27353 13175
rect 27387 13172 27399 13175
rect 28074 13172 28080 13184
rect 27387 13144 28080 13172
rect 27387 13141 27399 13144
rect 27341 13135 27399 13141
rect 28074 13132 28080 13144
rect 28132 13132 28138 13184
rect 28184 13181 28212 13212
rect 28169 13175 28227 13181
rect 28169 13141 28181 13175
rect 28215 13141 28227 13175
rect 28169 13135 28227 13141
rect 28813 13175 28871 13181
rect 28813 13141 28825 13175
rect 28859 13172 28871 13175
rect 29840 13172 29868 13212
rect 28859 13144 29868 13172
rect 28859 13141 28871 13144
rect 28813 13135 28871 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 7558 12968 7564 12980
rect 2792 12940 7564 12968
rect 2792 12909 2820 12940
rect 7558 12928 7564 12940
rect 7616 12968 7622 12980
rect 12342 12968 12348 12980
rect 7616 12940 12348 12968
rect 7616 12928 7622 12940
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 18693 12971 18751 12977
rect 18693 12937 18705 12971
rect 18739 12968 18751 12971
rect 18966 12968 18972 12980
rect 18739 12940 18972 12968
rect 18739 12937 18751 12940
rect 18693 12931 18751 12937
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 26421 12971 26479 12977
rect 26421 12968 26433 12971
rect 22112 12940 26433 12968
rect 2777 12903 2835 12909
rect 2777 12869 2789 12903
rect 2823 12869 2835 12903
rect 2777 12863 2835 12869
rect 3234 12860 3240 12912
rect 3292 12860 3298 12912
rect 10962 12900 10968 12912
rect 8418 12872 10968 12900
rect 10962 12860 10968 12872
rect 11020 12860 11026 12912
rect 13354 12900 13360 12912
rect 13315 12872 13360 12900
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 14734 12900 14740 12912
rect 14582 12872 14740 12900
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 16022 12900 16028 12912
rect 15983 12872 16028 12900
rect 16022 12860 16028 12872
rect 16080 12860 16086 12912
rect 17405 12903 17463 12909
rect 17405 12869 17417 12903
rect 17451 12900 17463 12903
rect 18598 12900 18604 12912
rect 17451 12872 18604 12900
rect 17451 12869 17463 12872
rect 17405 12863 17463 12869
rect 18598 12860 18604 12872
rect 18656 12860 18662 12912
rect 20898 12900 20904 12912
rect 20859 12872 20904 12900
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 22112 12909 22140 12940
rect 26421 12937 26433 12940
rect 26467 12937 26479 12971
rect 26421 12931 26479 12937
rect 29089 12971 29147 12977
rect 29089 12937 29101 12971
rect 29135 12968 29147 12971
rect 30834 12968 30840 12980
rect 29135 12940 30840 12968
rect 29135 12937 29147 12940
rect 29089 12931 29147 12937
rect 30834 12928 30840 12940
rect 30892 12928 30898 12980
rect 22097 12903 22155 12909
rect 22097 12869 22109 12903
rect 22143 12869 22155 12903
rect 22097 12863 22155 12869
rect 22189 12903 22247 12909
rect 22189 12869 22201 12903
rect 22235 12900 22247 12903
rect 23293 12903 23351 12909
rect 23293 12900 23305 12903
rect 22235 12872 23305 12900
rect 22235 12869 22247 12872
rect 22189 12863 22247 12869
rect 23293 12869 23305 12872
rect 23339 12869 23351 12903
rect 23293 12863 23351 12869
rect 24854 12860 24860 12912
rect 24912 12900 24918 12912
rect 24912 12872 25820 12900
rect 24912 12860 24918 12872
rect 25792 12844 25820 12872
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 9217 12835 9275 12841
rect 9217 12801 9229 12835
rect 9263 12832 9275 12835
rect 11606 12832 11612 12844
rect 9263 12804 11612 12832
rect 9263 12801 9275 12804
rect 9217 12795 9275 12801
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15746 12832 15752 12844
rect 15344 12804 15752 12832
rect 15344 12792 15350 12804
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 18874 12832 18880 12844
rect 18835 12804 18880 12832
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 23198 12832 23204 12844
rect 23159 12804 23204 12832
rect 23198 12792 23204 12804
rect 23256 12792 23262 12844
rect 24394 12832 24400 12844
rect 24355 12804 24400 12832
rect 24394 12792 24400 12804
rect 24452 12792 24458 12844
rect 25225 12835 25283 12841
rect 25225 12801 25237 12835
rect 25271 12832 25283 12835
rect 25271 12804 25728 12832
rect 25271 12801 25283 12804
rect 25225 12795 25283 12801
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12764 4307 12767
rect 6270 12764 6276 12776
rect 4295 12736 6276 12764
rect 4295 12733 4307 12736
rect 4249 12727 4307 12733
rect 6270 12724 6276 12736
rect 6328 12724 6334 12776
rect 6822 12724 6828 12776
rect 6880 12764 6886 12776
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 6880 12736 6929 12764
rect 6880 12724 6886 12736
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12764 7251 12767
rect 7239 12736 9674 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 8570 12588 8576 12640
rect 8628 12628 8634 12640
rect 8665 12631 8723 12637
rect 8665 12628 8677 12631
rect 8628 12600 8677 12628
rect 8628 12588 8634 12600
rect 8665 12597 8677 12600
rect 8711 12597 8723 12631
rect 9306 12628 9312 12640
rect 9267 12600 9312 12628
rect 8665 12591 8723 12597
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 9646 12628 9674 12736
rect 12894 12724 12900 12776
rect 12952 12764 12958 12776
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 12952 12736 13093 12764
rect 12952 12724 12958 12736
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 13504 12736 14412 12764
rect 13504 12724 13510 12736
rect 14384 12696 14412 12736
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 15105 12767 15163 12773
rect 15105 12764 15117 12767
rect 14608 12736 15117 12764
rect 14608 12724 14614 12736
rect 15105 12733 15117 12736
rect 15151 12733 15163 12767
rect 17310 12764 17316 12776
rect 17271 12736 17316 12764
rect 15105 12727 15163 12733
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 17586 12764 17592 12776
rect 17499 12736 17592 12764
rect 17586 12724 17592 12736
rect 17644 12724 17650 12776
rect 20806 12764 20812 12776
rect 20767 12736 20812 12764
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 21174 12764 21180 12776
rect 21135 12736 21180 12764
rect 21174 12724 21180 12736
rect 21232 12724 21238 12776
rect 22370 12764 22376 12776
rect 22331 12736 22376 12764
rect 22370 12724 22376 12736
rect 22428 12724 22434 12776
rect 16022 12696 16028 12708
rect 14384 12668 16028 12696
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 16942 12656 16948 12708
rect 17000 12696 17006 12708
rect 17604 12696 17632 12724
rect 17000 12668 17632 12696
rect 17000 12656 17006 12668
rect 23842 12656 23848 12708
rect 23900 12696 23906 12708
rect 25700 12705 25728 12804
rect 25774 12792 25780 12844
rect 25832 12832 25838 12844
rect 25869 12835 25927 12841
rect 25869 12832 25881 12835
rect 25832 12804 25881 12832
rect 25832 12792 25838 12804
rect 25869 12801 25881 12804
rect 25915 12801 25927 12835
rect 26326 12832 26332 12844
rect 26287 12804 26332 12832
rect 25869 12795 25927 12801
rect 26326 12792 26332 12804
rect 26384 12792 26390 12844
rect 26786 12792 26792 12844
rect 26844 12832 26850 12844
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 26844 12804 27169 12832
rect 26844 12792 26850 12804
rect 27157 12801 27169 12804
rect 27203 12801 27215 12835
rect 27798 12832 27804 12844
rect 27759 12804 27804 12832
rect 27157 12795 27215 12801
rect 27798 12792 27804 12804
rect 27856 12792 27862 12844
rect 27893 12835 27951 12841
rect 27893 12801 27905 12835
rect 27939 12832 27951 12835
rect 28629 12835 28687 12841
rect 28629 12832 28641 12835
rect 27939 12804 28641 12832
rect 27939 12801 27951 12804
rect 27893 12795 27951 12801
rect 28629 12801 28641 12804
rect 28675 12801 28687 12835
rect 28629 12795 28687 12801
rect 28074 12724 28080 12776
rect 28132 12764 28138 12776
rect 28445 12767 28503 12773
rect 28445 12764 28457 12767
rect 28132 12736 28457 12764
rect 28132 12724 28138 12736
rect 28445 12733 28457 12736
rect 28491 12733 28503 12767
rect 28445 12727 28503 12733
rect 25041 12699 25099 12705
rect 25041 12696 25053 12699
rect 23900 12668 25053 12696
rect 23900 12656 23906 12668
rect 25041 12665 25053 12668
rect 25087 12665 25099 12699
rect 25041 12659 25099 12665
rect 25685 12699 25743 12705
rect 25685 12665 25697 12699
rect 25731 12665 25743 12699
rect 25685 12659 25743 12665
rect 14642 12628 14648 12640
rect 9646 12600 14648 12628
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 24489 12631 24547 12637
rect 24489 12597 24501 12631
rect 24535 12628 24547 12631
rect 24946 12628 24952 12640
rect 24535 12600 24952 12628
rect 24535 12597 24547 12600
rect 24489 12591 24547 12597
rect 24946 12588 24952 12600
rect 25004 12588 25010 12640
rect 27246 12628 27252 12640
rect 27207 12600 27252 12628
rect 27246 12588 27252 12600
rect 27304 12588 27310 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 3234 12424 3240 12436
rect 3195 12396 3240 12424
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 16206 12424 16212 12436
rect 12216 12396 16212 12424
rect 12216 12384 12222 12396
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 18233 12427 18291 12433
rect 16632 12396 16677 12424
rect 16632 12384 16638 12396
rect 18233 12393 18245 12427
rect 18279 12424 18291 12427
rect 18874 12424 18880 12436
rect 18279 12396 18880 12424
rect 18279 12393 18291 12396
rect 18233 12387 18291 12393
rect 18874 12384 18880 12396
rect 18932 12384 18938 12436
rect 20806 12424 20812 12436
rect 20767 12396 20812 12424
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 21726 12384 21732 12436
rect 21784 12424 21790 12436
rect 22005 12427 22063 12433
rect 22005 12424 22017 12427
rect 21784 12396 22017 12424
rect 21784 12384 21790 12396
rect 22005 12393 22017 12396
rect 22051 12393 22063 12427
rect 22005 12387 22063 12393
rect 12618 12316 12624 12368
rect 12676 12356 12682 12368
rect 12676 12328 14412 12356
rect 12676 12316 12682 12328
rect 6362 12288 6368 12300
rect 6323 12260 6368 12288
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 13630 12288 13636 12300
rect 12759 12260 13636 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 13630 12248 13636 12260
rect 13688 12248 13694 12300
rect 14384 12288 14412 12328
rect 16040 12328 17540 12356
rect 15286 12288 15292 12300
rect 14384 12260 15292 12288
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12220 3203 12223
rect 3326 12220 3332 12232
rect 3191 12192 3332 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 5684 12192 6101 12220
rect 5684 12180 5690 12192
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 7926 12180 7932 12232
rect 7984 12220 7990 12232
rect 11701 12223 11759 12229
rect 11701 12220 11713 12223
rect 7984 12192 11713 12220
rect 7984 12180 7990 12192
rect 11701 12189 11713 12192
rect 11747 12189 11759 12223
rect 12618 12220 12624 12232
rect 12579 12192 12624 12220
rect 11701 12183 11759 12189
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 13504 12192 13553 12220
rect 13504 12180 13510 12192
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13872 12192 14289 12220
rect 13872 12180 13878 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 9306 12152 9312 12164
rect 7590 12124 9312 12152
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 14550 12152 14556 12164
rect 14511 12124 14556 12152
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 15194 12112 15200 12164
rect 15252 12112 15258 12164
rect 7834 12084 7840 12096
rect 7795 12056 7840 12084
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 11517 12087 11575 12093
rect 11517 12053 11529 12087
rect 11563 12084 11575 12087
rect 12802 12084 12808 12096
rect 11563 12056 12808 12084
rect 11563 12053 11575 12056
rect 11517 12047 11575 12053
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 13633 12087 13691 12093
rect 13633 12053 13645 12087
rect 13679 12084 13691 12087
rect 14918 12084 14924 12096
rect 13679 12056 14924 12084
rect 13679 12053 13691 12056
rect 13633 12047 13691 12053
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 16040 12093 16068 12328
rect 17310 12288 17316 12300
rect 17271 12260 17316 12288
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 16482 12220 16488 12232
rect 16443 12192 16488 12220
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 17512 12152 17540 12328
rect 17586 12316 17592 12368
rect 17644 12356 17650 12368
rect 27338 12356 27344 12368
rect 17644 12328 27344 12356
rect 17644 12316 17650 12328
rect 27338 12316 27344 12328
rect 27396 12316 27402 12368
rect 20349 12291 20407 12297
rect 20349 12257 20361 12291
rect 20395 12288 20407 12291
rect 21453 12291 21511 12297
rect 21453 12288 21465 12291
rect 20395 12260 21465 12288
rect 20395 12257 20407 12260
rect 20349 12251 20407 12257
rect 21453 12257 21465 12260
rect 21499 12257 21511 12291
rect 21453 12251 21511 12257
rect 22112 12260 25912 12288
rect 18414 12220 18420 12232
rect 18375 12192 18420 12220
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12220 20223 12223
rect 20438 12220 20444 12232
rect 20211 12192 20444 12220
rect 20211 12189 20223 12192
rect 20165 12183 20223 12189
rect 20438 12180 20444 12192
rect 20496 12180 20502 12232
rect 21358 12220 21364 12232
rect 21271 12192 21364 12220
rect 21358 12180 21364 12192
rect 21416 12220 21422 12232
rect 22112 12220 22140 12260
rect 21416 12192 22140 12220
rect 22189 12223 22247 12229
rect 21416 12180 21422 12192
rect 22189 12189 22201 12223
rect 22235 12189 22247 12223
rect 22189 12183 22247 12189
rect 23477 12223 23535 12229
rect 23477 12189 23489 12223
rect 23523 12220 23535 12223
rect 24394 12220 24400 12232
rect 23523 12192 24400 12220
rect 23523 12189 23535 12192
rect 23477 12183 23535 12189
rect 21634 12152 21640 12164
rect 17512 12124 21640 12152
rect 21634 12112 21640 12124
rect 21692 12152 21698 12164
rect 22204 12152 22232 12183
rect 24394 12180 24400 12192
rect 24452 12180 24458 12232
rect 25884 12229 25912 12260
rect 25869 12223 25927 12229
rect 25869 12189 25881 12223
rect 25915 12220 25927 12223
rect 26050 12220 26056 12232
rect 25915 12192 26056 12220
rect 25915 12189 25927 12192
rect 25869 12183 25927 12189
rect 26050 12180 26056 12192
rect 26108 12180 26114 12232
rect 30834 12180 30840 12232
rect 30892 12220 30898 12232
rect 32125 12223 32183 12229
rect 32125 12220 32137 12223
rect 30892 12192 32137 12220
rect 30892 12180 30898 12192
rect 32125 12189 32137 12192
rect 32171 12189 32183 12223
rect 32125 12183 32183 12189
rect 21692 12124 22232 12152
rect 21692 12112 21698 12124
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 15344 12056 16037 12084
rect 15344 12044 15350 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 16025 12047 16083 12053
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 22370 12084 22376 12096
rect 18196 12056 22376 12084
rect 18196 12044 18202 12056
rect 22370 12044 22376 12056
rect 22428 12044 22434 12096
rect 22649 12087 22707 12093
rect 22649 12053 22661 12087
rect 22695 12084 22707 12087
rect 23198 12084 23204 12096
rect 22695 12056 23204 12084
rect 22695 12053 22707 12056
rect 22649 12047 22707 12053
rect 23198 12044 23204 12056
rect 23256 12044 23262 12096
rect 23293 12087 23351 12093
rect 23293 12053 23305 12087
rect 23339 12084 23351 12087
rect 23566 12084 23572 12096
rect 23339 12056 23572 12084
rect 23339 12053 23351 12056
rect 23293 12047 23351 12053
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 25685 12087 25743 12093
rect 25685 12053 25697 12087
rect 25731 12084 25743 12087
rect 26142 12084 26148 12096
rect 25731 12056 26148 12084
rect 25731 12053 25743 12056
rect 25685 12047 25743 12053
rect 26142 12044 26148 12056
rect 26200 12044 26206 12096
rect 32217 12087 32275 12093
rect 32217 12053 32229 12087
rect 32263 12084 32275 12087
rect 32490 12084 32496 12096
rect 32263 12056 32496 12084
rect 32263 12053 32275 12056
rect 32217 12047 32275 12053
rect 32490 12044 32496 12056
rect 32548 12044 32554 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 5721 11883 5779 11889
rect 5721 11880 5733 11883
rect 5592 11852 5733 11880
rect 5592 11840 5598 11852
rect 5721 11849 5733 11852
rect 5767 11880 5779 11883
rect 5810 11880 5816 11892
rect 5767 11852 5816 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 10686 11880 10692 11892
rect 8404 11852 10692 11880
rect 6730 11812 6736 11824
rect 5474 11784 6736 11812
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 8404 11821 8432 11852
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 12894 11840 12900 11892
rect 12952 11840 12958 11892
rect 14734 11880 14740 11892
rect 14695 11852 14740 11880
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 16206 11880 16212 11892
rect 16167 11852 16212 11880
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 18138 11880 18144 11892
rect 17788 11852 18144 11880
rect 8389 11815 8447 11821
rect 8389 11781 8401 11815
rect 8435 11781 8447 11815
rect 12912 11812 12940 11840
rect 12912 11784 13584 11812
rect 8389 11775 8447 11781
rect 2498 11704 2504 11756
rect 2556 11744 2562 11756
rect 3970 11744 3976 11756
rect 2556 11716 3976 11744
rect 2556 11704 2562 11716
rect 3970 11704 3976 11716
rect 4028 11704 4034 11756
rect 6822 11704 6828 11756
rect 6880 11744 6886 11756
rect 6914 11744 6920 11756
rect 6880 11716 6920 11744
rect 6880 11704 6886 11716
rect 6914 11704 6920 11716
rect 6972 11744 6978 11756
rect 13556 11753 13584 11784
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 15381 11815 15439 11821
rect 15381 11812 15393 11815
rect 14516 11784 15393 11812
rect 14516 11772 14522 11784
rect 15381 11781 15393 11784
rect 15427 11781 15439 11815
rect 16482 11812 16488 11824
rect 15381 11775 15439 11781
rect 16132 11784 16488 11812
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 6972 11716 8125 11744
rect 6972 11704 6978 11716
rect 8113 11713 8125 11716
rect 8159 11713 8171 11747
rect 13541 11747 13599 11753
rect 8113 11707 8171 11713
rect 4249 11679 4307 11685
rect 4249 11645 4261 11679
rect 4295 11676 4307 11679
rect 7374 11676 7380 11688
rect 4295 11648 7380 11676
rect 4295 11645 4307 11648
rect 4249 11639 4307 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 9508 11608 9536 11730
rect 9582 11636 9588 11688
rect 9640 11676 9646 11688
rect 12176 11676 12204 11730
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 13814 11744 13820 11756
rect 13587 11716 13820 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 14645 11747 14703 11753
rect 14645 11713 14657 11747
rect 14691 11744 14703 11747
rect 15010 11744 15016 11756
rect 14691 11716 15016 11744
rect 14691 11713 14703 11716
rect 14645 11707 14703 11713
rect 15010 11704 15016 11716
rect 15068 11704 15074 11756
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11744 15347 11747
rect 15654 11744 15660 11756
rect 15335 11716 15660 11744
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 15654 11704 15660 11716
rect 15712 11744 15718 11756
rect 16132 11753 16160 11784
rect 16482 11772 16488 11784
rect 16540 11772 16546 11824
rect 17788 11821 17816 11852
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18414 11840 18420 11892
rect 18472 11880 18478 11892
rect 27062 11880 27068 11892
rect 18472 11852 27068 11880
rect 18472 11840 18478 11852
rect 27062 11840 27068 11852
rect 27120 11840 27126 11892
rect 27801 11883 27859 11889
rect 27801 11849 27813 11883
rect 27847 11880 27859 11883
rect 28074 11880 28080 11892
rect 27847 11852 28080 11880
rect 27847 11849 27859 11852
rect 27801 11843 27859 11849
rect 28074 11840 28080 11852
rect 28132 11840 28138 11892
rect 32398 11840 32404 11892
rect 32456 11880 32462 11892
rect 38105 11883 38163 11889
rect 38105 11880 38117 11883
rect 32456 11852 38117 11880
rect 32456 11840 32462 11852
rect 38105 11849 38117 11852
rect 38151 11849 38163 11883
rect 38105 11843 38163 11849
rect 17773 11815 17831 11821
rect 17773 11781 17785 11815
rect 17819 11781 17831 11815
rect 17773 11775 17831 11781
rect 17865 11815 17923 11821
rect 17865 11781 17877 11815
rect 17911 11812 17923 11815
rect 18230 11812 18236 11824
rect 17911 11784 18236 11812
rect 17911 11781 17923 11784
rect 17865 11775 17923 11781
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 18966 11812 18972 11824
rect 18927 11784 18972 11812
rect 18966 11772 18972 11784
rect 19024 11772 19030 11824
rect 19061 11815 19119 11821
rect 19061 11781 19073 11815
rect 19107 11812 19119 11815
rect 19978 11812 19984 11824
rect 19107 11784 19984 11812
rect 19107 11781 19119 11784
rect 19061 11775 19119 11781
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 25593 11815 25651 11821
rect 25593 11781 25605 11815
rect 25639 11812 25651 11815
rect 25958 11812 25964 11824
rect 25639 11784 25964 11812
rect 25639 11781 25651 11784
rect 25593 11775 25651 11781
rect 25958 11772 25964 11784
rect 26016 11772 26022 11824
rect 27706 11812 27712 11824
rect 26206 11784 27712 11812
rect 16117 11747 16175 11753
rect 16117 11744 16129 11747
rect 15712 11716 16129 11744
rect 15712 11704 15718 11716
rect 16117 11713 16129 11716
rect 16163 11713 16175 11747
rect 17586 11744 17592 11756
rect 16117 11707 16175 11713
rect 16546 11716 17592 11744
rect 9640 11648 12204 11676
rect 9640 11636 9646 11648
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 12584 11648 13277 11676
rect 12584 11636 12590 11648
rect 13265 11645 13277 11648
rect 13311 11676 13323 11679
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13311 11648 13921 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13909 11645 13921 11648
rect 13955 11676 13967 11679
rect 16546 11676 16574 11716
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11744 19671 11747
rect 20254 11744 20260 11756
rect 19659 11716 20260 11744
rect 19659 11713 19671 11716
rect 19613 11707 19671 11713
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 23198 11744 23204 11756
rect 23159 11716 23204 11744
rect 23198 11704 23204 11716
rect 23256 11704 23262 11756
rect 13955 11648 16574 11676
rect 17037 11679 17095 11685
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 17037 11645 17049 11679
rect 17083 11676 17095 11679
rect 17494 11676 17500 11688
rect 17083 11648 17500 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 17920 11648 18061 11676
rect 17920 11636 17926 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 21358 11676 21364 11688
rect 18049 11639 18107 11645
rect 18892 11648 21364 11676
rect 9508 11580 12296 11608
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 6822 11540 6828 11552
rect 6420 11512 6828 11540
rect 6420 11500 6426 11512
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 11606 11540 11612 11552
rect 9907 11512 11612 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 11606 11500 11612 11512
rect 11664 11500 11670 11552
rect 11790 11540 11796 11552
rect 11751 11512 11796 11540
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12268 11540 12296 11580
rect 13740 11580 14504 11608
rect 13740 11540 13768 11580
rect 12268 11512 13768 11540
rect 14476 11540 14504 11580
rect 14550 11568 14556 11620
rect 14608 11608 14614 11620
rect 18892 11608 18920 11648
rect 21358 11636 21364 11648
rect 21416 11636 21422 11688
rect 23382 11676 23388 11688
rect 23343 11648 23388 11676
rect 23382 11636 23388 11648
rect 23440 11636 23446 11688
rect 25501 11679 25559 11685
rect 25501 11645 25513 11679
rect 25547 11645 25559 11679
rect 25774 11676 25780 11688
rect 25735 11648 25780 11676
rect 25501 11639 25559 11645
rect 14608 11580 18920 11608
rect 14608 11568 14614 11580
rect 18966 11568 18972 11620
rect 19024 11608 19030 11620
rect 19024 11580 22968 11608
rect 19024 11568 19030 11580
rect 15286 11540 15292 11552
rect 14476 11512 15292 11540
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 16022 11540 16028 11552
rect 15436 11512 16028 11540
rect 15436 11500 15442 11512
rect 16022 11500 16028 11512
rect 16080 11540 16086 11552
rect 22646 11540 22652 11552
rect 16080 11512 22652 11540
rect 16080 11500 16086 11512
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 22940 11540 22968 11580
rect 23014 11568 23020 11620
rect 23072 11608 23078 11620
rect 23569 11611 23627 11617
rect 23569 11608 23581 11611
rect 23072 11580 23581 11608
rect 23072 11568 23078 11580
rect 23569 11577 23581 11580
rect 23615 11608 23627 11611
rect 25222 11608 25228 11620
rect 23615 11580 25228 11608
rect 23615 11577 23627 11580
rect 23569 11571 23627 11577
rect 25222 11568 25228 11580
rect 25280 11568 25286 11620
rect 25516 11608 25544 11639
rect 25774 11636 25780 11648
rect 25832 11676 25838 11688
rect 26206 11676 26234 11784
rect 27706 11772 27712 11784
rect 27764 11772 27770 11824
rect 27246 11704 27252 11756
rect 27304 11744 27310 11756
rect 27341 11747 27399 11753
rect 27341 11744 27353 11747
rect 27304 11716 27353 11744
rect 27304 11704 27310 11716
rect 27341 11713 27353 11716
rect 27387 11713 27399 11747
rect 32490 11744 32496 11756
rect 32451 11716 32496 11744
rect 27341 11707 27399 11713
rect 32490 11704 32496 11716
rect 32548 11704 32554 11756
rect 38286 11744 38292 11756
rect 38247 11716 38292 11744
rect 38286 11704 38292 11716
rect 38344 11704 38350 11756
rect 27154 11676 27160 11688
rect 25832 11648 26234 11676
rect 27067 11648 27160 11676
rect 25832 11636 25838 11648
rect 27154 11636 27160 11648
rect 27212 11676 27218 11688
rect 31754 11676 31760 11688
rect 27212 11648 31760 11676
rect 27212 11636 27218 11648
rect 31754 11636 31760 11648
rect 31812 11636 31818 11688
rect 25866 11608 25872 11620
rect 25516 11580 25872 11608
rect 25866 11568 25872 11580
rect 25924 11568 25930 11620
rect 25038 11540 25044 11552
rect 22940 11512 25044 11540
rect 25038 11500 25044 11512
rect 25096 11500 25102 11552
rect 32309 11543 32367 11549
rect 32309 11509 32321 11543
rect 32355 11540 32367 11543
rect 34054 11540 34060 11552
rect 32355 11512 34060 11540
rect 32355 11509 32367 11512
rect 32309 11503 32367 11509
rect 34054 11500 34060 11512
rect 34112 11500 34118 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 15749 11339 15807 11345
rect 15749 11336 15761 11339
rect 4120 11308 15761 11336
rect 4120 11296 4126 11308
rect 15749 11305 15761 11308
rect 15795 11305 15807 11339
rect 18414 11336 18420 11348
rect 15749 11299 15807 11305
rect 15856 11308 18420 11336
rect 6733 11271 6791 11277
rect 6733 11237 6745 11271
rect 6779 11268 6791 11271
rect 9214 11268 9220 11280
rect 6779 11240 9220 11268
rect 6779 11237 6791 11240
rect 6733 11231 6791 11237
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 11606 11228 11612 11280
rect 11664 11268 11670 11280
rect 14090 11268 14096 11280
rect 11664 11240 14096 11268
rect 11664 11228 11670 11240
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 15102 11268 15108 11280
rect 15063 11240 15108 11268
rect 15102 11228 15108 11240
rect 15160 11228 15166 11280
rect 1670 11160 1676 11212
rect 1728 11200 1734 11212
rect 1857 11203 1915 11209
rect 1857 11200 1869 11203
rect 1728 11172 1869 11200
rect 1728 11160 1734 11172
rect 1857 11169 1869 11172
rect 1903 11169 1915 11203
rect 1857 11163 1915 11169
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4985 11203 5043 11209
rect 4985 11200 4997 11203
rect 4028 11172 4997 11200
rect 4028 11160 4034 11172
rect 4985 11169 4997 11172
rect 5031 11200 5043 11203
rect 5626 11200 5632 11212
rect 5031 11172 5632 11200
rect 5031 11169 5043 11172
rect 4985 11163 5043 11169
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11200 10563 11203
rect 13722 11200 13728 11212
rect 10551 11172 13728 11200
rect 10551 11169 10563 11172
rect 10505 11163 10563 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 15856 11200 15884 11308
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 18598 11336 18604 11348
rect 18559 11308 18604 11336
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 23382 11336 23388 11348
rect 23343 11308 23388 11336
rect 23382 11296 23388 11308
rect 23440 11296 23446 11348
rect 25222 11336 25228 11348
rect 25183 11308 25228 11336
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 25958 11336 25964 11348
rect 25919 11308 25964 11336
rect 25958 11296 25964 11308
rect 26016 11296 26022 11348
rect 27522 11296 27528 11348
rect 27580 11336 27586 11348
rect 27801 11339 27859 11345
rect 27801 11336 27813 11339
rect 27580 11308 27813 11336
rect 27580 11296 27586 11308
rect 27801 11305 27813 11308
rect 27847 11305 27859 11339
rect 27801 11299 27859 11305
rect 25774 11268 25780 11280
rect 20548 11240 25780 11268
rect 14936 11172 15884 11200
rect 16577 11203 16635 11209
rect 1578 11132 1584 11144
rect 1539 11104 1584 11132
rect 1578 11092 1584 11104
rect 1636 11092 1642 11144
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 9824 11104 10241 11132
rect 9824 11092 9830 11104
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 14936 11132 14964 11172
rect 16577 11169 16589 11203
rect 16623 11200 16635 11203
rect 16666 11200 16672 11212
rect 16623 11172 16672 11200
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 16666 11160 16672 11172
rect 16724 11160 16730 11212
rect 17494 11200 17500 11212
rect 17455 11172 17500 11200
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 17678 11160 17684 11212
rect 17736 11200 17742 11212
rect 20548 11209 20576 11240
rect 25774 11228 25780 11240
rect 25832 11228 25838 11280
rect 20533 11203 20591 11209
rect 17736 11172 18828 11200
rect 17736 11160 17742 11172
rect 11848 11104 14964 11132
rect 11848 11092 11854 11104
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 15654 11132 15660 11144
rect 15068 11104 15113 11132
rect 15615 11104 15660 11132
rect 15068 11092 15074 11104
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 16301 11135 16359 11141
rect 16301 11132 16313 11135
rect 15896 11104 16313 11132
rect 15896 11092 15902 11104
rect 16301 11101 16313 11104
rect 16347 11132 16359 11135
rect 16482 11132 16488 11144
rect 16347 11104 16488 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 18800 11141 18828 11172
rect 20533 11169 20545 11203
rect 20579 11169 20591 11203
rect 20533 11163 20591 11169
rect 24946 11160 24952 11212
rect 25004 11200 25010 11212
rect 25041 11203 25099 11209
rect 25041 11200 25053 11203
rect 25004 11172 25053 11200
rect 25004 11160 25010 11172
rect 25041 11169 25053 11172
rect 25087 11169 25099 11203
rect 25041 11163 25099 11169
rect 26970 11160 26976 11212
rect 27028 11200 27034 11212
rect 27028 11172 31340 11200
rect 27028 11160 27034 11172
rect 18785 11135 18843 11141
rect 18785 11101 18797 11135
rect 18831 11101 18843 11135
rect 18785 11095 18843 11101
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 19484 11104 19625 11132
rect 19484 11092 19490 11104
rect 19613 11101 19625 11104
rect 19659 11101 19671 11135
rect 21634 11132 21640 11144
rect 21595 11104 21640 11132
rect 19613 11095 19671 11101
rect 21634 11092 21640 11104
rect 21692 11092 21698 11144
rect 22646 11092 22652 11144
rect 22704 11132 22710 11144
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 22704 11104 22753 11132
rect 22704 11092 22710 11104
rect 22741 11101 22753 11104
rect 22787 11101 22799 11135
rect 23566 11132 23572 11144
rect 23527 11104 23572 11132
rect 22741 11095 22799 11101
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5534 11064 5540 11076
rect 5307 11036 5540 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 5718 11024 5724 11076
rect 5776 11024 5782 11076
rect 12986 11064 12992 11076
rect 11730 11036 12992 11064
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 17586 11064 17592 11076
rect 17547 11036 17592 11064
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 17862 11024 17868 11076
rect 17920 11064 17926 11076
rect 18141 11067 18199 11073
rect 18141 11064 18153 11067
rect 17920 11036 18153 11064
rect 17920 11024 17926 11036
rect 18141 11033 18153 11036
rect 18187 11033 18199 11067
rect 18141 11027 18199 11033
rect 20625 11067 20683 11073
rect 20625 11033 20637 11067
rect 20671 11064 20683 11067
rect 21174 11064 21180 11076
rect 20671 11036 21036 11064
rect 21135 11036 21180 11064
rect 20671 11033 20683 11036
rect 20625 11027 20683 11033
rect 11514 10956 11520 11008
rect 11572 10996 11578 11008
rect 11977 10999 12035 11005
rect 11977 10996 11989 10999
rect 11572 10968 11989 10996
rect 11572 10956 11578 10968
rect 11977 10965 11989 10968
rect 12023 10965 12035 10999
rect 11977 10959 12035 10965
rect 19334 10956 19340 11008
rect 19392 10996 19398 11008
rect 19429 10999 19487 11005
rect 19429 10996 19441 10999
rect 19392 10968 19441 10996
rect 19392 10956 19398 10968
rect 19429 10965 19441 10968
rect 19475 10965 19487 10999
rect 21008 10996 21036 11036
rect 21174 11024 21180 11036
rect 21232 11024 21238 11076
rect 21729 11067 21787 11073
rect 21729 11064 21741 11067
rect 21284 11036 21741 11064
rect 21284 10996 21312 11036
rect 21729 11033 21741 11036
rect 21775 11033 21787 11067
rect 22756 11064 22784 11095
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 24857 11135 24915 11141
rect 24857 11101 24869 11135
rect 24903 11101 24915 11135
rect 26142 11132 26148 11144
rect 26103 11104 26148 11132
rect 24857 11095 24915 11101
rect 24762 11064 24768 11076
rect 22756 11036 24768 11064
rect 21729 11027 21787 11033
rect 24762 11024 24768 11036
rect 24820 11024 24826 11076
rect 24872 11064 24900 11095
rect 26142 11092 26148 11104
rect 26200 11092 26206 11144
rect 27709 11135 27767 11141
rect 27709 11101 27721 11135
rect 27755 11132 27767 11135
rect 29730 11132 29736 11144
rect 27755 11104 29736 11132
rect 27755 11101 27767 11104
rect 27709 11095 27767 11101
rect 29730 11092 29736 11104
rect 29788 11092 29794 11144
rect 31312 11141 31340 11172
rect 31297 11135 31355 11141
rect 31297 11101 31309 11135
rect 31343 11101 31355 11135
rect 31297 11095 31355 11101
rect 26694 11064 26700 11076
rect 24872 11036 26700 11064
rect 26694 11024 26700 11036
rect 26752 11024 26758 11076
rect 22830 10996 22836 11008
rect 21008 10968 21312 10996
rect 22791 10968 22836 10996
rect 19429 10959 19487 10965
rect 22830 10956 22836 10968
rect 22888 10956 22894 11008
rect 31386 10996 31392 11008
rect 31347 10968 31392 10996
rect 31386 10956 31392 10968
rect 31444 10956 31450 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 8754 10792 8760 10804
rect 8715 10764 8760 10792
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 9398 10752 9404 10804
rect 9456 10792 9462 10804
rect 15010 10792 15016 10804
rect 9456 10764 15016 10792
rect 9456 10752 9462 10764
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 16117 10795 16175 10801
rect 16117 10761 16129 10795
rect 16163 10792 16175 10795
rect 17678 10792 17684 10804
rect 16163 10764 17684 10792
rect 16163 10761 16175 10764
rect 16117 10755 16175 10761
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 18325 10795 18383 10801
rect 18325 10792 18337 10795
rect 18288 10764 18337 10792
rect 18288 10752 18294 10764
rect 18325 10761 18337 10764
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 36906 10752 36912 10804
rect 36964 10792 36970 10804
rect 38105 10795 38163 10801
rect 38105 10792 38117 10795
rect 36964 10764 38117 10792
rect 36964 10752 36970 10764
rect 38105 10761 38117 10764
rect 38151 10761 38163 10795
rect 38105 10755 38163 10761
rect 7558 10684 7564 10736
rect 7616 10724 7622 10736
rect 7616 10696 7774 10724
rect 7616 10684 7622 10696
rect 13998 10684 14004 10736
rect 14056 10724 14062 10736
rect 14056 10696 14582 10724
rect 14056 10684 14062 10696
rect 16206 10684 16212 10736
rect 16264 10724 16270 10736
rect 16482 10724 16488 10736
rect 16264 10696 16488 10724
rect 16264 10684 16270 10696
rect 16482 10684 16488 10696
rect 16540 10724 16546 10736
rect 16853 10727 16911 10733
rect 16853 10724 16865 10727
rect 16540 10696 16865 10724
rect 16540 10684 16546 10696
rect 16853 10693 16865 10696
rect 16899 10693 16911 10727
rect 19334 10724 19340 10736
rect 19295 10696 19340 10724
rect 16853 10687 16911 10693
rect 19334 10684 19340 10696
rect 19392 10684 19398 10736
rect 19889 10727 19947 10733
rect 19889 10693 19901 10727
rect 19935 10724 19947 10727
rect 20254 10724 20260 10736
rect 19935 10696 20260 10724
rect 19935 10693 19947 10696
rect 19889 10687 19947 10693
rect 20254 10684 20260 10696
rect 20312 10684 20318 10736
rect 26050 10724 26056 10736
rect 24228 10696 26056 10724
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 4614 10656 4620 10668
rect 1627 10628 4620 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 5684 10628 7021 10656
rect 5684 10616 5690 10628
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 13814 10656 13820 10668
rect 13775 10628 13820 10656
rect 7009 10619 7067 10625
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 15746 10616 15752 10668
rect 15804 10656 15810 10668
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 15804 10628 16313 10656
rect 15804 10616 15810 10628
rect 16301 10625 16313 10628
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 17494 10616 17500 10668
rect 17552 10656 17558 10668
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 17552 10628 18245 10656
rect 17552 10616 17558 10628
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 22830 10616 22836 10668
rect 22888 10656 22894 10668
rect 24228 10665 24256 10696
rect 26050 10684 26056 10696
rect 26108 10684 26114 10736
rect 23109 10659 23167 10665
rect 23109 10656 23121 10659
rect 22888 10628 23121 10656
rect 22888 10616 22894 10628
rect 23109 10625 23121 10628
rect 23155 10625 23167 10659
rect 23109 10619 23167 10625
rect 24213 10659 24271 10665
rect 24213 10625 24225 10659
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 24673 10659 24731 10665
rect 24673 10625 24685 10659
rect 24719 10625 24731 10659
rect 24673 10619 24731 10625
rect 7282 10588 7288 10600
rect 7195 10560 7288 10588
rect 7282 10548 7288 10560
rect 7340 10588 7346 10600
rect 11422 10588 11428 10600
rect 7340 10560 11428 10588
rect 7340 10548 7346 10560
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 14090 10588 14096 10600
rect 14051 10560 14096 10588
rect 14090 10548 14096 10560
rect 14148 10548 14154 10600
rect 14826 10548 14832 10600
rect 14884 10588 14890 10600
rect 17589 10591 17647 10597
rect 17589 10588 17601 10591
rect 14884 10560 17601 10588
rect 14884 10548 14890 10560
rect 17589 10557 17601 10560
rect 17635 10557 17647 10591
rect 17589 10551 17647 10557
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 16574 10480 16580 10532
rect 16632 10520 16638 10532
rect 17402 10520 17408 10532
rect 16632 10492 17408 10520
rect 16632 10480 16638 10492
rect 17402 10480 17408 10492
rect 17460 10520 17466 10532
rect 19260 10520 19288 10551
rect 22738 10548 22744 10600
rect 22796 10588 22802 10600
rect 22925 10591 22983 10597
rect 22925 10588 22937 10591
rect 22796 10560 22937 10588
rect 22796 10548 22802 10560
rect 22925 10557 22937 10560
rect 22971 10557 22983 10591
rect 24688 10588 24716 10619
rect 24762 10616 24768 10668
rect 24820 10656 24826 10668
rect 25501 10659 25559 10665
rect 25501 10656 25513 10659
rect 24820 10628 25513 10656
rect 24820 10616 24826 10628
rect 25501 10625 25513 10628
rect 25547 10625 25559 10659
rect 25501 10619 25559 10625
rect 27157 10659 27215 10665
rect 27157 10625 27169 10659
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 24946 10588 24952 10600
rect 24688 10560 24952 10588
rect 22925 10551 22983 10557
rect 24946 10548 24952 10560
rect 25004 10588 25010 10600
rect 25682 10588 25688 10600
rect 25004 10560 25688 10588
rect 25004 10548 25010 10560
rect 25682 10548 25688 10560
rect 25740 10548 25746 10600
rect 27172 10588 27200 10619
rect 27614 10616 27620 10668
rect 27672 10656 27678 10668
rect 30837 10659 30895 10665
rect 30837 10656 30849 10659
rect 27672 10628 30849 10656
rect 27672 10616 27678 10628
rect 30837 10625 30849 10628
rect 30883 10625 30895 10659
rect 38286 10656 38292 10668
rect 38247 10628 38292 10656
rect 30837 10619 30895 10625
rect 38286 10616 38292 10628
rect 38344 10616 38350 10668
rect 32306 10588 32312 10600
rect 27172 10560 32312 10588
rect 32306 10548 32312 10560
rect 32364 10548 32370 10600
rect 17460 10492 19288 10520
rect 17460 10480 17466 10492
rect 25866 10480 25872 10532
rect 25924 10520 25930 10532
rect 27249 10523 27307 10529
rect 27249 10520 27261 10523
rect 25924 10492 27261 10520
rect 25924 10480 25930 10492
rect 27249 10489 27261 10492
rect 27295 10489 27307 10523
rect 27249 10483 27307 10489
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 15562 10452 15568 10464
rect 9732 10424 15568 10452
rect 9732 10412 9738 10424
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 23566 10452 23572 10464
rect 23527 10424 23572 10452
rect 23566 10412 23572 10424
rect 23624 10412 23630 10464
rect 24026 10452 24032 10464
rect 23987 10424 24032 10452
rect 24026 10412 24032 10424
rect 24084 10412 24090 10464
rect 24765 10455 24823 10461
rect 24765 10421 24777 10455
rect 24811 10452 24823 10455
rect 24854 10452 24860 10464
rect 24811 10424 24860 10452
rect 24811 10421 24823 10424
rect 24765 10415 24823 10421
rect 24854 10412 24860 10424
rect 24912 10412 24918 10464
rect 25314 10452 25320 10464
rect 25275 10424 25320 10452
rect 25314 10412 25320 10424
rect 25372 10412 25378 10464
rect 30929 10455 30987 10461
rect 30929 10421 30941 10455
rect 30975 10452 30987 10455
rect 33134 10452 33140 10464
rect 30975 10424 33140 10452
rect 30975 10421 30987 10424
rect 30929 10415 30987 10421
rect 33134 10412 33140 10424
rect 33192 10412 33198 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 4065 10251 4123 10257
rect 4065 10248 4077 10251
rect 3936 10220 4077 10248
rect 3936 10208 3942 10220
rect 4065 10217 4077 10220
rect 4111 10217 4123 10251
rect 8570 10248 8576 10260
rect 4065 10211 4123 10217
rect 6886 10220 8576 10248
rect 3329 10183 3387 10189
rect 3329 10149 3341 10183
rect 3375 10180 3387 10183
rect 4982 10180 4988 10192
rect 3375 10152 4988 10180
rect 3375 10149 3387 10152
rect 3329 10143 3387 10149
rect 4982 10140 4988 10152
rect 5040 10140 5046 10192
rect 1578 10112 1584 10124
rect 1491 10084 1584 10112
rect 1578 10072 1584 10084
rect 1636 10112 1642 10124
rect 2498 10112 2504 10124
rect 1636 10084 2504 10112
rect 1636 10072 1642 10084
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 6886 10112 6914 10220
rect 8570 10208 8576 10220
rect 8628 10248 8634 10260
rect 15470 10248 15476 10260
rect 8628 10220 15476 10248
rect 8628 10208 8634 10220
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 17586 10208 17592 10260
rect 17644 10248 17650 10260
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 17644 10220 17785 10248
rect 17644 10208 17650 10220
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 18601 10251 18659 10257
rect 18601 10217 18613 10251
rect 18647 10248 18659 10251
rect 19426 10248 19432 10260
rect 18647 10220 19432 10248
rect 18647 10217 18659 10220
rect 18601 10211 18659 10217
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 23106 10248 23112 10260
rect 23067 10220 23112 10248
rect 23106 10208 23112 10220
rect 23164 10208 23170 10260
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 11572 10152 18828 10180
rect 11572 10140 11578 10152
rect 3252 10084 6914 10112
rect 7469 10115 7527 10121
rect 1857 9979 1915 9985
rect 1857 9945 1869 9979
rect 1903 9945 1915 9979
rect 3142 9976 3148 9988
rect 3082 9948 3148 9976
rect 1857 9939 1915 9945
rect 1872 9908 1900 9939
rect 3142 9936 3148 9948
rect 3200 9936 3206 9988
rect 3252 9908 3280 10084
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 12342 10112 12348 10124
rect 7515 10084 12348 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 15010 10072 15016 10124
rect 15068 10112 15074 10124
rect 17129 10115 17187 10121
rect 17129 10112 17141 10115
rect 15068 10084 17141 10112
rect 15068 10072 15074 10084
rect 17129 10081 17141 10084
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 3326 10004 3332 10056
rect 3384 10044 3390 10056
rect 3970 10044 3976 10056
rect 3384 10016 3976 10044
rect 3384 10004 3390 10016
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 5460 9976 5488 10007
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 9861 10047 9919 10053
rect 9861 10044 9873 10047
rect 9824 10016 9873 10044
rect 9824 10004 9830 10016
rect 9861 10013 9873 10016
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 11422 10004 11428 10056
rect 11480 10044 11486 10056
rect 17954 10044 17960 10056
rect 11480 10016 16574 10044
rect 17915 10016 17960 10044
rect 11480 10004 11486 10016
rect 5626 9976 5632 9988
rect 5460 9948 5632 9976
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 5721 9979 5779 9985
rect 5721 9945 5733 9979
rect 5767 9945 5779 9979
rect 5721 9939 5779 9945
rect 1872 9880 3280 9908
rect 5736 9908 5764 9939
rect 6270 9936 6276 9988
rect 6328 9936 6334 9988
rect 10134 9976 10140 9988
rect 10095 9948 10140 9976
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 13262 9976 13268 9988
rect 11362 9948 13268 9976
rect 13262 9936 13268 9948
rect 13320 9936 13326 9988
rect 16206 9936 16212 9988
rect 16264 9976 16270 9988
rect 16393 9979 16451 9985
rect 16393 9976 16405 9979
rect 16264 9948 16405 9976
rect 16264 9936 16270 9948
rect 16393 9945 16405 9948
rect 16439 9945 16451 9979
rect 16546 9976 16574 10016
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 18800 10053 18828 10152
rect 20070 10112 20076 10124
rect 19983 10084 20076 10112
rect 20070 10072 20076 10084
rect 20128 10112 20134 10124
rect 20438 10112 20444 10124
rect 20128 10084 20444 10112
rect 20128 10072 20134 10084
rect 20438 10072 20444 10084
rect 20496 10072 20502 10124
rect 24854 10112 24860 10124
rect 24815 10084 24860 10112
rect 24854 10072 24860 10084
rect 24912 10072 24918 10124
rect 26510 10112 26516 10124
rect 26471 10084 26516 10112
rect 26510 10072 26516 10084
rect 26568 10072 26574 10124
rect 18785 10047 18843 10053
rect 18785 10013 18797 10047
rect 18831 10044 18843 10047
rect 19242 10044 19248 10056
rect 18831 10016 19248 10044
rect 18831 10013 18843 10016
rect 18785 10007 18843 10013
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 20257 10047 20315 10053
rect 20257 10013 20269 10047
rect 20303 10044 20315 10047
rect 20806 10044 20812 10056
rect 20303 10016 20812 10044
rect 20303 10013 20315 10016
rect 20257 10007 20315 10013
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 21729 10047 21787 10053
rect 21729 10013 21741 10047
rect 21775 10013 21787 10047
rect 21910 10044 21916 10056
rect 21871 10016 21916 10044
rect 21729 10007 21787 10013
rect 18322 9976 18328 9988
rect 16546 9948 18328 9976
rect 16393 9939 16451 9945
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 21744 9976 21772 10007
rect 21910 10004 21916 10016
rect 21968 10004 21974 10056
rect 23293 10047 23351 10053
rect 23293 10013 23305 10047
rect 23339 10044 23351 10047
rect 24026 10044 24032 10056
rect 23339 10016 24032 10044
rect 23339 10013 23351 10016
rect 23293 10007 23351 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 24670 10044 24676 10056
rect 24631 10016 24676 10044
rect 24670 10004 24676 10016
rect 24728 10004 24734 10056
rect 31386 10044 31392 10056
rect 31347 10016 31392 10044
rect 31386 10004 31392 10016
rect 31444 10004 31450 10056
rect 33134 10044 33140 10056
rect 33095 10016 33140 10044
rect 33134 10004 33140 10016
rect 33192 10004 33198 10056
rect 25866 9976 25872 9988
rect 21744 9948 25872 9976
rect 25866 9936 25872 9948
rect 25924 9936 25930 9988
rect 25961 9979 26019 9985
rect 25961 9945 25973 9979
rect 26007 9976 26019 9979
rect 26234 9976 26240 9988
rect 26007 9948 26240 9976
rect 26007 9945 26019 9948
rect 25961 9939 26019 9945
rect 26234 9936 26240 9948
rect 26292 9936 26298 9988
rect 6362 9908 6368 9920
rect 5736 9880 6368 9908
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 11609 9911 11667 9917
rect 11609 9877 11621 9911
rect 11655 9908 11667 9911
rect 11974 9908 11980 9920
rect 11655 9880 11980 9908
rect 11655 9877 11667 9880
rect 11609 9871 11667 9877
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 17494 9908 17500 9920
rect 13780 9880 17500 9908
rect 13780 9868 13786 9880
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 20254 9868 20260 9920
rect 20312 9908 20318 9920
rect 20717 9911 20775 9917
rect 20717 9908 20729 9911
rect 20312 9880 20729 9908
rect 20312 9868 20318 9880
rect 20717 9877 20729 9880
rect 20763 9877 20775 9911
rect 22370 9908 22376 9920
rect 22331 9880 22376 9908
rect 20717 9871 20775 9877
rect 22370 9868 22376 9880
rect 22428 9868 22434 9920
rect 25317 9911 25375 9917
rect 25317 9877 25329 9911
rect 25363 9908 25375 9911
rect 25498 9908 25504 9920
rect 25363 9880 25504 9908
rect 25363 9877 25375 9880
rect 25317 9871 25375 9877
rect 25498 9868 25504 9880
rect 25556 9868 25562 9920
rect 31205 9911 31263 9917
rect 31205 9877 31217 9911
rect 31251 9908 31263 9911
rect 32858 9908 32864 9920
rect 31251 9880 32864 9908
rect 31251 9877 31263 9880
rect 31205 9871 31263 9877
rect 32858 9868 32864 9880
rect 32916 9868 32922 9920
rect 32953 9911 33011 9917
rect 32953 9877 32965 9911
rect 32999 9908 33011 9911
rect 38010 9908 38016 9920
rect 32999 9880 38016 9908
rect 32999 9877 33011 9880
rect 32953 9871 33011 9877
rect 38010 9868 38016 9880
rect 38068 9868 38074 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 4172 9676 6132 9704
rect 3786 9636 3792 9648
rect 3082 9608 3792 9636
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 4172 9636 4200 9676
rect 3896 9608 4200 9636
rect 1578 9568 1584 9580
rect 1539 9540 1584 9568
rect 1578 9528 1584 9540
rect 1636 9528 1642 9580
rect 3896 9577 3924 9608
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 5994 9568 6000 9580
rect 5290 9540 6000 9568
rect 3881 9531 3939 9537
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6104 9568 6132 9676
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 9674 9704 9680 9716
rect 6420 9676 9680 9704
rect 6420 9664 6426 9676
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 9824 9676 10732 9704
rect 9824 9664 9830 9676
rect 9030 9636 9036 9648
rect 8326 9608 9036 9636
rect 9030 9596 9036 9608
rect 9088 9596 9094 9648
rect 9784 9636 9812 9664
rect 9140 9608 9812 9636
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6104 9540 6837 9568
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 1854 9500 1860 9512
rect 1815 9472 1860 9500
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 6454 9500 6460 9512
rect 4203 9472 6460 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 6454 9460 6460 9472
rect 6512 9460 6518 9512
rect 3326 9364 3332 9376
rect 3287 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 5626 9364 5632 9376
rect 5587 9336 5632 9364
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 6840 9364 6868 9531
rect 7101 9503 7159 9509
rect 7101 9469 7113 9503
rect 7147 9500 7159 9503
rect 8386 9500 8392 9512
rect 7147 9472 8392 9500
rect 7147 9469 7159 9472
rect 7101 9463 7159 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 9140 9509 9168 9608
rect 10704 9568 10732 9676
rect 17052 9676 17540 9704
rect 10778 9596 10784 9648
rect 10836 9636 10842 9648
rect 11149 9639 11207 9645
rect 11149 9636 11161 9639
rect 10836 9608 11161 9636
rect 10836 9596 10842 9608
rect 11149 9605 11161 9608
rect 11195 9605 11207 9639
rect 11149 9599 11207 9605
rect 12526 9596 12532 9648
rect 12584 9596 12590 9648
rect 14918 9596 14924 9648
rect 14976 9596 14982 9648
rect 15746 9596 15752 9648
rect 15804 9636 15810 9648
rect 16666 9636 16672 9648
rect 15804 9608 16672 9636
rect 15804 9596 15810 9608
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 10534 9540 10640 9568
rect 10704 9540 11713 9568
rect 9125 9503 9183 9509
rect 9125 9500 9137 9503
rect 8496 9472 9137 9500
rect 6914 9364 6920 9376
rect 6840 9336 6920 9364
rect 6914 9324 6920 9336
rect 6972 9364 6978 9376
rect 8496 9364 8524 9472
rect 9125 9469 9137 9472
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 10612 9500 10640 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 13814 9528 13820 9580
rect 13872 9568 13878 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13872 9540 14197 9568
rect 13872 9528 13878 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 16942 9568 16948 9580
rect 15988 9540 16948 9568
rect 15988 9528 15994 9540
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 11974 9500 11980 9512
rect 9447 9472 10456 9500
rect 10612 9472 11836 9500
rect 11935 9472 11980 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 6972 9336 8524 9364
rect 8573 9367 8631 9373
rect 6972 9324 6978 9336
rect 8573 9333 8585 9367
rect 8619 9364 8631 9367
rect 10042 9364 10048 9376
rect 8619 9336 10048 9364
rect 8619 9333 8631 9336
rect 8573 9327 8631 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10428 9364 10456 9472
rect 11514 9364 11520 9376
rect 10428 9336 11520 9364
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 11808 9364 11836 9472
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 13722 9500 13728 9512
rect 13635 9472 13728 9500
rect 13722 9460 13728 9472
rect 13780 9500 13786 9512
rect 14461 9503 14519 9509
rect 13780 9472 14320 9500
rect 13780 9460 13786 9472
rect 13170 9364 13176 9376
rect 11808 9336 13176 9364
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 14292 9364 14320 9472
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 17052 9500 17080 9676
rect 17313 9639 17371 9645
rect 17313 9605 17325 9639
rect 17359 9636 17371 9639
rect 17402 9636 17408 9648
rect 17359 9608 17408 9636
rect 17359 9605 17371 9608
rect 17313 9599 17371 9605
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 17512 9636 17540 9676
rect 23566 9664 23572 9716
rect 23624 9704 23630 9716
rect 24673 9707 24731 9713
rect 24673 9704 24685 9707
rect 23624 9676 24685 9704
rect 23624 9664 23630 9676
rect 24673 9673 24685 9676
rect 24719 9704 24731 9707
rect 24762 9704 24768 9716
rect 24719 9676 24768 9704
rect 24719 9673 24731 9676
rect 24673 9667 24731 9673
rect 24762 9664 24768 9676
rect 24820 9664 24826 9716
rect 26234 9664 26240 9716
rect 26292 9704 26298 9716
rect 27157 9707 27215 9713
rect 27157 9704 27169 9707
rect 26292 9676 27169 9704
rect 26292 9664 26298 9676
rect 27157 9673 27169 9676
rect 27203 9673 27215 9707
rect 27157 9667 27215 9673
rect 18230 9636 18236 9648
rect 17512 9608 18236 9636
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 19334 9636 19340 9648
rect 18340 9608 19340 9636
rect 18340 9577 18368 9608
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 19705 9639 19763 9645
rect 19705 9605 19717 9639
rect 19751 9636 19763 9639
rect 19978 9636 19984 9648
rect 19751 9608 19984 9636
rect 19751 9605 19763 9608
rect 19705 9599 19763 9605
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 25498 9636 25504 9648
rect 20456 9608 22048 9636
rect 18325 9571 18383 9577
rect 18325 9537 18337 9571
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 18800 9540 19196 9568
rect 17218 9500 17224 9512
rect 14507 9472 17080 9500
rect 17179 9472 17224 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 17310 9460 17316 9512
rect 17368 9500 17374 9512
rect 17497 9503 17555 9509
rect 17497 9500 17509 9503
rect 17368 9472 17509 9500
rect 17368 9460 17374 9472
rect 17497 9469 17509 9472
rect 17543 9469 17555 9503
rect 18800 9500 18828 9540
rect 18966 9500 18972 9512
rect 17880 9488 18828 9500
rect 17497 9463 17555 9469
rect 17696 9472 18828 9488
rect 18927 9472 18972 9500
rect 17696 9460 17908 9472
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 19168 9500 19196 9540
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 19613 9571 19671 9577
rect 19613 9568 19625 9571
rect 19300 9540 19625 9568
rect 19300 9528 19306 9540
rect 19613 9537 19625 9540
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 20456 9500 20484 9608
rect 22020 9577 22048 9608
rect 24044 9608 25504 9636
rect 22005 9571 22063 9577
rect 22005 9537 22017 9571
rect 22051 9568 22063 9571
rect 23014 9568 23020 9580
rect 22051 9540 23020 9568
rect 22051 9537 22063 9540
rect 22005 9531 22063 9537
rect 23014 9528 23020 9540
rect 23072 9528 23078 9580
rect 24044 9577 24072 9608
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 29089 9639 29147 9645
rect 29089 9605 29101 9639
rect 29135 9636 29147 9639
rect 29546 9636 29552 9648
rect 29135 9608 29552 9636
rect 29135 9605 29147 9608
rect 29089 9599 29147 9605
rect 29546 9596 29552 9608
rect 29604 9596 29610 9648
rect 24029 9571 24087 9577
rect 24029 9537 24041 9571
rect 24075 9537 24087 9571
rect 25314 9568 25320 9580
rect 25275 9540 25320 9568
rect 24029 9531 24087 9537
rect 25314 9528 25320 9540
rect 25372 9528 25378 9580
rect 27341 9571 27399 9577
rect 27341 9537 27353 9571
rect 27387 9568 27399 9571
rect 27387 9540 27844 9568
rect 27387 9537 27399 9540
rect 27341 9531 27399 9537
rect 20622 9500 20628 9512
rect 19168 9472 20484 9500
rect 20583 9472 20628 9500
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 20809 9503 20867 9509
rect 20809 9500 20821 9503
rect 20772 9472 20821 9500
rect 20772 9460 20778 9472
rect 20809 9469 20821 9472
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 22741 9503 22799 9509
rect 22741 9469 22753 9503
rect 22787 9500 22799 9503
rect 23198 9500 23204 9512
rect 22787 9472 23204 9500
rect 22787 9469 22799 9472
rect 22741 9463 22799 9469
rect 23198 9460 23204 9472
rect 23256 9460 23262 9512
rect 24213 9503 24271 9509
rect 24213 9469 24225 9503
rect 24259 9500 24271 9503
rect 24259 9472 25176 9500
rect 24259 9469 24271 9472
rect 24213 9463 24271 9469
rect 15562 9392 15568 9444
rect 15620 9432 15626 9444
rect 17696 9432 17724 9460
rect 15620 9404 17724 9432
rect 18417 9435 18475 9441
rect 15620 9392 15626 9404
rect 18417 9401 18429 9435
rect 18463 9432 18475 9435
rect 20530 9432 20536 9444
rect 18463 9404 20536 9432
rect 18463 9401 18475 9404
rect 18417 9395 18475 9401
rect 20530 9392 20536 9404
rect 20588 9392 20594 9444
rect 25148 9441 25176 9472
rect 27816 9441 27844 9540
rect 27890 9528 27896 9580
rect 27948 9568 27954 9580
rect 27985 9571 28043 9577
rect 27985 9568 27997 9571
rect 27948 9540 27997 9568
rect 27948 9528 27954 9540
rect 27985 9537 27997 9540
rect 28031 9537 28043 9571
rect 27985 9531 28043 9537
rect 28997 9571 29055 9577
rect 28997 9537 29009 9571
rect 29043 9568 29055 9571
rect 33042 9568 33048 9580
rect 29043 9540 33048 9568
rect 29043 9537 29055 9540
rect 28997 9531 29055 9537
rect 33042 9528 33048 9540
rect 33100 9528 33106 9580
rect 25133 9435 25191 9441
rect 25133 9401 25145 9435
rect 25179 9401 25191 9435
rect 25133 9395 25191 9401
rect 27801 9435 27859 9441
rect 27801 9401 27813 9435
rect 27847 9401 27859 9435
rect 27801 9395 27859 9401
rect 15838 9364 15844 9376
rect 14292 9336 15844 9364
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 15933 9367 15991 9373
rect 15933 9333 15945 9367
rect 15979 9364 15991 9367
rect 16022 9364 16028 9376
rect 15979 9336 16028 9364
rect 15979 9333 15991 9336
rect 15933 9327 15991 9333
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17770 9364 17776 9376
rect 16816 9336 17776 9364
rect 16816 9324 16822 9336
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 18046 9324 18052 9376
rect 18104 9364 18110 9376
rect 20714 9364 20720 9376
rect 18104 9336 20720 9364
rect 18104 9324 18110 9336
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 20990 9364 20996 9376
rect 20951 9336 20996 9364
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 22094 9364 22100 9376
rect 22055 9336 22100 9364
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 4614 9160 4620 9172
rect 4571 9132 4620 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 5442 9160 5448 9172
rect 5403 9132 5448 9160
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6730 9160 6736 9172
rect 6691 9132 6736 9160
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 17129 9163 17187 9169
rect 6880 9132 16574 9160
rect 6880 9120 6886 9132
rect 1854 9052 1860 9104
rect 1912 9092 1918 9104
rect 11790 9092 11796 9104
rect 1912 9064 11796 9092
rect 1912 9052 1918 9064
rect 11790 9052 11796 9064
rect 11848 9052 11854 9104
rect 15102 9092 15108 9104
rect 14016 9064 15108 9092
rect 7837 9027 7895 9033
rect 7837 9024 7849 9027
rect 4724 8996 7849 9024
rect 4724 8965 4752 8996
rect 7837 8993 7849 8996
rect 7883 8993 7895 9027
rect 7837 8987 7895 8993
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 14016 9024 14044 9064
rect 15102 9052 15108 9064
rect 15160 9052 15166 9104
rect 15286 9092 15292 9104
rect 15247 9064 15292 9092
rect 15286 9052 15292 9064
rect 15344 9052 15350 9104
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 16390 9092 16396 9104
rect 15436 9064 16396 9092
rect 15436 9052 15442 9064
rect 16390 9052 16396 9064
rect 16448 9052 16454 9104
rect 16546 9092 16574 9132
rect 17129 9129 17141 9163
rect 17175 9160 17187 9163
rect 17954 9160 17960 9172
rect 17175 9132 17960 9160
rect 17175 9129 17187 9132
rect 17129 9123 17187 9129
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 18230 9120 18236 9172
rect 18288 9160 18294 9172
rect 24946 9160 24952 9172
rect 18288 9132 20852 9160
rect 18288 9120 18294 9132
rect 16942 9092 16948 9104
rect 16546 9064 16948 9092
rect 16942 9052 16948 9064
rect 17000 9052 17006 9104
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 18417 9095 18475 9101
rect 18417 9092 18429 9095
rect 17092 9064 18429 9092
rect 17092 9052 17098 9064
rect 18417 9061 18429 9064
rect 18463 9061 18475 9095
rect 20824 9092 20852 9132
rect 22480 9132 24952 9160
rect 22480 9092 22508 9132
rect 24946 9120 24952 9132
rect 25004 9120 25010 9172
rect 25038 9120 25044 9172
rect 25096 9160 25102 9172
rect 26237 9163 26295 9169
rect 26237 9160 26249 9163
rect 25096 9132 26249 9160
rect 25096 9120 25102 9132
rect 26237 9129 26249 9132
rect 26283 9129 26295 9163
rect 26237 9123 26295 9129
rect 20824 9064 22508 9092
rect 22557 9095 22615 9101
rect 18417 9055 18475 9061
rect 22557 9061 22569 9095
rect 22603 9092 22615 9095
rect 22603 9064 23520 9092
rect 22603 9061 22615 9064
rect 22557 9055 22615 9061
rect 8444 8996 14044 9024
rect 8444 8984 8450 8996
rect 14090 8984 14096 9036
rect 14148 9024 14154 9036
rect 15933 9027 15991 9033
rect 14148 8996 15884 9024
rect 14148 8984 14154 8996
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8925 4767 8959
rect 5350 8956 5356 8968
rect 5311 8928 5356 8956
rect 4709 8919 4767 8925
rect 5350 8916 5356 8928
rect 5408 8956 5414 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5408 8928 6009 8956
rect 5408 8916 5414 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 6822 8956 6828 8968
rect 6687 8928 6828 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8956 7803 8959
rect 15102 8956 15108 8968
rect 7791 8928 15108 8956
rect 7791 8925 7803 8928
rect 7745 8919 7803 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 15197 8959 15255 8965
rect 15197 8925 15209 8959
rect 15243 8956 15255 8959
rect 15746 8956 15752 8968
rect 15243 8928 15752 8956
rect 15243 8925 15255 8928
rect 15197 8919 15255 8925
rect 15746 8916 15752 8928
rect 15804 8916 15810 8968
rect 15856 8965 15884 8996
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16022 9024 16028 9036
rect 15979 8996 16028 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 17865 9027 17923 9033
rect 17865 9024 17877 9027
rect 17696 8996 17877 9024
rect 17696 8968 17724 8996
rect 17865 8993 17877 8996
rect 17911 8993 17923 9027
rect 17865 8987 17923 8993
rect 18966 8984 18972 9036
rect 19024 9024 19030 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19024 8996 19625 9024
rect 19024 8984 19030 8996
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 19797 9027 19855 9033
rect 19797 8993 19809 9027
rect 19843 9024 19855 9027
rect 22002 9024 22008 9036
rect 19843 8996 22008 9024
rect 19843 8993 19855 8996
rect 19797 8987 19855 8993
rect 22002 8984 22008 8996
rect 22060 8984 22066 9036
rect 23198 9024 23204 9036
rect 23159 8996 23204 9024
rect 23198 8984 23204 8996
rect 23256 8984 23262 9036
rect 23492 9033 23520 9064
rect 23477 9027 23535 9033
rect 23477 8993 23489 9027
rect 23523 9024 23535 9027
rect 23523 8996 24256 9024
rect 23523 8993 23535 8996
rect 23477 8987 23535 8993
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 16485 8959 16543 8965
rect 16485 8925 16497 8959
rect 16531 8956 16543 8959
rect 16666 8956 16672 8968
rect 16531 8928 16672 8956
rect 16531 8925 16543 8928
rect 16485 8919 16543 8925
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8956 17371 8959
rect 17494 8956 17500 8968
rect 17359 8928 17500 8956
rect 17359 8925 17371 8928
rect 17313 8919 17371 8925
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 17678 8916 17684 8968
rect 17736 8916 17742 8968
rect 20717 8959 20775 8965
rect 20717 8956 20729 8959
rect 19352 8928 20729 8956
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 5368 8888 5396 8916
rect 4028 8860 5396 8888
rect 6089 8891 6147 8897
rect 4028 8848 4034 8860
rect 6089 8857 6101 8891
rect 6135 8888 6147 8891
rect 7558 8888 7564 8900
rect 6135 8860 7564 8888
rect 6135 8857 6147 8860
rect 6089 8851 6147 8857
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 15930 8888 15936 8900
rect 8260 8860 15936 8888
rect 8260 8848 8266 8860
rect 15930 8848 15936 8860
rect 15988 8848 15994 8900
rect 16577 8891 16635 8897
rect 16577 8857 16589 8891
rect 16623 8888 16635 8891
rect 17934 8891 17992 8897
rect 17934 8888 17946 8891
rect 16623 8860 17946 8888
rect 16623 8857 16635 8860
rect 16577 8851 16635 8857
rect 17934 8857 17946 8860
rect 17980 8857 17992 8891
rect 17934 8851 17992 8857
rect 5994 8780 6000 8832
rect 6052 8820 6058 8832
rect 11514 8820 11520 8832
rect 6052 8792 11520 8820
rect 6052 8780 6058 8792
rect 11514 8780 11520 8792
rect 11572 8780 11578 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 16482 8820 16488 8832
rect 12032 8792 16488 8820
rect 12032 8780 12038 8792
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 19352 8820 19380 8928
rect 20717 8925 20729 8928
rect 20763 8925 20775 8959
rect 20717 8919 20775 8925
rect 17000 8792 19380 8820
rect 17000 8780 17006 8792
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 20254 8820 20260 8832
rect 19484 8792 20260 8820
rect 19484 8780 19490 8792
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 20732 8820 20760 8919
rect 20806 8916 20812 8968
rect 20864 8956 20870 8968
rect 20864 8928 20909 8956
rect 20864 8916 20870 8928
rect 20990 8848 20996 8900
rect 21048 8888 21054 8900
rect 22005 8891 22063 8897
rect 22005 8888 22017 8891
rect 21048 8860 22017 8888
rect 21048 8848 21054 8860
rect 22005 8857 22017 8860
rect 22051 8857 22063 8891
rect 22005 8851 22063 8857
rect 22094 8848 22100 8900
rect 22152 8888 22158 8900
rect 23293 8891 23351 8897
rect 22152 8860 22197 8888
rect 22152 8848 22158 8860
rect 23293 8857 23305 8891
rect 23339 8888 23351 8891
rect 23566 8888 23572 8900
rect 23339 8860 23572 8888
rect 23339 8857 23351 8860
rect 23293 8851 23351 8857
rect 23566 8848 23572 8860
rect 23624 8848 23630 8900
rect 24228 8888 24256 8996
rect 24762 8984 24768 9036
rect 24820 9024 24826 9036
rect 24820 8996 27568 9024
rect 24820 8984 24826 8996
rect 24946 8916 24952 8968
rect 25004 8956 25010 8968
rect 25409 8959 25467 8965
rect 25409 8956 25421 8959
rect 25004 8928 25421 8956
rect 25004 8916 25010 8928
rect 25409 8925 25421 8928
rect 25455 8925 25467 8959
rect 26142 8956 26148 8968
rect 26103 8928 26148 8956
rect 25409 8919 25467 8925
rect 26142 8916 26148 8928
rect 26200 8916 26206 8968
rect 27540 8965 27568 8996
rect 27525 8959 27583 8965
rect 27525 8925 27537 8959
rect 27571 8925 27583 8959
rect 27525 8919 27583 8925
rect 32858 8916 32864 8968
rect 32916 8956 32922 8968
rect 38013 8959 38071 8965
rect 38013 8956 38025 8959
rect 32916 8928 38025 8956
rect 32916 8916 32922 8928
rect 38013 8925 38025 8928
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 28718 8888 28724 8900
rect 24228 8860 28724 8888
rect 28718 8848 28724 8860
rect 28776 8848 28782 8900
rect 22830 8820 22836 8832
rect 20732 8792 22836 8820
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 25222 8820 25228 8832
rect 25183 8792 25228 8820
rect 25222 8780 25228 8792
rect 25280 8780 25286 8832
rect 27617 8823 27675 8829
rect 27617 8789 27629 8823
rect 27663 8820 27675 8823
rect 30282 8820 30288 8832
rect 27663 8792 30288 8820
rect 27663 8789 27675 8792
rect 27617 8783 27675 8789
rect 30282 8780 30288 8792
rect 30340 8780 30346 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 1596 8588 6561 8616
rect 1596 8489 1624 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 6549 8579 6607 8585
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 6696 8588 16957 8616
rect 6696 8576 6702 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 16945 8579 17003 8585
rect 19429 8619 19487 8625
rect 19429 8585 19441 8619
rect 19475 8616 19487 8619
rect 21910 8616 21916 8628
rect 19475 8588 21916 8616
rect 19475 8585 19487 8588
rect 19429 8579 19487 8585
rect 21910 8576 21916 8588
rect 21968 8576 21974 8628
rect 23566 8616 23572 8628
rect 23527 8588 23572 8616
rect 23566 8576 23572 8588
rect 23624 8576 23630 8628
rect 8202 8548 8208 8560
rect 5828 8520 8208 8548
rect 5828 8489 5856 8520
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 8389 8551 8447 8557
rect 8389 8517 8401 8551
rect 8435 8548 8447 8551
rect 9582 8548 9588 8560
rect 8435 8520 9588 8548
rect 8435 8517 8447 8520
rect 8389 8511 8447 8517
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 13814 8548 13820 8560
rect 13280 8520 13820 8548
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 5951 8452 6745 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 6733 8449 6745 8452
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 8294 8480 8300 8492
rect 6880 8452 8300 8480
rect 6880 8440 6886 8452
rect 8294 8440 8300 8452
rect 8352 8480 8358 8492
rect 9398 8480 9404 8492
rect 8352 8452 9404 8480
rect 8352 8440 8358 8452
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 13280 8489 13308 8520
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 17494 8548 17500 8560
rect 15028 8520 17500 8548
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 3326 8372 3332 8424
rect 3384 8412 3390 8424
rect 10134 8412 10140 8424
rect 3384 8384 10140 8412
rect 3384 8372 3390 8384
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 13538 8412 13544 8424
rect 13499 8384 13544 8412
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 13630 8372 13636 8424
rect 13688 8412 13694 8424
rect 14660 8412 14688 8466
rect 15028 8421 15056 8520
rect 17494 8508 17500 8520
rect 17552 8508 17558 8560
rect 17678 8508 17684 8560
rect 17736 8548 17742 8560
rect 18141 8551 18199 8557
rect 18141 8548 18153 8551
rect 17736 8520 18153 8548
rect 17736 8508 17742 8520
rect 18141 8517 18153 8520
rect 18187 8548 18199 8551
rect 22370 8548 22376 8560
rect 18187 8520 22376 8548
rect 18187 8517 18199 8520
rect 18141 8511 18199 8517
rect 22370 8508 22376 8520
rect 22428 8508 22434 8560
rect 22830 8508 22836 8560
rect 22888 8548 22894 8560
rect 27890 8548 27896 8560
rect 22888 8520 27896 8548
rect 22888 8508 22894 8520
rect 27890 8508 27896 8520
rect 27948 8508 27954 8560
rect 15470 8480 15476 8492
rect 15383 8452 15476 8480
rect 15470 8440 15476 8452
rect 15528 8480 15534 8492
rect 16022 8480 16028 8492
rect 15528 8452 16028 8480
rect 15528 8440 15534 8452
rect 16022 8440 16028 8452
rect 16080 8440 16086 8492
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8478 16175 8483
rect 16163 8450 16252 8478
rect 16163 8449 16175 8450
rect 16117 8443 16175 8449
rect 13688 8384 14688 8412
rect 15013 8415 15071 8421
rect 13688 8372 13694 8384
rect 15013 8381 15025 8415
rect 15059 8381 15071 8415
rect 16224 8412 16252 8450
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16816 8452 16865 8480
rect 16816 8440 16822 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 18785 8483 18843 8489
rect 18785 8480 18797 8483
rect 16853 8443 16911 8449
rect 17328 8452 18797 8480
rect 17328 8412 17356 8452
rect 18785 8449 18797 8452
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8449 19671 8483
rect 23014 8480 23020 8492
rect 22975 8452 23020 8480
rect 19613 8443 19671 8449
rect 17494 8412 17500 8424
rect 15013 8375 15071 8381
rect 15488 8384 17356 8412
rect 17455 8384 17500 8412
rect 1762 8344 1768 8356
rect 1723 8316 1768 8344
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 3142 8304 3148 8356
rect 3200 8344 3206 8356
rect 6638 8344 6644 8356
rect 3200 8316 6644 8344
rect 3200 8304 3206 8316
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 10152 8344 10180 8372
rect 15488 8344 15516 8384
rect 17494 8372 17500 8384
rect 17552 8372 17558 8424
rect 17681 8415 17739 8421
rect 17681 8381 17693 8415
rect 17727 8381 17739 8415
rect 19628 8412 19656 8443
rect 23014 8440 23020 8452
rect 23072 8440 23078 8492
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 23768 8412 23796 8443
rect 25222 8440 25228 8492
rect 25280 8480 25286 8492
rect 26421 8483 26479 8489
rect 26421 8480 26433 8483
rect 25280 8452 26433 8480
rect 25280 8440 25286 8452
rect 26421 8449 26433 8452
rect 26467 8449 26479 8483
rect 26421 8443 26479 8449
rect 25130 8412 25136 8424
rect 17681 8375 17739 8381
rect 18616 8384 19656 8412
rect 22848 8384 23796 8412
rect 25091 8384 25136 8412
rect 10152 8316 13400 8344
rect 13372 8276 13400 8316
rect 14568 8316 15516 8344
rect 15565 8347 15623 8353
rect 14568 8276 14596 8316
rect 15565 8313 15577 8347
rect 15611 8344 15623 8347
rect 15746 8344 15752 8356
rect 15611 8316 15752 8344
rect 15611 8313 15623 8316
rect 15565 8307 15623 8313
rect 15746 8304 15752 8316
rect 15804 8304 15810 8356
rect 16209 8347 16267 8353
rect 16209 8313 16221 8347
rect 16255 8344 16267 8347
rect 17696 8344 17724 8375
rect 18616 8353 18644 8384
rect 22848 8353 22876 8384
rect 25130 8372 25136 8384
rect 25188 8372 25194 8424
rect 25317 8415 25375 8421
rect 25317 8381 25329 8415
rect 25363 8412 25375 8415
rect 25363 8384 25820 8412
rect 25363 8381 25375 8384
rect 25317 8375 25375 8381
rect 16255 8316 17724 8344
rect 18601 8347 18659 8353
rect 16255 8313 16267 8316
rect 16209 8307 16267 8313
rect 18601 8313 18613 8347
rect 18647 8313 18659 8347
rect 18601 8307 18659 8313
rect 22833 8347 22891 8353
rect 22833 8313 22845 8347
rect 22879 8313 22891 8347
rect 25498 8344 25504 8356
rect 25459 8316 25504 8344
rect 22833 8307 22891 8313
rect 25498 8304 25504 8316
rect 25556 8304 25562 8356
rect 25792 8344 25820 8384
rect 26237 8347 26295 8353
rect 26237 8344 26249 8347
rect 25792 8316 26249 8344
rect 26237 8313 26249 8316
rect 26283 8313 26295 8347
rect 26237 8307 26295 8313
rect 13372 8248 14596 8276
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16390 8276 16396 8288
rect 16080 8248 16396 8276
rect 16080 8236 16086 8248
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 16482 8236 16488 8288
rect 16540 8276 16546 8288
rect 16666 8276 16672 8288
rect 16540 8248 16672 8276
rect 16540 8236 16546 8248
rect 16666 8236 16672 8248
rect 16724 8276 16730 8288
rect 17678 8276 17684 8288
rect 16724 8248 17684 8276
rect 16724 8236 16730 8248
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 5353 8075 5411 8081
rect 5353 8041 5365 8075
rect 5399 8072 5411 8075
rect 8662 8072 8668 8084
rect 5399 8044 8668 8072
rect 5399 8041 5411 8044
rect 5353 8035 5411 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 9088 8044 9689 8072
rect 9088 8032 9094 8044
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 13170 8072 13176 8084
rect 13131 8044 13176 8072
rect 9677 8035 9735 8041
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 16666 8072 16672 8084
rect 14700 8044 16672 8072
rect 14700 8032 14706 8044
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 17497 8075 17555 8081
rect 17497 8041 17509 8075
rect 17543 8072 17555 8075
rect 23937 8075 23995 8081
rect 17543 8044 18368 8072
rect 17543 8041 17555 8044
rect 17497 8035 17555 8041
rect 3786 7964 3792 8016
rect 3844 8004 3850 8016
rect 16942 8004 16948 8016
rect 3844 7976 16948 8004
rect 3844 7964 3850 7976
rect 16942 7964 16948 7976
rect 17000 7964 17006 8016
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 17770 7936 17776 7948
rect 5868 7908 10272 7936
rect 5868 7896 5874 7908
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5350 7868 5356 7880
rect 5307 7840 5356 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5350 7828 5356 7840
rect 5408 7868 5414 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 5408 7840 9597 7868
rect 5408 7828 5414 7840
rect 9585 7837 9597 7840
rect 9631 7868 9643 7871
rect 9766 7868 9772 7880
rect 9631 7840 9772 7868
rect 9631 7837 9643 7840
rect 9585 7831 9643 7837
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 10244 7877 10272 7908
rect 10888 7908 17776 7936
rect 10888 7877 10916 7908
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10873 7871 10931 7877
rect 10873 7837 10885 7871
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 12529 7871 12587 7877
rect 12529 7837 12541 7871
rect 12575 7837 12587 7871
rect 12529 7831 12587 7837
rect 10244 7800 10272 7831
rect 12544 7800 12572 7831
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 12676 7840 13093 7868
rect 12676 7828 12682 7840
rect 13081 7837 13093 7840
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7868 17003 7871
rect 17034 7868 17040 7880
rect 16991 7840 17040 7868
rect 16991 7837 17003 7840
rect 16945 7831 17003 7837
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 17678 7868 17684 7880
rect 17639 7840 17684 7868
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 18340 7877 18368 8044
rect 23937 8041 23949 8075
rect 23983 8072 23995 8075
rect 24670 8072 24676 8084
rect 23983 8044 24676 8072
rect 23983 8041 23995 8044
rect 23937 8035 23995 8041
rect 24670 8032 24676 8044
rect 24728 8032 24734 8084
rect 26694 8072 26700 8084
rect 26655 8044 26700 8072
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 25130 7936 25136 7948
rect 25091 7908 25136 7936
rect 25130 7896 25136 7908
rect 25188 7896 25194 7948
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 23842 7868 23848 7880
rect 23803 7840 23848 7868
rect 18325 7831 18383 7837
rect 23842 7828 23848 7840
rect 23900 7828 23906 7880
rect 26605 7871 26663 7877
rect 26605 7837 26617 7871
rect 26651 7868 26663 7871
rect 27890 7868 27896 7880
rect 26651 7840 27896 7868
rect 26651 7837 26663 7840
rect 26605 7831 26663 7837
rect 27890 7828 27896 7840
rect 27948 7828 27954 7880
rect 28718 7868 28724 7880
rect 28679 7840 28724 7868
rect 28718 7828 28724 7840
rect 28776 7828 28782 7880
rect 14458 7800 14464 7812
rect 10244 7772 12572 7800
rect 14419 7772 14464 7800
rect 14458 7760 14464 7772
rect 14516 7760 14522 7812
rect 14553 7803 14611 7809
rect 14553 7769 14565 7803
rect 14599 7769 14611 7803
rect 15102 7800 15108 7812
rect 15063 7772 15108 7800
rect 14553 7763 14611 7769
rect 10318 7732 10324 7744
rect 10279 7704 10324 7732
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7732 12403 7735
rect 13078 7732 13084 7744
rect 12391 7704 13084 7732
rect 12391 7701 12403 7704
rect 12345 7695 12403 7701
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 14568 7732 14596 7763
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 15565 7803 15623 7809
rect 15565 7769 15577 7803
rect 15611 7800 15623 7803
rect 16301 7803 16359 7809
rect 16301 7800 16313 7803
rect 15611 7772 16313 7800
rect 15611 7769 15623 7772
rect 15565 7763 15623 7769
rect 16301 7769 16313 7772
rect 16347 7769 16359 7803
rect 16301 7763 16359 7769
rect 16393 7803 16451 7809
rect 16393 7769 16405 7803
rect 16439 7800 16451 7803
rect 16439 7772 16574 7800
rect 16439 7769 16451 7772
rect 16393 7763 16451 7769
rect 15470 7732 15476 7744
rect 14568 7704 15476 7732
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 16546 7732 16574 7772
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 23474 7800 23480 7812
rect 16724 7772 23480 7800
rect 16724 7760 16730 7772
rect 23474 7760 23480 7772
rect 23532 7760 23538 7812
rect 18141 7735 18199 7741
rect 18141 7732 18153 7735
rect 16546 7704 18153 7732
rect 18141 7701 18153 7704
rect 18187 7701 18199 7735
rect 18141 7695 18199 7701
rect 28813 7735 28871 7741
rect 28813 7701 28825 7735
rect 28859 7732 28871 7735
rect 31662 7732 31668 7744
rect 28859 7704 31668 7732
rect 28859 7701 28871 7704
rect 28813 7695 28871 7701
rect 31662 7692 31668 7704
rect 31720 7692 31726 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 12986 7528 12992 7540
rect 12947 7500 12992 7528
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 14458 7528 14464 7540
rect 14419 7500 14464 7528
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 16942 7528 16948 7540
rect 16903 7500 16948 7528
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 19334 7528 19340 7540
rect 17052 7500 19340 7528
rect 9858 7460 9864 7472
rect 4816 7432 9864 7460
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 4816 7401 4844 7432
rect 9858 7420 9864 7432
rect 9916 7420 9922 7472
rect 10318 7420 10324 7472
rect 10376 7460 10382 7472
rect 11885 7463 11943 7469
rect 11885 7460 11897 7463
rect 10376 7432 11897 7460
rect 10376 7420 10382 7432
rect 11885 7429 11897 7432
rect 11931 7429 11943 7463
rect 17052 7460 17080 7500
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 22002 7528 22008 7540
rect 21963 7500 22008 7528
rect 22002 7488 22008 7500
rect 22060 7488 22066 7540
rect 22186 7488 22192 7540
rect 22244 7488 22250 7540
rect 11885 7423 11943 7429
rect 16546 7432 17080 7460
rect 19245 7463 19303 7469
rect 4801 7395 4859 7401
rect 4801 7392 4813 7395
rect 3476 7364 4813 7392
rect 3476 7352 3482 7364
rect 4801 7361 4813 7364
rect 4847 7361 4859 7395
rect 5994 7392 6000 7404
rect 5955 7364 6000 7392
rect 4801 7355 4859 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 12894 7392 12900 7404
rect 12676 7364 12900 7392
rect 12676 7352 12682 7364
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 13136 7364 15485 7392
rect 13136 7352 13142 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7392 15991 7395
rect 16546 7392 16574 7432
rect 19245 7429 19257 7463
rect 19291 7460 19303 7463
rect 20346 7460 20352 7472
rect 19291 7432 20352 7460
rect 19291 7429 19303 7432
rect 19245 7423 19303 7429
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 22204 7460 22232 7488
rect 22204 7432 23244 7460
rect 15979 7364 16574 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16816 7364 16865 7392
rect 16816 7352 16822 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 17034 7352 17040 7404
rect 17092 7392 17098 7404
rect 17497 7395 17555 7401
rect 17497 7392 17509 7395
rect 17092 7364 17509 7392
rect 17092 7352 17098 7364
rect 17497 7361 17509 7364
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22830 7392 22836 7404
rect 22235 7364 22692 7392
rect 22791 7364 22836 7392
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 9214 7324 9220 7336
rect 9175 7296 9220 7324
rect 9214 7284 9220 7296
rect 9272 7284 9278 7336
rect 11793 7327 11851 7333
rect 11793 7293 11805 7327
rect 11839 7324 11851 7327
rect 11974 7324 11980 7336
rect 11839 7296 11980 7324
rect 11839 7293 11851 7296
rect 11793 7287 11851 7293
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 17310 7324 17316 7336
rect 12299 7296 17316 7324
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 10778 7216 10784 7268
rect 10836 7256 10842 7268
rect 12268 7256 12296 7287
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 19153 7327 19211 7333
rect 19153 7293 19165 7327
rect 19199 7324 19211 7327
rect 20622 7324 20628 7336
rect 19199 7296 20628 7324
rect 19199 7293 19211 7296
rect 19153 7287 19211 7293
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 10836 7228 12296 7256
rect 15289 7259 15347 7265
rect 10836 7216 10842 7228
rect 15289 7225 15301 7259
rect 15335 7256 15347 7259
rect 17402 7256 17408 7268
rect 15335 7228 17408 7256
rect 15335 7225 15347 7228
rect 15289 7219 15347 7225
rect 17402 7216 17408 7228
rect 17460 7216 17466 7268
rect 19334 7216 19340 7268
rect 19392 7256 19398 7268
rect 22664 7265 22692 7364
rect 22830 7352 22836 7364
rect 22888 7352 22894 7404
rect 23216 7324 23244 7432
rect 23382 7392 23388 7404
rect 23343 7364 23388 7392
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 24213 7395 24271 7401
rect 24213 7392 24225 7395
rect 23523 7364 24225 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 24213 7361 24225 7364
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 34054 7352 34060 7404
rect 34112 7392 34118 7404
rect 38013 7395 38071 7401
rect 38013 7392 38025 7395
rect 34112 7364 38025 7392
rect 34112 7352 34118 7364
rect 38013 7361 38025 7364
rect 38059 7361 38071 7395
rect 38013 7355 38071 7361
rect 24026 7324 24032 7336
rect 23216 7296 24032 7324
rect 24026 7284 24032 7296
rect 24084 7284 24090 7336
rect 19705 7259 19763 7265
rect 19705 7256 19717 7259
rect 19392 7228 19717 7256
rect 19392 7216 19398 7228
rect 19705 7225 19717 7228
rect 19751 7225 19763 7259
rect 19705 7219 19763 7225
rect 22649 7259 22707 7265
rect 22649 7225 22661 7259
rect 22695 7225 22707 7259
rect 22649 7219 22707 7225
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 4893 7191 4951 7197
rect 4893 7188 4905 7191
rect 4672 7160 4905 7188
rect 4672 7148 4678 7160
rect 4893 7157 4905 7160
rect 4939 7157 4951 7191
rect 4893 7151 4951 7157
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 5592 7160 5825 7188
rect 5592 7148 5598 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 5813 7151 5871 7157
rect 16025 7191 16083 7197
rect 16025 7157 16037 7191
rect 16071 7188 16083 7191
rect 16298 7188 16304 7200
rect 16071 7160 16304 7188
rect 16071 7157 16083 7160
rect 16025 7151 16083 7157
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 17589 7191 17647 7197
rect 17589 7157 17601 7191
rect 17635 7188 17647 7191
rect 17862 7188 17868 7200
rect 17635 7160 17868 7188
rect 17635 7157 17647 7160
rect 17589 7151 17647 7157
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 24394 7188 24400 7200
rect 24355 7160 24400 7188
rect 24394 7148 24400 7160
rect 24452 7148 24458 7200
rect 38194 7188 38200 7200
rect 38155 7160 38200 7188
rect 38194 7148 38200 7160
rect 38252 7148 38258 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 5994 6984 6000 6996
rect 5955 6956 6000 6984
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 7834 6984 7840 6996
rect 7248 6956 7840 6984
rect 7248 6944 7254 6956
rect 7834 6944 7840 6956
rect 7892 6984 7898 6996
rect 15470 6984 15476 6996
rect 7892 6956 11100 6984
rect 15431 6956 15476 6984
rect 7892 6944 7898 6956
rect 10962 6916 10968 6928
rect 8956 6888 9352 6916
rect 8956 6848 8984 6888
rect 9214 6848 9220 6860
rect 2884 6820 8984 6848
rect 9175 6820 9220 6848
rect 2884 6789 2912 6820
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 9324 6848 9352 6888
rect 9646 6888 10968 6916
rect 9646 6848 9674 6888
rect 10962 6876 10968 6888
rect 11020 6876 11026 6928
rect 11072 6916 11100 6956
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 16942 6944 16948 6996
rect 17000 6984 17006 6996
rect 19242 6984 19248 6996
rect 17000 6956 19248 6984
rect 17000 6944 17006 6956
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 17034 6916 17040 6928
rect 11072 6888 17040 6916
rect 17034 6876 17040 6888
rect 17092 6876 17098 6928
rect 20622 6876 20628 6928
rect 20680 6876 20686 6928
rect 9858 6848 9864 6860
rect 9324 6820 9674 6848
rect 9819 6820 9864 6848
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 17494 6848 17500 6860
rect 11664 6820 17500 6848
rect 11664 6808 11670 6820
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 19518 6848 19524 6860
rect 19479 6820 19524 6848
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 20640 6848 20668 6876
rect 25133 6851 25191 6857
rect 25133 6848 25145 6851
rect 20640 6820 25145 6848
rect 25133 6817 25145 6820
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 2869 6743 2927 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 5994 6780 6000 6792
rect 5955 6752 6000 6780
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6730 6780 6736 6792
rect 6691 6752 6736 6780
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7374 6780 7380 6792
rect 7335 6752 7380 6780
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 11698 6780 11704 6792
rect 11659 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 12250 6780 12256 6792
rect 11931 6752 12256 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 15654 6780 15660 6792
rect 15615 6752 15660 6780
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 16114 6740 16120 6792
rect 16172 6740 16178 6792
rect 16298 6780 16304 6792
rect 16259 6752 16304 6780
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 18432 6752 19380 6780
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 9309 6715 9367 6721
rect 5684 6684 9260 6712
rect 5684 6672 5690 6684
rect 2682 6644 2688 6656
rect 2643 6616 2688 6644
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 4801 6647 4859 6653
rect 4801 6613 4813 6647
rect 4847 6644 4859 6647
rect 5810 6644 5816 6656
rect 4847 6616 5816 6644
rect 4847 6613 4859 6616
rect 4801 6607 4859 6613
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 6549 6647 6607 6653
rect 6549 6644 6561 6647
rect 6512 6616 6561 6644
rect 6512 6604 6518 6616
rect 6549 6613 6561 6616
rect 6595 6613 6607 6647
rect 7190 6644 7196 6656
rect 7151 6616 7196 6644
rect 6549 6607 6607 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 7926 6644 7932 6656
rect 7432 6616 7932 6644
rect 7432 6604 7438 6616
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 9232 6644 9260 6684
rect 9309 6681 9321 6715
rect 9355 6712 9367 6715
rect 13538 6712 13544 6724
rect 9355 6684 13544 6712
rect 9355 6681 9367 6684
rect 9309 6675 9367 6681
rect 13538 6672 13544 6684
rect 13596 6672 13602 6724
rect 16132 6712 16160 6740
rect 17770 6712 17776 6724
rect 16132 6684 17632 6712
rect 17731 6684 17776 6712
rect 12158 6644 12164 6656
rect 9232 6616 12164 6644
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 12345 6647 12403 6653
rect 12345 6613 12357 6647
rect 12391 6644 12403 6647
rect 14550 6644 14556 6656
rect 12391 6616 14556 6644
rect 12391 6613 12403 6616
rect 12345 6607 12403 6613
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 16117 6647 16175 6653
rect 16117 6613 16129 6647
rect 16163 6644 16175 6647
rect 16758 6644 16764 6656
rect 16163 6616 16764 6644
rect 16163 6613 16175 6616
rect 16117 6607 16175 6613
rect 16758 6604 16764 6616
rect 16816 6604 16822 6656
rect 17604 6644 17632 6684
rect 17770 6672 17776 6684
rect 17828 6672 17834 6724
rect 17862 6672 17868 6724
rect 17920 6712 17926 6724
rect 17920 6684 17965 6712
rect 17920 6672 17926 6684
rect 18046 6672 18052 6724
rect 18104 6712 18110 6724
rect 18432 6721 18460 6752
rect 18417 6715 18475 6721
rect 18417 6712 18429 6715
rect 18104 6684 18429 6712
rect 18104 6672 18110 6684
rect 18417 6681 18429 6684
rect 18463 6681 18475 6715
rect 18417 6675 18475 6681
rect 19058 6644 19064 6656
rect 17604 6616 19064 6644
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 19352 6644 19380 6752
rect 20530 6740 20536 6792
rect 20588 6780 20594 6792
rect 22189 6783 22247 6789
rect 22189 6780 22201 6783
rect 20588 6752 22201 6780
rect 20588 6740 20594 6752
rect 22189 6749 22201 6752
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6780 22891 6783
rect 23382 6780 23388 6792
rect 22879 6752 23388 6780
rect 22879 6749 22891 6752
rect 22833 6743 22891 6749
rect 19518 6672 19524 6724
rect 19576 6712 19582 6724
rect 19613 6715 19671 6721
rect 19613 6712 19625 6715
rect 19576 6684 19625 6712
rect 19576 6672 19582 6684
rect 19613 6681 19625 6684
rect 19659 6681 19671 6715
rect 19613 6675 19671 6681
rect 20165 6715 20223 6721
rect 20165 6681 20177 6715
rect 20211 6681 20223 6715
rect 22664 6712 22692 6743
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 23474 6740 23480 6792
rect 23532 6780 23538 6792
rect 23937 6783 23995 6789
rect 23937 6780 23949 6783
rect 23532 6752 23949 6780
rect 23532 6740 23538 6752
rect 23937 6749 23949 6752
rect 23983 6749 23995 6783
rect 23937 6743 23995 6749
rect 25041 6783 25099 6789
rect 25041 6749 25053 6783
rect 25087 6780 25099 6783
rect 27522 6780 27528 6792
rect 25087 6752 27528 6780
rect 25087 6749 25099 6752
rect 25041 6743 25099 6749
rect 27522 6740 27528 6752
rect 27580 6740 27586 6792
rect 29822 6712 29828 6724
rect 22664 6684 29828 6712
rect 20165 6675 20223 6681
rect 20180 6644 20208 6675
rect 29822 6672 29828 6684
rect 29880 6672 29886 6724
rect 19352 6616 20208 6644
rect 22005 6647 22063 6653
rect 22005 6613 22017 6647
rect 22051 6644 22063 6647
rect 22278 6644 22284 6656
rect 22051 6616 22284 6644
rect 22051 6613 22063 6616
rect 22005 6607 22063 6613
rect 22278 6604 22284 6616
rect 22336 6604 22342 6656
rect 23293 6647 23351 6653
rect 23293 6613 23305 6647
rect 23339 6644 23351 6647
rect 23474 6644 23480 6656
rect 23339 6616 23480 6644
rect 23339 6613 23351 6616
rect 23293 6607 23351 6613
rect 23474 6604 23480 6616
rect 23532 6604 23538 6656
rect 23750 6644 23756 6656
rect 23711 6616 23756 6644
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 6730 6440 6736 6452
rect 6691 6412 6736 6440
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 10778 6440 10784 6452
rect 6886 6412 10784 6440
rect 5534 6372 5540 6384
rect 1596 6344 5540 6372
rect 1596 6313 1624 6344
rect 5534 6332 5540 6344
rect 5592 6332 5598 6384
rect 6886 6372 6914 6412
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 13998 6440 14004 6452
rect 13959 6412 14004 6440
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 16853 6443 16911 6449
rect 16853 6440 16865 6443
rect 15712 6412 16865 6440
rect 15712 6400 15718 6412
rect 16853 6409 16865 6412
rect 16899 6409 16911 6443
rect 16853 6403 16911 6409
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 19426 6440 19432 6452
rect 17000 6412 19432 6440
rect 17000 6400 17006 6412
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 19705 6443 19763 6449
rect 19705 6409 19717 6443
rect 19751 6409 19763 6443
rect 20346 6440 20352 6452
rect 20307 6412 20352 6440
rect 19705 6403 19763 6409
rect 7742 6372 7748 6384
rect 5644 6344 6914 6372
rect 7116 6344 7748 6372
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6273 1639 6307
rect 2314 6304 2320 6316
rect 2275 6276 2320 6304
rect 1581 6267 1639 6273
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 5644 6313 5672 6344
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 7116 6304 7144 6344
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 7834 6332 7840 6384
rect 7892 6372 7898 6384
rect 8573 6375 8631 6381
rect 8573 6372 8585 6375
rect 7892 6344 8585 6372
rect 7892 6332 7898 6344
rect 8573 6341 8585 6344
rect 8619 6341 8631 6375
rect 8573 6335 8631 6341
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 9953 6375 10011 6381
rect 9953 6372 9965 6375
rect 9824 6344 9965 6372
rect 9824 6332 9830 6344
rect 9953 6341 9965 6344
rect 9999 6341 10011 6375
rect 9953 6335 10011 6341
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 15013 6375 15071 6381
rect 15013 6372 15025 6375
rect 13320 6344 15025 6372
rect 13320 6332 13326 6344
rect 15013 6341 15025 6344
rect 15059 6341 15071 6375
rect 15746 6372 15752 6384
rect 15707 6344 15752 6372
rect 15013 6335 15071 6341
rect 15746 6332 15752 6344
rect 15804 6332 15810 6384
rect 19720 6372 19748 6403
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 23382 6440 23388 6452
rect 23343 6412 23388 6440
rect 23382 6400 23388 6412
rect 23440 6400 23446 6452
rect 24026 6400 24032 6452
rect 24084 6440 24090 6452
rect 25777 6443 25835 6449
rect 25777 6440 25789 6443
rect 24084 6412 25789 6440
rect 24084 6400 24090 6412
rect 25777 6409 25789 6412
rect 25823 6409 25835 6443
rect 25777 6403 25835 6409
rect 19720 6344 20576 6372
rect 6779 6276 7144 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 5000 6236 5028 6267
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7248 6276 7573 6304
rect 7248 6264 7254 6276
rect 7561 6273 7573 6276
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6304 9735 6307
rect 10134 6304 10140 6316
rect 9723 6276 10140 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 12216 6276 12265 6304
rect 12216 6264 12222 6276
rect 12253 6273 12265 6276
rect 12299 6304 12311 6307
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12299 6276 13001 6304
rect 12299 6273 12311 6276
rect 12253 6267 12311 6273
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6304 13967 6307
rect 14918 6304 14924 6316
rect 13955 6276 14924 6304
rect 13955 6273 13967 6276
rect 13909 6267 13967 6273
rect 14918 6264 14924 6276
rect 14976 6264 14982 6316
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 16448 6276 17049 6304
rect 16448 6264 16454 6276
rect 17037 6273 17049 6276
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 17126 6264 17132 6316
rect 17184 6304 17190 6316
rect 17589 6307 17647 6313
rect 17589 6304 17601 6307
rect 17184 6276 17601 6304
rect 17184 6264 17190 6276
rect 17589 6273 17601 6276
rect 17635 6273 17647 6307
rect 17589 6267 17647 6273
rect 18601 6307 18659 6313
rect 18601 6273 18613 6307
rect 18647 6304 18659 6307
rect 18966 6304 18972 6316
rect 18647 6276 18972 6304
rect 18647 6273 18659 6276
rect 18601 6267 18659 6273
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19058 6264 19064 6316
rect 19116 6304 19122 6316
rect 20548 6313 20576 6344
rect 23474 6332 23480 6384
rect 23532 6372 23538 6384
rect 24394 6372 24400 6384
rect 23532 6344 24400 6372
rect 23532 6332 23538 6344
rect 24394 6332 24400 6344
rect 24452 6332 24458 6384
rect 19889 6307 19947 6313
rect 19889 6304 19901 6307
rect 19116 6276 19901 6304
rect 19116 6264 19122 6276
rect 19889 6273 19901 6276
rect 19935 6273 19947 6307
rect 19889 6267 19947 6273
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 23569 6307 23627 6313
rect 23569 6273 23581 6307
rect 23615 6304 23627 6307
rect 23750 6304 23756 6316
rect 23615 6276 23756 6304
rect 23615 6273 23627 6276
rect 23569 6267 23627 6273
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 25685 6307 25743 6313
rect 25685 6273 25697 6307
rect 25731 6304 25743 6307
rect 27154 6304 27160 6316
rect 25731 6276 27160 6304
rect 25731 6273 25743 6276
rect 25685 6267 25743 6273
rect 27154 6264 27160 6276
rect 27212 6264 27218 6316
rect 5000 6208 5488 6236
rect 1762 6168 1768 6180
rect 1723 6140 1768 6168
rect 1762 6128 1768 6140
rect 1820 6128 1826 6180
rect 5460 6177 5488 6208
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 5868 6208 8493 6236
rect 5868 6196 5874 6208
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 12066 6236 12072 6248
rect 9171 6208 12072 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 12066 6196 12072 6208
rect 12124 6196 12130 6248
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 13722 6236 13728 6248
rect 12492 6208 13728 6236
rect 12492 6196 12498 6208
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 15657 6239 15715 6245
rect 15657 6205 15669 6239
rect 15703 6236 15715 6239
rect 17402 6236 17408 6248
rect 15703 6208 17408 6236
rect 15703 6205 15715 6208
rect 15657 6199 15715 6205
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 17681 6239 17739 6245
rect 17681 6205 17693 6239
rect 17727 6236 17739 6239
rect 20070 6236 20076 6248
rect 17727 6208 20076 6236
rect 17727 6205 17739 6208
rect 17681 6199 17739 6205
rect 20070 6196 20076 6208
rect 20128 6196 20134 6248
rect 5445 6171 5503 6177
rect 5445 6137 5457 6171
rect 5491 6137 5503 6171
rect 5445 6131 5503 6137
rect 7190 6128 7196 6180
rect 7248 6168 7254 6180
rect 11606 6168 11612 6180
rect 7248 6140 11612 6168
rect 7248 6128 7254 6140
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 15102 6168 15108 6180
rect 11900 6140 15108 6168
rect 2406 6100 2412 6112
rect 2367 6072 2412 6100
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 7374 6100 7380 6112
rect 7335 6072 7380 6100
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 11900 6100 11928 6140
rect 15102 6128 15108 6140
rect 15160 6168 15166 6180
rect 16209 6171 16267 6177
rect 16209 6168 16221 6171
rect 15160 6140 16221 6168
rect 15160 6128 15166 6140
rect 16209 6137 16221 6140
rect 16255 6137 16267 6171
rect 16209 6131 16267 6137
rect 17770 6128 17776 6180
rect 17828 6168 17834 6180
rect 26510 6168 26516 6180
rect 17828 6140 26516 6168
rect 17828 6128 17834 6140
rect 26510 6128 26516 6140
rect 26568 6128 26574 6180
rect 12066 6100 12072 6112
rect 7800 6072 11928 6100
rect 12027 6072 12072 6100
rect 7800 6060 7806 6072
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 13081 6103 13139 6109
rect 13081 6069 13093 6103
rect 13127 6100 13139 6103
rect 14458 6100 14464 6112
rect 13127 6072 14464 6100
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 18874 6100 18880 6112
rect 18739 6072 18880 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 18874 6060 18880 6072
rect 18932 6060 18938 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 6328 5868 6377 5896
rect 6328 5856 6334 5868
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 7834 5896 7840 5908
rect 7795 5868 7840 5896
rect 6365 5859 6423 5865
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 12250 5896 12256 5908
rect 7984 5868 11836 5896
rect 12211 5868 12256 5896
rect 7984 5856 7990 5868
rect 2406 5788 2412 5840
rect 2464 5828 2470 5840
rect 7190 5828 7196 5840
rect 2464 5800 7196 5828
rect 2464 5788 2470 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 11698 5828 11704 5840
rect 7300 5800 11704 5828
rect 4893 5763 4951 5769
rect 4893 5729 4905 5763
rect 4939 5760 4951 5763
rect 7300 5760 7328 5800
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 11808 5828 11836 5868
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 12400 5868 14657 5896
rect 12400 5856 12406 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 21361 5899 21419 5905
rect 17460 5868 21312 5896
rect 17460 5856 17466 5868
rect 12434 5828 12440 5840
rect 11808 5800 12440 5828
rect 12434 5788 12440 5800
rect 12492 5788 12498 5840
rect 12897 5831 12955 5837
rect 12897 5797 12909 5831
rect 12943 5797 12955 5831
rect 13538 5828 13544 5840
rect 13499 5800 13544 5828
rect 12897 5791 12955 5797
rect 8294 5760 8300 5772
rect 4939 5732 7328 5760
rect 7392 5732 8300 5760
rect 4939 5729 4951 5732
rect 4893 5723 4951 5729
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 4614 5692 4620 5704
rect 4387 5664 4620 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5692 6331 5695
rect 7101 5695 7159 5701
rect 7101 5692 7113 5695
rect 6319 5664 7113 5692
rect 6319 5661 6331 5664
rect 6273 5655 6331 5661
rect 7101 5661 7113 5664
rect 7147 5692 7159 5695
rect 7392 5692 7420 5732
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 7147 5664 7420 5692
rect 7745 5695 7803 5701
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 8478 5692 8484 5704
rect 7791 5664 8484 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 4816 5624 4844 5655
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5692 12495 5695
rect 12912 5692 12940 5791
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 19334 5828 19340 5840
rect 14292 5800 19340 5828
rect 14182 5760 14188 5772
rect 13096 5732 14188 5760
rect 13096 5701 13124 5732
rect 14182 5720 14188 5732
rect 14240 5720 14246 5772
rect 14292 5769 14320 5800
rect 19334 5788 19340 5800
rect 19392 5788 19398 5840
rect 21284 5828 21312 5868
rect 21361 5865 21373 5899
rect 21407 5896 21419 5899
rect 26602 5896 26608 5908
rect 21407 5868 26608 5896
rect 21407 5865 21419 5868
rect 21361 5859 21419 5865
rect 26602 5856 26608 5868
rect 26660 5856 26666 5908
rect 29822 5896 29828 5908
rect 29783 5868 29828 5896
rect 29822 5856 29828 5868
rect 29880 5856 29886 5908
rect 23474 5828 23480 5840
rect 21284 5800 23480 5828
rect 23474 5788 23480 5800
rect 23532 5788 23538 5840
rect 14277 5763 14335 5769
rect 14277 5729 14289 5763
rect 14323 5729 14335 5763
rect 14458 5760 14464 5772
rect 14419 5732 14464 5760
rect 14277 5723 14335 5729
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 20990 5760 20996 5772
rect 14608 5732 20996 5760
rect 14608 5720 14614 5732
rect 20990 5720 20996 5732
rect 21048 5720 21054 5772
rect 26326 5720 26332 5772
rect 26384 5760 26390 5772
rect 37737 5763 37795 5769
rect 37737 5760 37749 5763
rect 26384 5732 37749 5760
rect 26384 5720 26390 5732
rect 37737 5729 37749 5732
rect 37783 5729 37795 5763
rect 37737 5723 37795 5729
rect 12483 5664 12940 5692
rect 13081 5695 13139 5701
rect 12483 5661 12495 5664
rect 12437 5655 12495 5661
rect 13081 5661 13093 5695
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 2832 5596 4844 5624
rect 7193 5627 7251 5633
rect 2832 5584 2838 5596
rect 7193 5593 7205 5627
rect 7239 5624 7251 5627
rect 12526 5624 12532 5636
rect 7239 5596 12532 5624
rect 7239 5593 7251 5596
rect 7193 5587 7251 5593
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 12802 5584 12808 5636
rect 12860 5624 12866 5636
rect 13740 5624 13768 5655
rect 14918 5652 14924 5704
rect 14976 5692 14982 5704
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 14976 5664 15853 5692
rect 14976 5652 14982 5664
rect 15841 5661 15853 5664
rect 15887 5692 15899 5695
rect 16485 5695 16543 5701
rect 16485 5692 16497 5695
rect 15887 5664 16497 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 16485 5661 16497 5664
rect 16531 5692 16543 5695
rect 16850 5692 16856 5704
rect 16531 5664 16856 5692
rect 16531 5661 16543 5664
rect 16485 5655 16543 5661
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 18874 5692 18880 5704
rect 18835 5664 18880 5692
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 21266 5692 21272 5704
rect 21227 5664 21272 5692
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 29733 5695 29791 5701
rect 29733 5661 29745 5695
rect 29779 5692 29791 5695
rect 36722 5692 36728 5704
rect 29779 5664 36728 5692
rect 29779 5661 29791 5664
rect 29733 5655 29791 5661
rect 36722 5652 36728 5664
rect 36780 5652 36786 5704
rect 37182 5652 37188 5704
rect 37240 5692 37246 5704
rect 37461 5695 37519 5701
rect 37461 5692 37473 5695
rect 37240 5664 37473 5692
rect 37240 5652 37246 5664
rect 37461 5661 37473 5664
rect 37507 5661 37519 5695
rect 37461 5655 37519 5661
rect 12860 5596 13768 5624
rect 12860 5584 12866 5596
rect 16574 5584 16580 5636
rect 16632 5624 16638 5636
rect 16632 5596 16677 5624
rect 16632 5584 16638 5596
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 4157 5559 4215 5565
rect 4157 5556 4169 5559
rect 2924 5528 4169 5556
rect 2924 5516 2930 5528
rect 4157 5525 4169 5528
rect 4203 5525 4215 5559
rect 4157 5519 4215 5525
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 15933 5559 15991 5565
rect 15933 5556 15945 5559
rect 11572 5528 15945 5556
rect 11572 5516 11578 5528
rect 15933 5525 15945 5528
rect 15979 5525 15991 5559
rect 15933 5519 15991 5525
rect 18693 5559 18751 5565
rect 18693 5525 18705 5559
rect 18739 5556 18751 5559
rect 20070 5556 20076 5568
rect 18739 5528 20076 5556
rect 18739 5525 18751 5528
rect 18693 5519 18751 5525
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 17862 5352 17868 5364
rect 6886 5324 17868 5352
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5216 1639 5219
rect 6454 5216 6460 5228
rect 1627 5188 6460 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 6454 5176 6460 5188
rect 6512 5176 6518 5228
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6886 5216 6914 5324
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 7374 5284 7380 5296
rect 7335 5256 7380 5284
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 10413 5287 10471 5293
rect 10413 5253 10425 5287
rect 10459 5284 10471 5287
rect 12894 5284 12900 5296
rect 10459 5256 12900 5284
rect 10459 5253 10471 5256
rect 10413 5247 10471 5253
rect 12894 5244 12900 5256
rect 12952 5244 12958 5296
rect 30282 5244 30288 5296
rect 30340 5284 30346 5296
rect 30340 5256 32536 5284
rect 30340 5244 30346 5256
rect 10134 5216 10140 5228
rect 6595 5188 6914 5216
rect 10095 5188 10140 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 12342 5216 12348 5228
rect 11747 5188 12348 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 18414 5216 18420 5228
rect 15335 5188 18420 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 7282 5148 7288 5160
rect 7243 5120 7288 5148
rect 7282 5108 7288 5120
rect 7340 5108 7346 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 11974 5148 11980 5160
rect 7975 5120 11980 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 14016 5148 14044 5179
rect 18414 5176 18420 5188
rect 18472 5176 18478 5228
rect 31662 5216 31668 5228
rect 31623 5188 31668 5216
rect 31662 5176 31668 5188
rect 31720 5176 31726 5228
rect 32508 5225 32536 5256
rect 32493 5219 32551 5225
rect 32493 5185 32505 5219
rect 32539 5185 32551 5219
rect 32493 5179 32551 5185
rect 15381 5151 15439 5157
rect 15381 5148 15393 5151
rect 14016 5120 15393 5148
rect 15381 5117 15393 5120
rect 15427 5117 15439 5151
rect 15381 5111 15439 5117
rect 31481 5083 31539 5089
rect 31481 5049 31493 5083
rect 31527 5080 31539 5083
rect 33686 5080 33692 5092
rect 31527 5052 33692 5080
rect 31527 5049 31539 5052
rect 31481 5043 31539 5049
rect 33686 5040 33692 5052
rect 33744 5040 33750 5092
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 6638 5012 6644 5024
rect 6599 4984 6644 5012
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 11790 5012 11796 5024
rect 11751 4984 11796 5012
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 13817 5015 13875 5021
rect 13817 4981 13829 5015
rect 13863 5012 13875 5015
rect 14274 5012 14280 5024
rect 13863 4984 14280 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 32309 5015 32367 5021
rect 32309 4981 32321 5015
rect 32355 5012 32367 5015
rect 34054 5012 34060 5024
rect 32355 4984 34060 5012
rect 32355 4981 32367 4984
rect 32309 4975 32367 4981
rect 34054 4972 34060 4984
rect 34112 4972 34118 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 12066 4604 12072 4616
rect 12027 4576 12072 4604
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 17681 4607 17739 4613
rect 17681 4604 17693 4607
rect 13780 4576 17693 4604
rect 13780 4564 13786 4576
rect 17681 4573 17693 4576
rect 17727 4573 17739 4607
rect 17681 4567 17739 4573
rect 27709 4607 27767 4613
rect 27709 4573 27721 4607
rect 27755 4604 27767 4607
rect 35618 4604 35624 4616
rect 27755 4576 35624 4604
rect 27755 4573 27767 4576
rect 27709 4567 27767 4573
rect 35618 4564 35624 4576
rect 35676 4564 35682 4616
rect 11146 4468 11152 4480
rect 11107 4440 11152 4468
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 11882 4468 11888 4480
rect 11843 4440 11888 4468
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 17773 4471 17831 4477
rect 17773 4437 17785 4471
rect 17819 4468 17831 4471
rect 18322 4468 18328 4480
rect 17819 4440 18328 4468
rect 17819 4437 17831 4440
rect 17773 4431 17831 4437
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 27798 4468 27804 4480
rect 27759 4440 27804 4468
rect 27798 4428 27804 4440
rect 27856 4428 27862 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 12342 4264 12348 4276
rect 12303 4236 12348 4264
rect 12342 4224 12348 4236
rect 12400 4224 12406 4276
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11204 4100 11713 4128
rect 11204 4088 11210 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11882 4128 11888 4140
rect 11843 4100 11888 4128
rect 11701 4091 11759 4097
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 16850 4088 16856 4140
rect 16908 4128 16914 4140
rect 17037 4131 17095 4137
rect 17037 4128 17049 4131
rect 16908 4100 17049 4128
rect 16908 4088 16914 4100
rect 17037 4097 17049 4100
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 16853 3995 16911 4001
rect 16853 3961 16865 3995
rect 16899 3992 16911 3995
rect 16942 3992 16948 4004
rect 16899 3964 16948 3992
rect 16899 3961 16911 3964
rect 16853 3955 16911 3961
rect 16942 3952 16948 3964
rect 17000 3952 17006 4004
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 2774 3720 2780 3732
rect 1627 3692 2780 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 1762 3516 1768 3528
rect 1723 3488 1768 3516
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 6638 3516 6644 3528
rect 6599 3488 6644 3516
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3516 11207 3519
rect 11195 3488 16574 3516
rect 11195 3485 11207 3488
rect 11149 3479 11207 3485
rect 16546 3448 16574 3488
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 17644 3488 18613 3516
rect 17644 3476 17650 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 38010 3516 38016 3528
rect 37971 3488 38016 3516
rect 18601 3479 18659 3485
rect 38010 3476 38016 3488
rect 38068 3476 38074 3528
rect 21174 3448 21180 3460
rect 16546 3420 21180 3448
rect 21174 3408 21180 3420
rect 21232 3408 21238 3460
rect 6457 3383 6515 3389
rect 6457 3349 6469 3383
rect 6503 3380 6515 3383
rect 6546 3380 6552 3392
rect 6503 3352 6552 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 11054 3340 11060 3392
rect 11112 3380 11118 3392
rect 11241 3383 11299 3389
rect 11241 3380 11253 3383
rect 11112 3352 11253 3380
rect 11112 3340 11118 3352
rect 11241 3349 11253 3352
rect 11287 3349 11299 3383
rect 11241 3343 11299 3349
rect 18417 3383 18475 3389
rect 18417 3349 18429 3383
rect 18463 3380 18475 3383
rect 18598 3380 18604 3392
rect 18463 3352 18604 3380
rect 18463 3349 18475 3352
rect 18417 3343 18475 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 7282 3176 7288 3188
rect 6687 3148 7288 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 13357 3179 13415 3185
rect 13357 3145 13369 3179
rect 13403 3176 13415 3179
rect 16666 3176 16672 3188
rect 13403 3148 16672 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 16850 3176 16856 3188
rect 16811 3148 16856 3176
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17586 3176 17592 3188
rect 17547 3148 17592 3176
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 36722 3176 36728 3188
rect 36683 3148 36728 3176
rect 36722 3136 36728 3148
rect 36780 3136 36786 3188
rect 2866 3108 2872 3120
rect 1596 3080 2872 3108
rect 1596 3049 1624 3080
rect 2866 3068 2872 3080
rect 2924 3068 2930 3120
rect 11790 3108 11796 3120
rect 9692 3080 11796 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2774 3040 2780 3052
rect 2547 3012 2780 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 9692 3049 9720 3080
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 18322 3108 18328 3120
rect 18283 3080 18328 3108
rect 18322 3068 18328 3080
rect 18380 3068 18386 3120
rect 34054 3068 34060 3120
rect 34112 3108 34118 3120
rect 34112 3080 38056 3108
rect 34112 3068 34118 3080
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3009 9735 3043
rect 11054 3040 11060 3052
rect 11015 3012 11060 3040
rect 9677 3003 9735 3009
rect 6564 2972 6592 3003
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 13265 3043 13323 3049
rect 13265 3040 13277 3043
rect 11204 3012 13277 3040
rect 11204 3000 11210 3012
rect 13265 3009 13277 3012
rect 13311 3009 13323 3043
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 13265 3003 13323 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 17218 3000 17224 3052
rect 17276 3040 17282 3052
rect 17497 3043 17555 3049
rect 17497 3040 17509 3043
rect 17276 3012 17509 3040
rect 17276 3000 17282 3012
rect 17497 3009 17509 3012
rect 17543 3009 17555 3043
rect 36906 3040 36912 3052
rect 36867 3012 36912 3040
rect 17497 3003 17555 3009
rect 36906 3000 36912 3012
rect 36964 3000 36970 3052
rect 38028 3049 38056 3080
rect 38013 3043 38071 3049
rect 38013 3009 38025 3043
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 2332 2944 6592 2972
rect 18233 2975 18291 2981
rect 2332 2913 2360 2944
rect 18233 2941 18245 2975
rect 18279 2972 18291 2975
rect 27798 2972 27804 2984
rect 18279 2944 27804 2972
rect 18279 2941 18291 2944
rect 18233 2935 18291 2941
rect 27798 2932 27804 2944
rect 27856 2932 27862 2984
rect 2317 2907 2375 2913
rect 2317 2873 2329 2907
rect 2363 2873 2375 2907
rect 2317 2867 2375 2873
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 10873 2907 10931 2913
rect 10873 2904 10885 2907
rect 8352 2876 10885 2904
rect 8352 2864 8358 2876
rect 10873 2873 10885 2876
rect 10919 2873 10931 2907
rect 10873 2867 10931 2873
rect 11974 2864 11980 2916
rect 12032 2904 12038 2916
rect 18785 2907 18843 2913
rect 18785 2904 18797 2907
rect 12032 2876 18797 2904
rect 12032 2864 12038 2876
rect 18785 2873 18797 2876
rect 18831 2873 18843 2907
rect 18785 2867 18843 2873
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 72 2808 1777 2836
rect 72 2796 78 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 9493 2839 9551 2845
rect 9493 2836 9505 2839
rect 9180 2808 9505 2836
rect 9180 2796 9186 2808
rect 9493 2805 9505 2808
rect 9539 2805 9551 2839
rect 38194 2836 38200 2848
rect 38155 2808 38200 2836
rect 9493 2799 9551 2805
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2685 2635 2743 2641
rect 2685 2601 2697 2635
rect 2731 2632 2743 2635
rect 4706 2632 4712 2644
rect 2731 2604 4712 2632
rect 2731 2601 2743 2604
rect 2685 2595 2743 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 11146 2632 11152 2644
rect 10459 2604 11152 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 15565 2635 15623 2641
rect 15565 2601 15577 2635
rect 15611 2632 15623 2635
rect 17126 2632 17132 2644
rect 15611 2604 17132 2632
rect 15611 2601 15623 2604
rect 15565 2595 15623 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 21266 2592 21272 2644
rect 21324 2632 21330 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 21324 2604 22017 2632
rect 21324 2592 21330 2604
rect 22005 2601 22017 2604
rect 22051 2601 22063 2635
rect 22005 2595 22063 2601
rect 23842 2592 23848 2644
rect 23900 2632 23906 2644
rect 24581 2635 24639 2641
rect 24581 2632 24593 2635
rect 23900 2604 24593 2632
rect 23900 2592 23906 2604
rect 24581 2601 24593 2604
rect 24627 2601 24639 2635
rect 27154 2632 27160 2644
rect 27115 2604 27160 2632
rect 24581 2595 24639 2601
rect 27154 2592 27160 2604
rect 27212 2592 27218 2644
rect 27522 2592 27528 2644
rect 27580 2632 27586 2644
rect 27801 2635 27859 2641
rect 27801 2632 27813 2635
rect 27580 2604 27813 2632
rect 27580 2592 27586 2604
rect 27801 2601 27813 2604
rect 27847 2601 27859 2635
rect 29730 2632 29736 2644
rect 29691 2604 29736 2632
rect 27801 2595 27859 2601
rect 29730 2592 29736 2604
rect 29788 2592 29794 2644
rect 32306 2632 32312 2644
rect 32267 2604 32312 2632
rect 32306 2592 32312 2604
rect 32364 2592 32370 2644
rect 33042 2592 33048 2644
rect 33100 2632 33106 2644
rect 35529 2635 35587 2641
rect 35529 2632 35541 2635
rect 33100 2604 35541 2632
rect 33100 2592 33106 2604
rect 35529 2601 35541 2604
rect 35575 2601 35587 2635
rect 35529 2595 35587 2601
rect 35618 2592 35624 2644
rect 35676 2632 35682 2644
rect 36725 2635 36783 2641
rect 36725 2632 36737 2635
rect 35676 2604 36737 2632
rect 35676 2592 35682 2604
rect 36725 2601 36737 2604
rect 36771 2601 36783 2635
rect 36725 2595 36783 2601
rect 4798 2564 4804 2576
rect 1596 2536 4804 2564
rect 1596 2437 1624 2536
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 10134 2524 10140 2576
rect 10192 2564 10198 2576
rect 12345 2567 12403 2573
rect 12345 2564 12357 2567
rect 10192 2536 12357 2564
rect 10192 2524 10198 2536
rect 12345 2533 12357 2536
rect 12391 2533 12403 2567
rect 12345 2527 12403 2533
rect 27890 2524 27896 2576
rect 27948 2564 27954 2576
rect 31021 2567 31079 2573
rect 31021 2564 31033 2567
rect 27948 2536 31033 2564
rect 27948 2524 27954 2536
rect 31021 2533 31033 2536
rect 31067 2533 31079 2567
rect 31021 2527 31079 2533
rect 7098 2496 7104 2508
rect 4632 2468 7104 2496
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 4632 2437 4660 2468
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 33686 2456 33692 2508
rect 33744 2496 33750 2508
rect 33744 2468 37504 2496
rect 33744 2456 33750 2468
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2648 2400 2881 2428
rect 2648 2388 2654 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 4617 2391 4675 2397
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8294 2428 8300 2440
rect 7883 2400 8300 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12308 2400 12541 2428
rect 12308 2388 12314 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 14274 2428 14280 2440
rect 14235 2400 14280 2428
rect 12529 2391 12587 2397
rect 14274 2388 14280 2400
rect 14332 2388 14338 2440
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15528 2400 15761 2428
rect 15528 2388 15534 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 18598 2428 18604 2440
rect 18559 2400 18604 2428
rect 16853 2391 16911 2397
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21324 2400 22201 2428
rect 21324 2388 21330 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 23293 2431 23351 2437
rect 23293 2428 23305 2431
rect 22336 2400 23305 2428
rect 22336 2388 22342 2400
rect 23293 2397 23305 2400
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24544 2400 24777 2428
rect 24544 2388 24550 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 26476 2400 27353 2428
rect 26476 2388 26482 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 27985 2431 28043 2437
rect 27985 2428 27997 2431
rect 27764 2400 27997 2428
rect 27764 2388 27770 2400
rect 27985 2397 27997 2400
rect 28031 2397 28043 2431
rect 27985 2391 28043 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 30926 2388 30932 2440
rect 30984 2428 30990 2440
rect 31205 2431 31263 2437
rect 31205 2428 31217 2431
rect 30984 2400 31217 2428
rect 30984 2388 30990 2400
rect 31205 2397 31217 2400
rect 31251 2397 31263 2431
rect 31205 2391 31263 2397
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 32272 2400 32505 2428
rect 32272 2388 32278 2400
rect 32493 2397 32505 2400
rect 32539 2397 32551 2431
rect 32493 2391 32551 2397
rect 34146 2388 34152 2440
rect 34204 2428 34210 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34204 2400 35081 2428
rect 34204 2388 34210 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35069 2391 35127 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 37476 2437 37504 2468
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 36909 2431 36967 2437
rect 36909 2397 36921 2431
rect 36955 2397 36967 2431
rect 36909 2391 36967 2397
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 26142 2320 26148 2372
rect 26200 2360 26206 2372
rect 36924 2360 36952 2391
rect 38654 2360 38660 2372
rect 26200 2332 34928 2360
rect 36924 2332 38660 2360
rect 26200 2320 26206 2332
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1765 2295 1823 2301
rect 1765 2292 1777 2295
rect 1360 2264 1777 2292
rect 1360 2252 1366 2264
rect 1765 2261 1777 2264
rect 1811 2261 1823 2295
rect 1765 2255 1823 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4580 2264 4813 2292
rect 4580 2252 4586 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 5868 2264 6745 2292
rect 5868 2252 5874 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 14461 2295 14519 2301
rect 14461 2292 14473 2295
rect 13596 2264 14473 2292
rect 13596 2252 13602 2264
rect 14461 2261 14473 2264
rect 14507 2261 14519 2295
rect 14461 2255 14519 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18748 2264 18797 2292
rect 18748 2252 18754 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 18785 2255 18843 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 20036 2264 20269 2292
rect 20036 2252 20042 2264
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 34900 2301 34928 2332
rect 38654 2320 38660 2332
rect 38712 2320 38718 2372
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23256 2264 23489 2292
rect 23256 2252 23262 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 34885 2295 34943 2301
rect 34885 2261 34897 2295
rect 34931 2261 34943 2295
rect 34885 2255 34943 2261
rect 37366 2252 37372 2304
rect 37424 2292 37430 2304
rect 37645 2295 37703 2301
rect 37645 2292 37657 2295
rect 37424 2264 37657 2292
rect 37424 2252 37430 2264
rect 37645 2261 37657 2264
rect 37691 2261 37703 2295
rect 37645 2255 37703 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 39304 37408 39356 37460
rect 37464 37315 37516 37324
rect 37464 37281 37473 37315
rect 37473 37281 37507 37315
rect 37507 37281 37516 37315
rect 37464 37272 37516 37281
rect 1584 37247 1636 37256
rect 1584 37213 1593 37247
rect 1593 37213 1627 37247
rect 1627 37213 1636 37247
rect 1584 37204 1636 37213
rect 1952 37204 2004 37256
rect 3148 37247 3200 37256
rect 3148 37213 3157 37247
rect 3157 37213 3191 37247
rect 3191 37213 3200 37247
rect 3148 37204 3200 37213
rect 4160 37247 4212 37256
rect 4160 37213 4169 37247
rect 4169 37213 4203 37247
rect 4203 37213 4212 37247
rect 4160 37204 4212 37213
rect 5172 37204 5224 37256
rect 7104 37204 7156 37256
rect 8392 37204 8444 37256
rect 10324 37204 10376 37256
rect 11612 37204 11664 37256
rect 11980 37204 12032 37256
rect 14832 37204 14884 37256
rect 16120 37204 16172 37256
rect 17224 37204 17276 37256
rect 18972 37204 19024 37256
rect 20812 37204 20864 37256
rect 22560 37204 22612 37256
rect 23296 37204 23348 37256
rect 25780 37204 25832 37256
rect 27160 37247 27212 37256
rect 27160 37213 27169 37247
rect 27169 37213 27203 37247
rect 27203 37213 27212 37247
rect 27160 37204 27212 37213
rect 29000 37204 29052 37256
rect 30380 37204 30432 37256
rect 31760 37204 31812 37256
rect 33508 37204 33560 37256
rect 34796 37204 34848 37256
rect 35440 37204 35492 37256
rect 36636 37247 36688 37256
rect 36636 37213 36645 37247
rect 36645 37213 36679 37247
rect 36679 37213 36688 37247
rect 36636 37204 36688 37213
rect 37740 37247 37792 37256
rect 37740 37213 37749 37247
rect 37749 37213 37783 37247
rect 37783 37213 37792 37247
rect 37740 37204 37792 37213
rect 2780 37136 2832 37188
rect 2320 37111 2372 37120
rect 2320 37077 2329 37111
rect 2329 37077 2363 37111
rect 2363 37077 2372 37111
rect 2320 37068 2372 37077
rect 3884 37068 3936 37120
rect 6828 37136 6880 37188
rect 23756 37136 23808 37188
rect 4620 37068 4672 37120
rect 7196 37111 7248 37120
rect 7196 37077 7205 37111
rect 7205 37077 7239 37111
rect 7239 37077 7248 37111
rect 7196 37068 7248 37077
rect 9128 37111 9180 37120
rect 9128 37077 9137 37111
rect 9137 37077 9171 37111
rect 9171 37077 9180 37111
rect 9128 37068 9180 37077
rect 10416 37111 10468 37120
rect 10416 37077 10425 37111
rect 10425 37077 10459 37111
rect 10459 37077 10468 37111
rect 10416 37068 10468 37077
rect 11704 37111 11756 37120
rect 11704 37077 11713 37111
rect 11713 37077 11747 37111
rect 11747 37077 11756 37111
rect 11704 37068 11756 37077
rect 12900 37068 12952 37120
rect 14740 37068 14792 37120
rect 16580 37068 16632 37120
rect 18052 37068 18104 37120
rect 19340 37068 19392 37120
rect 20720 37068 20772 37120
rect 20996 37068 21048 37120
rect 23848 37068 23900 37120
rect 27436 37136 27488 37188
rect 27068 37068 27120 37120
rect 29736 37111 29788 37120
rect 29736 37077 29745 37111
rect 29745 37077 29779 37111
rect 29779 37077 29788 37111
rect 29736 37068 29788 37077
rect 30380 37111 30432 37120
rect 30380 37077 30389 37111
rect 30389 37077 30423 37111
rect 30423 37077 30432 37111
rect 30380 37068 30432 37077
rect 32404 37068 32456 37120
rect 34612 37068 34664 37120
rect 36728 37068 36780 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 664 36864 716 36916
rect 2872 36728 2924 36780
rect 34336 36771 34388 36780
rect 34336 36737 34345 36771
rect 34345 36737 34379 36771
rect 34379 36737 34388 36771
rect 34336 36728 34388 36737
rect 38016 36864 38068 36916
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 36636 36320 36688 36372
rect 38200 36363 38252 36372
rect 38200 36329 38209 36363
rect 38209 36329 38243 36363
rect 38243 36329 38252 36363
rect 38200 36320 38252 36329
rect 1768 36159 1820 36168
rect 1768 36125 1777 36159
rect 1777 36125 1811 36159
rect 1811 36125 1820 36159
rect 1768 36116 1820 36125
rect 29828 36116 29880 36168
rect 38016 36159 38068 36168
rect 38016 36125 38025 36159
rect 38025 36125 38059 36159
rect 38059 36125 38068 36159
rect 38016 36116 38068 36125
rect 3516 35980 3568 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 34336 35776 34388 35828
rect 33324 35683 33376 35692
rect 33324 35649 33333 35683
rect 33333 35649 33367 35683
rect 33367 35649 33376 35683
rect 33324 35640 33376 35649
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 38292 35071 38344 35080
rect 38292 35037 38301 35071
rect 38301 35037 38335 35071
rect 38335 35037 38344 35071
rect 38292 35028 38344 35037
rect 37280 34892 37332 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1584 34688 1636 34740
rect 38016 34688 38068 34740
rect 1952 34595 2004 34604
rect 1952 34561 1961 34595
rect 1961 34561 1995 34595
rect 1995 34561 2004 34595
rect 1952 34552 2004 34561
rect 15292 34595 15344 34604
rect 15292 34561 15301 34595
rect 15301 34561 15335 34595
rect 15335 34561 15344 34595
rect 15292 34552 15344 34561
rect 36452 34552 36504 34604
rect 17408 34484 17460 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 35440 34144 35492 34196
rect 12164 34008 12216 34060
rect 1768 33983 1820 33992
rect 1768 33949 1777 33983
rect 1777 33949 1811 33983
rect 1811 33949 1820 33983
rect 1768 33940 1820 33949
rect 1676 33804 1728 33856
rect 12624 33847 12676 33856
rect 12624 33813 12633 33847
rect 12633 33813 12667 33847
rect 12667 33813 12676 33847
rect 12624 33804 12676 33813
rect 34520 33940 34572 33992
rect 13544 33804 13596 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1952 33643 2004 33652
rect 1952 33609 1961 33643
rect 1961 33609 1995 33643
rect 1995 33609 2004 33643
rect 1952 33600 2004 33609
rect 17224 33643 17276 33652
rect 17224 33609 17233 33643
rect 17233 33609 17267 33643
rect 17267 33609 17276 33643
rect 17224 33600 17276 33609
rect 23296 33643 23348 33652
rect 23296 33609 23305 33643
rect 23305 33609 23339 33643
rect 23339 33609 23348 33643
rect 23296 33600 23348 33609
rect 12624 33532 12676 33584
rect 2136 33464 2188 33516
rect 12164 33464 12216 33516
rect 13544 33507 13596 33516
rect 13544 33473 13553 33507
rect 13553 33473 13587 33507
rect 13587 33473 13596 33507
rect 13544 33464 13596 33473
rect 17408 33507 17460 33516
rect 17408 33473 17417 33507
rect 17417 33473 17451 33507
rect 17451 33473 17460 33507
rect 17408 33464 17460 33473
rect 22836 33464 22888 33516
rect 38292 33507 38344 33516
rect 38292 33473 38301 33507
rect 38301 33473 38335 33507
rect 38335 33473 38344 33507
rect 38292 33464 38344 33473
rect 3056 33396 3108 33448
rect 2228 33260 2280 33312
rect 11796 33303 11848 33312
rect 11796 33269 11805 33303
rect 11805 33269 11839 33303
rect 11839 33269 11848 33303
rect 11796 33260 11848 33269
rect 13912 33303 13964 33312
rect 13912 33269 13921 33303
rect 13921 33269 13955 33303
rect 13955 33269 13964 33303
rect 13912 33260 13964 33269
rect 15292 33260 15344 33312
rect 29460 33260 29512 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2872 33099 2924 33108
rect 2872 33065 2881 33099
rect 2881 33065 2915 33099
rect 2915 33065 2924 33099
rect 2872 33056 2924 33065
rect 27160 33056 27212 33108
rect 1768 32895 1820 32904
rect 1768 32861 1777 32895
rect 1777 32861 1811 32895
rect 1811 32861 1820 32895
rect 1768 32852 1820 32861
rect 6184 32852 6236 32904
rect 9128 32895 9180 32904
rect 9128 32861 9137 32895
rect 9137 32861 9171 32895
rect 9171 32861 9180 32895
rect 9128 32852 9180 32861
rect 13360 32852 13412 32904
rect 23296 32895 23348 32904
rect 23296 32861 23305 32895
rect 23305 32861 23339 32895
rect 23339 32861 23348 32895
rect 23296 32852 23348 32861
rect 1860 32716 1912 32768
rect 6552 32716 6604 32768
rect 11244 32716 11296 32768
rect 15384 32759 15436 32768
rect 15384 32725 15393 32759
rect 15393 32725 15427 32759
rect 15427 32725 15436 32759
rect 15384 32716 15436 32725
rect 15660 32716 15712 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 13912 32512 13964 32564
rect 18972 32555 19024 32564
rect 18972 32521 18981 32555
rect 18981 32521 19015 32555
rect 19015 32521 19024 32555
rect 18972 32512 19024 32521
rect 23296 32512 23348 32564
rect 1492 32376 1544 32428
rect 4620 32419 4672 32428
rect 4620 32385 4629 32419
rect 4629 32385 4663 32419
rect 4663 32385 4672 32419
rect 4620 32376 4672 32385
rect 6552 32419 6604 32428
rect 6552 32385 6561 32419
rect 6561 32385 6595 32419
rect 6595 32385 6604 32419
rect 6552 32376 6604 32385
rect 6828 32376 6880 32428
rect 5448 32351 5500 32360
rect 5448 32317 5457 32351
rect 5457 32317 5491 32351
rect 5491 32317 5500 32351
rect 5448 32308 5500 32317
rect 6736 32351 6788 32360
rect 6736 32317 6745 32351
rect 6745 32317 6779 32351
rect 6779 32317 6788 32351
rect 6736 32308 6788 32317
rect 11152 32376 11204 32428
rect 15384 32444 15436 32496
rect 11796 32376 11848 32428
rect 13452 32376 13504 32428
rect 14188 32419 14240 32428
rect 14188 32385 14197 32419
rect 14197 32385 14231 32419
rect 14231 32385 14240 32419
rect 14188 32376 14240 32385
rect 14740 32419 14792 32428
rect 14740 32385 14749 32419
rect 14749 32385 14783 32419
rect 14783 32385 14792 32419
rect 14740 32376 14792 32385
rect 15660 32419 15712 32428
rect 15660 32385 15669 32419
rect 15669 32385 15703 32419
rect 15703 32385 15712 32419
rect 15660 32376 15712 32385
rect 16396 32376 16448 32428
rect 19432 32376 19484 32428
rect 19340 32308 19392 32360
rect 34612 32376 34664 32428
rect 1952 32215 2004 32224
rect 1952 32181 1961 32215
rect 1961 32181 1995 32215
rect 1995 32181 2004 32215
rect 1952 32172 2004 32181
rect 7748 32215 7800 32224
rect 7748 32181 7757 32215
rect 7757 32181 7791 32215
rect 7791 32181 7800 32215
rect 7748 32172 7800 32181
rect 10140 32215 10192 32224
rect 10140 32181 10149 32215
rect 10149 32181 10183 32215
rect 10183 32181 10192 32215
rect 10140 32172 10192 32181
rect 11888 32172 11940 32224
rect 14004 32215 14056 32224
rect 14004 32181 14013 32215
rect 14013 32181 14047 32215
rect 14047 32181 14056 32215
rect 14004 32172 14056 32181
rect 14096 32172 14148 32224
rect 16028 32215 16080 32224
rect 16028 32181 16037 32215
rect 16037 32181 16071 32215
rect 16071 32181 16080 32215
rect 16028 32172 16080 32181
rect 17408 32172 17460 32224
rect 25044 32172 25096 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 5448 31968 5500 32020
rect 11980 31968 12032 32020
rect 16028 31968 16080 32020
rect 16948 31968 17000 32020
rect 2872 31900 2924 31952
rect 7380 31900 7432 31952
rect 7748 31900 7800 31952
rect 2780 31764 2832 31816
rect 9220 31832 9272 31884
rect 13636 31900 13688 31952
rect 15752 31900 15804 31952
rect 17592 31900 17644 31952
rect 21364 31875 21416 31884
rect 21364 31841 21373 31875
rect 21373 31841 21407 31875
rect 21407 31841 21416 31875
rect 21364 31832 21416 31841
rect 5264 31807 5316 31816
rect 5264 31773 5273 31807
rect 5273 31773 5307 31807
rect 5307 31773 5316 31807
rect 5264 31764 5316 31773
rect 10416 31764 10468 31816
rect 10876 31764 10928 31816
rect 12992 31807 13044 31816
rect 10600 31696 10652 31748
rect 12992 31773 13001 31807
rect 13001 31773 13035 31807
rect 13035 31773 13044 31807
rect 12992 31764 13044 31773
rect 14004 31764 14056 31816
rect 16396 31807 16448 31816
rect 16396 31773 16405 31807
rect 16405 31773 16439 31807
rect 16439 31773 16448 31807
rect 16396 31764 16448 31773
rect 16764 31764 16816 31816
rect 17408 31807 17460 31816
rect 17408 31773 17417 31807
rect 17417 31773 17451 31807
rect 17451 31773 17460 31807
rect 17408 31764 17460 31773
rect 20720 31807 20772 31816
rect 20720 31773 20729 31807
rect 20729 31773 20763 31807
rect 20763 31773 20772 31807
rect 20720 31764 20772 31773
rect 22928 31764 22980 31816
rect 29828 31832 29880 31884
rect 37372 31832 37424 31884
rect 38108 31807 38160 31816
rect 38108 31773 38117 31807
rect 38117 31773 38151 31807
rect 38151 31773 38160 31807
rect 38108 31764 38160 31773
rect 3700 31628 3752 31680
rect 11152 31628 11204 31680
rect 17224 31671 17276 31680
rect 17224 31637 17233 31671
rect 17233 31637 17267 31671
rect 17267 31637 17276 31671
rect 17224 31628 17276 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 5264 31424 5316 31476
rect 6736 31424 6788 31476
rect 10140 31356 10192 31408
rect 1952 31288 2004 31340
rect 5172 31331 5224 31340
rect 5172 31297 5181 31331
rect 5181 31297 5215 31331
rect 5215 31297 5224 31331
rect 5172 31288 5224 31297
rect 7196 31288 7248 31340
rect 10692 31331 10744 31340
rect 10692 31297 10701 31331
rect 10701 31297 10735 31331
rect 10735 31297 10744 31331
rect 10692 31288 10744 31297
rect 13452 31424 13504 31476
rect 16396 31424 16448 31476
rect 19432 31424 19484 31476
rect 20720 31467 20772 31476
rect 20720 31433 20729 31467
rect 20729 31433 20763 31467
rect 20763 31433 20772 31467
rect 20720 31424 20772 31433
rect 22928 31467 22980 31476
rect 13636 31331 13688 31340
rect 13636 31297 13645 31331
rect 13645 31297 13679 31331
rect 13679 31297 13688 31331
rect 13636 31288 13688 31297
rect 16580 31356 16632 31408
rect 16948 31399 17000 31408
rect 16948 31365 16957 31399
rect 16957 31365 16991 31399
rect 16991 31365 17000 31399
rect 16948 31356 17000 31365
rect 17224 31356 17276 31408
rect 22928 31433 22937 31467
rect 22937 31433 22971 31467
rect 22971 31433 22980 31467
rect 22928 31424 22980 31433
rect 16396 31288 16448 31340
rect 21364 31288 21416 31340
rect 22468 31331 22520 31340
rect 22468 31297 22477 31331
rect 22477 31297 22511 31331
rect 22511 31297 22520 31331
rect 22468 31288 22520 31297
rect 7380 31263 7432 31272
rect 7380 31229 7389 31263
rect 7389 31229 7423 31263
rect 7423 31229 7432 31263
rect 7380 31220 7432 31229
rect 7748 31220 7800 31272
rect 9588 31152 9640 31204
rect 11060 31220 11112 31272
rect 15568 31220 15620 31272
rect 17592 31263 17644 31272
rect 17592 31229 17601 31263
rect 17601 31229 17635 31263
rect 17635 31229 17644 31263
rect 17592 31220 17644 31229
rect 2504 31084 2556 31136
rect 5448 31084 5500 31136
rect 10416 31084 10468 31136
rect 12072 31084 12124 31136
rect 13084 31084 13136 31136
rect 14556 31152 14608 31204
rect 13728 31084 13780 31136
rect 13820 31084 13872 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1952 30923 2004 30932
rect 1952 30889 1961 30923
rect 1961 30889 1995 30923
rect 1995 30889 2004 30923
rect 1952 30880 2004 30889
rect 7748 30923 7800 30932
rect 7748 30889 7757 30923
rect 7757 30889 7791 30923
rect 7791 30889 7800 30923
rect 7748 30880 7800 30889
rect 10692 30880 10744 30932
rect 12992 30880 13044 30932
rect 13728 30880 13780 30932
rect 15660 30880 15712 30932
rect 20812 30923 20864 30932
rect 20812 30889 20821 30923
rect 20821 30889 20855 30923
rect 20855 30889 20864 30923
rect 20812 30880 20864 30889
rect 22836 30923 22888 30932
rect 22836 30889 22845 30923
rect 22845 30889 22879 30923
rect 22879 30889 22888 30923
rect 22836 30880 22888 30889
rect 2780 30676 2832 30728
rect 5724 30744 5776 30796
rect 7380 30744 7432 30796
rect 3884 30676 3936 30728
rect 11152 30812 11204 30864
rect 13360 30812 13412 30864
rect 10416 30744 10468 30796
rect 19340 30812 19392 30864
rect 15568 30787 15620 30796
rect 15568 30753 15577 30787
rect 15577 30753 15611 30787
rect 15611 30753 15620 30787
rect 15568 30744 15620 30753
rect 15752 30787 15804 30796
rect 15752 30753 15761 30787
rect 15761 30753 15795 30787
rect 15795 30753 15804 30787
rect 15752 30744 15804 30753
rect 23848 30744 23900 30796
rect 8576 30719 8628 30728
rect 8576 30685 8585 30719
rect 8585 30685 8619 30719
rect 8619 30685 8628 30719
rect 8576 30676 8628 30685
rect 9404 30719 9456 30728
rect 9404 30685 9413 30719
rect 9413 30685 9447 30719
rect 9447 30685 9456 30719
rect 9404 30676 9456 30685
rect 10140 30676 10192 30728
rect 10600 30719 10652 30728
rect 10600 30685 10609 30719
rect 10609 30685 10643 30719
rect 10643 30685 10652 30719
rect 10600 30676 10652 30685
rect 13360 30719 13412 30728
rect 13360 30685 13369 30719
rect 13369 30685 13403 30719
rect 13403 30685 13412 30719
rect 13360 30676 13412 30685
rect 16580 30676 16632 30728
rect 17868 30676 17920 30728
rect 19984 30676 20036 30728
rect 4620 30608 4672 30660
rect 6644 30651 6696 30660
rect 6644 30617 6653 30651
rect 6653 30617 6687 30651
rect 6687 30617 6696 30651
rect 6644 30608 6696 30617
rect 7472 30608 7524 30660
rect 11152 30608 11204 30660
rect 14464 30651 14516 30660
rect 2412 30540 2464 30592
rect 3148 30540 3200 30592
rect 4160 30583 4212 30592
rect 4160 30549 4169 30583
rect 4169 30549 4203 30583
rect 4203 30549 4212 30583
rect 4160 30540 4212 30549
rect 14464 30617 14473 30651
rect 14473 30617 14507 30651
rect 14507 30617 14516 30651
rect 14464 30608 14516 30617
rect 14556 30651 14608 30660
rect 14556 30617 14565 30651
rect 14565 30617 14599 30651
rect 14599 30617 14608 30651
rect 20444 30676 20496 30728
rect 22744 30719 22796 30728
rect 22744 30685 22753 30719
rect 22753 30685 22787 30719
rect 22787 30685 22796 30719
rect 22744 30676 22796 30685
rect 23572 30719 23624 30728
rect 23572 30685 23581 30719
rect 23581 30685 23615 30719
rect 23615 30685 23624 30719
rect 23572 30676 23624 30685
rect 32404 30676 32456 30728
rect 14556 30608 14608 30617
rect 17316 30540 17368 30592
rect 20168 30583 20220 30592
rect 20168 30549 20177 30583
rect 20177 30549 20211 30583
rect 20211 30549 20220 30583
rect 20168 30540 20220 30549
rect 24032 30583 24084 30592
rect 24032 30549 24041 30583
rect 24041 30549 24075 30583
rect 24075 30549 24084 30583
rect 24032 30540 24084 30549
rect 27896 30540 27948 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 9588 30336 9640 30388
rect 5448 30268 5500 30320
rect 6920 30268 6972 30320
rect 8576 30268 8628 30320
rect 9496 30268 9548 30320
rect 10876 30311 10928 30320
rect 10876 30277 10885 30311
rect 10885 30277 10919 30311
rect 10919 30277 10928 30311
rect 10876 30268 10928 30277
rect 1768 30243 1820 30252
rect 1768 30209 1777 30243
rect 1777 30209 1811 30243
rect 1811 30209 1820 30243
rect 1768 30200 1820 30209
rect 2596 30200 2648 30252
rect 6000 30243 6052 30252
rect 6000 30209 6009 30243
rect 6009 30209 6043 30243
rect 6043 30209 6052 30243
rect 6000 30200 6052 30209
rect 4160 30132 4212 30184
rect 10692 30200 10744 30252
rect 12348 30200 12400 30252
rect 2780 30064 2832 30116
rect 7472 30107 7524 30116
rect 7472 30073 7481 30107
rect 7481 30073 7515 30107
rect 7515 30073 7524 30107
rect 7472 30064 7524 30073
rect 11336 30132 11388 30184
rect 14096 30200 14148 30252
rect 11060 30064 11112 30116
rect 1584 30039 1636 30048
rect 1584 30005 1593 30039
rect 1593 30005 1627 30039
rect 1627 30005 1636 30039
rect 1584 29996 1636 30005
rect 6368 29996 6420 30048
rect 9312 30039 9364 30048
rect 9312 30005 9321 30039
rect 9321 30005 9355 30039
rect 9355 30005 9364 30039
rect 9312 29996 9364 30005
rect 9496 29996 9548 30048
rect 14188 30132 14240 30184
rect 16764 30268 16816 30320
rect 17592 30311 17644 30320
rect 17592 30277 17601 30311
rect 17601 30277 17635 30311
rect 17635 30277 17644 30311
rect 17592 30268 17644 30277
rect 34520 30268 34572 30320
rect 17868 30200 17920 30252
rect 21916 30200 21968 30252
rect 22468 30200 22520 30252
rect 30472 30200 30524 30252
rect 31760 30200 31812 30252
rect 11704 30064 11756 30116
rect 14280 30064 14332 30116
rect 11520 29996 11572 30048
rect 13176 29996 13228 30048
rect 13912 30039 13964 30048
rect 13912 30005 13921 30039
rect 13921 30005 13955 30039
rect 13955 30005 13964 30039
rect 13912 29996 13964 30005
rect 18972 29996 19024 30048
rect 21640 29996 21692 30048
rect 38200 30039 38252 30048
rect 38200 30005 38209 30039
rect 38209 30005 38243 30039
rect 38243 30005 38252 30039
rect 38200 29996 38252 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 6644 29792 6696 29844
rect 6920 29835 6972 29844
rect 6920 29801 6929 29835
rect 6929 29801 6963 29835
rect 6963 29801 6972 29835
rect 6920 29792 6972 29801
rect 9128 29792 9180 29844
rect 2780 29699 2832 29708
rect 2780 29665 2789 29699
rect 2789 29665 2823 29699
rect 2823 29665 2832 29699
rect 3056 29699 3108 29708
rect 2780 29656 2832 29665
rect 3056 29665 3065 29699
rect 3065 29665 3099 29699
rect 3099 29665 3108 29699
rect 3056 29656 3108 29665
rect 6000 29656 6052 29708
rect 9312 29699 9364 29708
rect 1860 29631 1912 29640
rect 1860 29597 1869 29631
rect 1869 29597 1903 29631
rect 1903 29597 1912 29631
rect 1860 29588 1912 29597
rect 3976 29631 4028 29640
rect 3976 29597 3985 29631
rect 3985 29597 4019 29631
rect 4019 29597 4028 29631
rect 3976 29588 4028 29597
rect 6368 29631 6420 29640
rect 6368 29597 6377 29631
rect 6377 29597 6411 29631
rect 6411 29597 6420 29631
rect 6368 29588 6420 29597
rect 9312 29665 9321 29699
rect 9321 29665 9355 29699
rect 9355 29665 9364 29699
rect 9312 29656 9364 29665
rect 11520 29699 11572 29708
rect 11520 29665 11529 29699
rect 11529 29665 11563 29699
rect 11563 29665 11572 29699
rect 11520 29656 11572 29665
rect 12992 29656 13044 29708
rect 20444 29792 20496 29844
rect 21364 29792 21416 29844
rect 23572 29792 23624 29844
rect 23848 29835 23900 29844
rect 23848 29801 23857 29835
rect 23857 29801 23891 29835
rect 23891 29801 23900 29835
rect 23848 29792 23900 29801
rect 7748 29588 7800 29640
rect 9128 29631 9180 29640
rect 9128 29597 9137 29631
rect 9137 29597 9171 29631
rect 9171 29597 9180 29631
rect 9128 29588 9180 29597
rect 11244 29588 11296 29640
rect 14280 29631 14332 29640
rect 2872 29563 2924 29572
rect 2872 29529 2881 29563
rect 2881 29529 2915 29563
rect 2915 29529 2924 29563
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 17316 29631 17368 29640
rect 17316 29597 17325 29631
rect 17325 29597 17359 29631
rect 17359 29597 17368 29631
rect 17316 29588 17368 29597
rect 19156 29588 19208 29640
rect 20168 29656 20220 29708
rect 21640 29699 21692 29708
rect 21640 29665 21649 29699
rect 21649 29665 21683 29699
rect 21683 29665 21692 29699
rect 21640 29656 21692 29665
rect 20628 29588 20680 29640
rect 20996 29588 21048 29640
rect 23020 29631 23072 29640
rect 2872 29520 2924 29529
rect 11520 29520 11572 29572
rect 2136 29452 2188 29504
rect 7564 29495 7616 29504
rect 7564 29461 7573 29495
rect 7573 29461 7607 29495
rect 7607 29461 7616 29495
rect 7564 29452 7616 29461
rect 10508 29452 10560 29504
rect 12072 29452 12124 29504
rect 12808 29520 12860 29572
rect 23020 29597 23029 29631
rect 23029 29597 23063 29631
rect 23063 29597 23072 29631
rect 23020 29588 23072 29597
rect 23756 29631 23808 29640
rect 23756 29597 23765 29631
rect 23765 29597 23799 29631
rect 23799 29597 23808 29631
rect 23756 29588 23808 29597
rect 24032 29520 24084 29572
rect 14372 29495 14424 29504
rect 14372 29461 14381 29495
rect 14381 29461 14415 29495
rect 14415 29461 14424 29495
rect 14372 29452 14424 29461
rect 17132 29495 17184 29504
rect 17132 29461 17141 29495
rect 17141 29461 17175 29495
rect 17175 29461 17184 29495
rect 17132 29452 17184 29461
rect 20076 29495 20128 29504
rect 20076 29461 20085 29495
rect 20085 29461 20119 29495
rect 20119 29461 20128 29495
rect 20076 29452 20128 29461
rect 22192 29452 22244 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 9128 29248 9180 29300
rect 12348 29291 12400 29300
rect 12348 29257 12357 29291
rect 12357 29257 12391 29291
rect 12391 29257 12400 29291
rect 12348 29248 12400 29257
rect 12532 29248 12584 29300
rect 12808 29248 12860 29300
rect 14464 29248 14516 29300
rect 36452 29248 36504 29300
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 2320 29112 2372 29164
rect 2596 29044 2648 29096
rect 8576 29180 8628 29232
rect 10600 29223 10652 29232
rect 10600 29189 10609 29223
rect 10609 29189 10643 29223
rect 10643 29189 10652 29223
rect 10600 29180 10652 29189
rect 5540 29112 5592 29164
rect 9864 29155 9916 29164
rect 8208 29044 8260 29096
rect 6828 28976 6880 29028
rect 9864 29121 9873 29155
rect 9873 29121 9907 29155
rect 9907 29121 9916 29155
rect 9864 29112 9916 29121
rect 11336 29112 11388 29164
rect 12440 29112 12492 29164
rect 13176 29155 13228 29164
rect 13176 29121 13185 29155
rect 13185 29121 13219 29155
rect 13219 29121 13228 29155
rect 13176 29112 13228 29121
rect 14096 29112 14148 29164
rect 16856 29112 16908 29164
rect 18972 29155 19024 29164
rect 18972 29121 18981 29155
rect 18981 29121 19015 29155
rect 19015 29121 19024 29155
rect 18972 29112 19024 29121
rect 25320 29155 25372 29164
rect 25320 29121 25329 29155
rect 25329 29121 25363 29155
rect 25363 29121 25372 29155
rect 25320 29112 25372 29121
rect 27988 29112 28040 29164
rect 36636 29112 36688 29164
rect 10508 29087 10560 29096
rect 10508 29053 10517 29087
rect 10517 29053 10551 29087
rect 10551 29053 10560 29087
rect 10508 29044 10560 29053
rect 10692 29044 10744 29096
rect 12992 29087 13044 29096
rect 12992 29053 13001 29087
rect 13001 29053 13035 29087
rect 13035 29053 13044 29087
rect 12992 29044 13044 29053
rect 20076 29044 20128 29096
rect 24216 29087 24268 29096
rect 24216 29053 24225 29087
rect 24225 29053 24259 29087
rect 24259 29053 24268 29087
rect 24216 29044 24268 29053
rect 19156 29019 19208 29028
rect 19156 28985 19165 29019
rect 19165 28985 19199 29019
rect 19199 28985 19208 29019
rect 19156 28976 19208 28985
rect 38200 29019 38252 29028
rect 38200 28985 38209 29019
rect 38209 28985 38243 29019
rect 38243 28985 38252 29019
rect 38200 28976 38252 28985
rect 1952 28908 2004 28960
rect 15016 28951 15068 28960
rect 15016 28917 15025 28951
rect 15025 28917 15059 28951
rect 15059 28917 15068 28951
rect 15016 28908 15068 28917
rect 16028 28951 16080 28960
rect 16028 28917 16037 28951
rect 16037 28917 16071 28951
rect 16071 28917 16080 28951
rect 16028 28908 16080 28917
rect 24676 28951 24728 28960
rect 24676 28917 24685 28951
rect 24685 28917 24719 28951
rect 24719 28917 24728 28951
rect 24676 28908 24728 28917
rect 24952 28908 25004 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 10600 28747 10652 28756
rect 10600 28713 10609 28747
rect 10609 28713 10643 28747
rect 10643 28713 10652 28747
rect 10600 28704 10652 28713
rect 16856 28747 16908 28756
rect 16856 28713 16865 28747
rect 16865 28713 16899 28747
rect 16899 28713 16908 28747
rect 16856 28704 16908 28713
rect 20076 28747 20128 28756
rect 20076 28713 20085 28747
rect 20085 28713 20119 28747
rect 20119 28713 20128 28747
rect 20076 28704 20128 28713
rect 24216 28704 24268 28756
rect 17592 28636 17644 28688
rect 3516 28568 3568 28620
rect 9220 28611 9272 28620
rect 1952 28543 2004 28552
rect 1952 28509 1961 28543
rect 1961 28509 1995 28543
rect 1995 28509 2004 28543
rect 1952 28500 2004 28509
rect 5080 28500 5132 28552
rect 9220 28577 9229 28611
rect 9229 28577 9263 28611
rect 9263 28577 9272 28611
rect 9220 28568 9272 28577
rect 12992 28568 13044 28620
rect 15660 28568 15712 28620
rect 16028 28568 16080 28620
rect 24584 28568 24636 28620
rect 9864 28500 9916 28552
rect 10876 28500 10928 28552
rect 8208 28432 8260 28484
rect 1952 28364 2004 28416
rect 5356 28364 5408 28416
rect 5448 28407 5500 28416
rect 5448 28373 5457 28407
rect 5457 28373 5491 28407
rect 5491 28373 5500 28407
rect 5448 28364 5500 28373
rect 5632 28364 5684 28416
rect 14464 28500 14516 28552
rect 15844 28500 15896 28552
rect 22008 28543 22060 28552
rect 14832 28432 14884 28484
rect 19432 28432 19484 28484
rect 22008 28509 22017 28543
rect 22017 28509 22051 28543
rect 22051 28509 22060 28543
rect 22008 28500 22060 28509
rect 24952 28543 25004 28552
rect 24952 28509 24961 28543
rect 24961 28509 24995 28543
rect 24995 28509 25004 28543
rect 24952 28500 25004 28509
rect 15752 28364 15804 28416
rect 19340 28364 19392 28416
rect 20812 28364 20864 28416
rect 21824 28407 21876 28416
rect 21824 28373 21833 28407
rect 21833 28373 21867 28407
rect 21867 28373 21876 28407
rect 21824 28364 21876 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 3056 28160 3108 28212
rect 3148 28135 3200 28144
rect 3148 28101 3157 28135
rect 3157 28101 3191 28135
rect 3191 28101 3200 28135
rect 3148 28092 3200 28101
rect 5448 28160 5500 28212
rect 14832 28203 14884 28212
rect 3792 28092 3844 28144
rect 9588 28092 9640 28144
rect 13912 28092 13964 28144
rect 1584 28024 1636 28076
rect 5356 28024 5408 28076
rect 14832 28169 14841 28203
rect 14841 28169 14875 28203
rect 14875 28169 14884 28203
rect 14832 28160 14884 28169
rect 19156 28160 19208 28212
rect 19432 28203 19484 28212
rect 19432 28169 19441 28203
rect 19441 28169 19475 28203
rect 19475 28169 19484 28203
rect 19432 28160 19484 28169
rect 22744 28160 22796 28212
rect 24032 28160 24084 28212
rect 24676 28160 24728 28212
rect 14464 28092 14516 28144
rect 15016 28067 15068 28076
rect 3056 27999 3108 28008
rect 3056 27965 3065 27999
rect 3065 27965 3099 27999
rect 3099 27965 3108 27999
rect 3056 27956 3108 27965
rect 3516 27956 3568 28008
rect 5816 27956 5868 28008
rect 14372 27956 14424 28008
rect 15016 28033 15025 28067
rect 15025 28033 15059 28067
rect 15059 28033 15068 28067
rect 15016 28024 15068 28033
rect 15568 28024 15620 28076
rect 15844 28024 15896 28076
rect 20536 28092 20588 28144
rect 16764 27956 16816 28008
rect 17132 28024 17184 28076
rect 19432 28024 19484 28076
rect 19984 28024 20036 28076
rect 20812 28067 20864 28076
rect 20812 28033 20821 28067
rect 20821 28033 20855 28067
rect 20855 28033 20864 28067
rect 20812 28024 20864 28033
rect 21824 28024 21876 28076
rect 29736 28092 29788 28144
rect 23020 28067 23072 28076
rect 23020 28033 23029 28067
rect 23029 28033 23063 28067
rect 23063 28033 23072 28067
rect 23020 28024 23072 28033
rect 25044 28067 25096 28076
rect 25044 28033 25053 28067
rect 25053 28033 25087 28067
rect 25087 28033 25096 28067
rect 25044 28024 25096 28033
rect 18144 27999 18196 28008
rect 3332 27820 3384 27872
rect 5908 27820 5960 27872
rect 17040 27888 17092 27940
rect 18144 27965 18153 27999
rect 18153 27965 18187 27999
rect 18187 27965 18196 27999
rect 18144 27956 18196 27965
rect 23848 27999 23900 28008
rect 23848 27965 23857 27999
rect 23857 27965 23891 27999
rect 23891 27965 23900 27999
rect 23848 27956 23900 27965
rect 25228 27999 25280 28008
rect 25228 27965 25237 27999
rect 25237 27965 25271 27999
rect 25271 27965 25280 27999
rect 25228 27956 25280 27965
rect 27160 27888 27212 27940
rect 15752 27820 15804 27872
rect 17408 27820 17460 27872
rect 20812 27820 20864 27872
rect 23572 27820 23624 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 13728 27616 13780 27668
rect 3976 27548 4028 27600
rect 19432 27616 19484 27668
rect 22008 27616 22060 27668
rect 23940 27616 23992 27668
rect 24584 27616 24636 27668
rect 25228 27616 25280 27668
rect 5632 27480 5684 27532
rect 5816 27523 5868 27532
rect 5816 27489 5825 27523
rect 5825 27489 5859 27523
rect 5859 27489 5868 27523
rect 5816 27480 5868 27489
rect 19340 27548 19392 27600
rect 19984 27548 20036 27600
rect 20536 27591 20588 27600
rect 20536 27557 20545 27591
rect 20545 27557 20579 27591
rect 20579 27557 20588 27591
rect 20536 27548 20588 27557
rect 23848 27548 23900 27600
rect 1768 27455 1820 27464
rect 1768 27421 1777 27455
rect 1777 27421 1811 27455
rect 1811 27421 1820 27455
rect 1768 27412 1820 27421
rect 9128 27412 9180 27464
rect 4068 27387 4120 27396
rect 4068 27353 4077 27387
rect 4077 27353 4111 27387
rect 4111 27353 4120 27387
rect 4068 27344 4120 27353
rect 4344 27344 4396 27396
rect 5908 27387 5960 27396
rect 5908 27353 5917 27387
rect 5917 27353 5951 27387
rect 5951 27353 5960 27387
rect 5908 27344 5960 27353
rect 6184 27344 6236 27396
rect 6460 27387 6512 27396
rect 6460 27353 6469 27387
rect 6469 27353 6503 27387
rect 6503 27353 6512 27387
rect 6460 27344 6512 27353
rect 11888 27344 11940 27396
rect 4252 27276 4304 27328
rect 12164 27276 12216 27328
rect 14648 27480 14700 27532
rect 16488 27412 16540 27464
rect 17040 27455 17092 27464
rect 17040 27421 17049 27455
rect 17049 27421 17083 27455
rect 17083 27421 17092 27455
rect 17040 27412 17092 27421
rect 17408 27480 17460 27532
rect 18144 27480 18196 27532
rect 20812 27480 20864 27532
rect 20720 27455 20772 27464
rect 20720 27421 20729 27455
rect 20729 27421 20763 27455
rect 20763 27421 20772 27455
rect 20720 27412 20772 27421
rect 21180 27412 21232 27464
rect 23572 27455 23624 27464
rect 23572 27421 23581 27455
rect 23581 27421 23615 27455
rect 23615 27421 23624 27455
rect 23572 27412 23624 27421
rect 30380 27548 30432 27600
rect 25228 27455 25280 27464
rect 25228 27421 25237 27455
rect 25237 27421 25271 27455
rect 25271 27421 25280 27455
rect 25228 27412 25280 27421
rect 27436 27455 27488 27464
rect 14924 27344 14976 27396
rect 27436 27421 27445 27455
rect 27445 27421 27479 27455
rect 27479 27421 27488 27455
rect 27436 27412 27488 27421
rect 37740 27412 37792 27464
rect 26240 27344 26292 27396
rect 12808 27276 12860 27328
rect 14004 27276 14056 27328
rect 16212 27319 16264 27328
rect 16212 27285 16221 27319
rect 16221 27285 16255 27319
rect 16255 27285 16264 27319
rect 16212 27276 16264 27285
rect 16856 27319 16908 27328
rect 16856 27285 16865 27319
rect 16865 27285 16899 27319
rect 16899 27285 16908 27319
rect 16856 27276 16908 27285
rect 24584 27276 24636 27328
rect 24768 27276 24820 27328
rect 27252 27276 27304 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4344 27115 4396 27124
rect 4344 27081 4353 27115
rect 4353 27081 4387 27115
rect 4387 27081 4396 27115
rect 4344 27072 4396 27081
rect 6644 27004 6696 27056
rect 12716 27072 12768 27124
rect 10968 27004 11020 27056
rect 11152 27004 11204 27056
rect 12532 27047 12584 27056
rect 12532 27013 12541 27047
rect 12541 27013 12575 27047
rect 12575 27013 12584 27047
rect 12532 27004 12584 27013
rect 1676 26936 1728 26988
rect 4252 26979 4304 26988
rect 4252 26945 4261 26979
rect 4261 26945 4295 26979
rect 4295 26945 4304 26979
rect 4252 26936 4304 26945
rect 10048 26911 10100 26920
rect 1860 26775 1912 26784
rect 1860 26741 1869 26775
rect 1869 26741 1903 26775
rect 1903 26741 1912 26775
rect 1860 26732 1912 26741
rect 10048 26877 10057 26911
rect 10057 26877 10091 26911
rect 10091 26877 10100 26911
rect 10048 26868 10100 26877
rect 12808 26936 12860 26988
rect 9312 26800 9364 26852
rect 14556 27072 14608 27124
rect 20720 27072 20772 27124
rect 22560 27072 22612 27124
rect 25228 27072 25280 27124
rect 15936 27004 15988 27056
rect 16396 26936 16448 26988
rect 22928 27004 22980 27056
rect 24768 27047 24820 27056
rect 24768 27013 24777 27047
rect 24777 27013 24811 27047
rect 24811 27013 24820 27047
rect 24768 27004 24820 27013
rect 12992 26911 13044 26920
rect 12992 26877 13001 26911
rect 13001 26877 13035 26911
rect 13035 26877 13044 26911
rect 13268 26911 13320 26920
rect 12992 26868 13044 26877
rect 13268 26877 13277 26911
rect 13277 26877 13311 26911
rect 13311 26877 13320 26911
rect 13268 26868 13320 26877
rect 13728 26868 13780 26920
rect 14556 26868 14608 26920
rect 19432 26936 19484 26988
rect 20260 26979 20312 26988
rect 20260 26945 20269 26979
rect 20269 26945 20303 26979
rect 20303 26945 20312 26979
rect 20260 26936 20312 26945
rect 21088 26936 21140 26988
rect 37280 26936 37332 26988
rect 38292 26979 38344 26988
rect 38292 26945 38301 26979
rect 38301 26945 38335 26979
rect 38335 26945 38344 26979
rect 38292 26936 38344 26945
rect 17316 26911 17368 26920
rect 17316 26877 17325 26911
rect 17325 26877 17359 26911
rect 17359 26877 17368 26911
rect 17316 26868 17368 26877
rect 17408 26868 17460 26920
rect 20720 26868 20772 26920
rect 16120 26800 16172 26852
rect 24492 26868 24544 26920
rect 24676 26911 24728 26920
rect 24676 26877 24685 26911
rect 24685 26877 24719 26911
rect 24719 26877 24728 26911
rect 24676 26868 24728 26877
rect 24124 26800 24176 26852
rect 31760 26800 31812 26852
rect 8300 26732 8352 26784
rect 10784 26732 10836 26784
rect 13820 26732 13872 26784
rect 14740 26775 14792 26784
rect 14740 26741 14749 26775
rect 14749 26741 14783 26775
rect 14783 26741 14792 26775
rect 14740 26732 14792 26741
rect 14832 26732 14884 26784
rect 19616 26732 19668 26784
rect 20812 26732 20864 26784
rect 25964 26732 26016 26784
rect 37280 26732 37332 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3056 26528 3108 26580
rect 16488 26503 16540 26512
rect 16488 26469 16497 26503
rect 16497 26469 16531 26503
rect 16531 26469 16540 26503
rect 16488 26460 16540 26469
rect 1860 26435 1912 26444
rect 1860 26401 1869 26435
rect 1869 26401 1903 26435
rect 1903 26401 1912 26435
rect 1860 26392 1912 26401
rect 2504 26392 2556 26444
rect 8300 26392 8352 26444
rect 9128 26392 9180 26444
rect 13176 26392 13228 26444
rect 14556 26435 14608 26444
rect 14556 26401 14565 26435
rect 14565 26401 14599 26435
rect 14599 26401 14608 26435
rect 14556 26392 14608 26401
rect 3148 26367 3200 26376
rect 3148 26333 3157 26367
rect 3157 26333 3191 26367
rect 3191 26333 3200 26367
rect 3148 26324 3200 26333
rect 9312 26324 9364 26376
rect 10784 26324 10836 26376
rect 2964 26231 3016 26240
rect 2964 26197 2973 26231
rect 2973 26197 3007 26231
rect 3007 26197 3016 26231
rect 2964 26188 3016 26197
rect 9772 26188 9824 26240
rect 11428 26299 11480 26308
rect 11428 26265 11437 26299
rect 11437 26265 11471 26299
rect 11471 26265 11480 26299
rect 11428 26256 11480 26265
rect 12164 26299 12216 26308
rect 12164 26265 12173 26299
rect 12173 26265 12207 26299
rect 12207 26265 12216 26299
rect 12164 26256 12216 26265
rect 12900 26256 12952 26308
rect 15016 26256 15068 26308
rect 16580 26324 16632 26376
rect 18696 26460 18748 26512
rect 19432 26460 19484 26512
rect 22744 26460 22796 26512
rect 24584 26503 24636 26512
rect 24584 26469 24593 26503
rect 24593 26469 24627 26503
rect 24627 26469 24636 26503
rect 24584 26460 24636 26469
rect 27804 26528 27856 26580
rect 17316 26435 17368 26444
rect 17316 26401 17325 26435
rect 17325 26401 17359 26435
rect 17359 26401 17368 26435
rect 17316 26392 17368 26401
rect 17592 26435 17644 26444
rect 17592 26401 17601 26435
rect 17601 26401 17635 26435
rect 17635 26401 17644 26435
rect 17592 26392 17644 26401
rect 16120 26256 16172 26308
rect 16212 26256 16264 26308
rect 19616 26299 19668 26308
rect 19616 26265 19625 26299
rect 19625 26265 19659 26299
rect 19659 26265 19668 26299
rect 20628 26435 20680 26444
rect 20628 26401 20637 26435
rect 20637 26401 20671 26435
rect 20671 26401 20680 26435
rect 20812 26435 20864 26444
rect 20628 26392 20680 26401
rect 20812 26401 20821 26435
rect 20821 26401 20855 26435
rect 20855 26401 20864 26435
rect 20812 26392 20864 26401
rect 27896 26435 27948 26444
rect 27896 26401 27905 26435
rect 27905 26401 27939 26435
rect 27939 26401 27948 26435
rect 27896 26392 27948 26401
rect 37372 26392 37424 26444
rect 21272 26367 21324 26376
rect 21272 26333 21281 26367
rect 21281 26333 21315 26367
rect 21315 26333 21324 26367
rect 21272 26324 21324 26333
rect 22100 26367 22152 26376
rect 22100 26333 22109 26367
rect 22109 26333 22143 26367
rect 22143 26333 22152 26367
rect 22100 26324 22152 26333
rect 22284 26324 22336 26376
rect 19616 26256 19668 26265
rect 22192 26256 22244 26308
rect 24492 26256 24544 26308
rect 27344 26324 27396 26376
rect 27620 26188 27672 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 3056 25984 3108 26036
rect 2412 25848 2464 25900
rect 5264 25984 5316 26036
rect 5356 25848 5408 25900
rect 9036 25984 9088 26036
rect 11428 25984 11480 26036
rect 12348 25984 12400 26036
rect 15016 25984 15068 26036
rect 22100 25984 22152 26036
rect 8208 25916 8260 25968
rect 14372 25916 14424 25968
rect 14648 25916 14700 25968
rect 16856 25916 16908 25968
rect 19340 25959 19392 25968
rect 19340 25925 19349 25959
rect 19349 25925 19383 25959
rect 19383 25925 19392 25959
rect 19340 25916 19392 25925
rect 28540 25916 28592 25968
rect 10048 25848 10100 25900
rect 1860 25823 1912 25832
rect 1860 25789 1869 25823
rect 1869 25789 1903 25823
rect 1903 25789 1912 25823
rect 1860 25780 1912 25789
rect 2228 25780 2280 25832
rect 3976 25823 4028 25832
rect 3976 25789 3985 25823
rect 3985 25789 4019 25823
rect 4019 25789 4028 25823
rect 3976 25780 4028 25789
rect 10600 25780 10652 25832
rect 11704 25780 11756 25832
rect 16212 25848 16264 25900
rect 16396 25848 16448 25900
rect 20720 25848 20772 25900
rect 21180 25848 21232 25900
rect 22376 25848 22428 25900
rect 27068 25848 27120 25900
rect 27160 25891 27212 25900
rect 27160 25857 27169 25891
rect 27169 25857 27203 25891
rect 27203 25857 27212 25891
rect 27160 25848 27212 25857
rect 29460 25891 29512 25900
rect 18512 25823 18564 25832
rect 18512 25789 18521 25823
rect 18521 25789 18555 25823
rect 18555 25789 18564 25823
rect 18512 25780 18564 25789
rect 19248 25823 19300 25832
rect 19248 25789 19257 25823
rect 19257 25789 19291 25823
rect 19291 25789 19300 25823
rect 19248 25780 19300 25789
rect 19524 25823 19576 25832
rect 19524 25789 19533 25823
rect 19533 25789 19567 25823
rect 19567 25789 19576 25823
rect 19524 25780 19576 25789
rect 29460 25857 29469 25891
rect 29469 25857 29503 25891
rect 29503 25857 29512 25891
rect 29460 25848 29512 25857
rect 17592 25712 17644 25764
rect 38108 25780 38160 25832
rect 3424 25687 3476 25696
rect 3424 25653 3433 25687
rect 3433 25653 3467 25687
rect 3467 25653 3476 25687
rect 3424 25644 3476 25653
rect 11152 25644 11204 25696
rect 16028 25644 16080 25696
rect 20628 25687 20680 25696
rect 20628 25653 20637 25687
rect 20637 25653 20671 25687
rect 20671 25653 20680 25687
rect 20628 25644 20680 25653
rect 23480 25644 23532 25696
rect 27620 25687 27672 25696
rect 27620 25653 27629 25687
rect 27629 25653 27663 25687
rect 27663 25653 27672 25687
rect 27620 25644 27672 25653
rect 28172 25644 28224 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3792 25440 3844 25492
rect 5356 25440 5408 25492
rect 13728 25440 13780 25492
rect 20260 25440 20312 25492
rect 22376 25483 22428 25492
rect 22376 25449 22385 25483
rect 22385 25449 22419 25483
rect 22419 25449 22428 25483
rect 22376 25440 22428 25449
rect 27068 25483 27120 25492
rect 27068 25449 27077 25483
rect 27077 25449 27111 25483
rect 27111 25449 27120 25483
rect 27068 25440 27120 25449
rect 36636 25440 36688 25492
rect 38108 25483 38160 25492
rect 38108 25449 38117 25483
rect 38117 25449 38151 25483
rect 38151 25449 38160 25483
rect 38108 25440 38160 25449
rect 3516 25372 3568 25424
rect 2964 25304 3016 25356
rect 3332 25304 3384 25356
rect 9128 25347 9180 25356
rect 9128 25313 9137 25347
rect 9137 25313 9171 25347
rect 9171 25313 9180 25347
rect 9128 25304 9180 25313
rect 10968 25372 11020 25424
rect 19524 25372 19576 25424
rect 19248 25304 19300 25356
rect 26240 25304 26292 25356
rect 28540 25347 28592 25356
rect 28540 25313 28549 25347
rect 28549 25313 28583 25347
rect 28583 25313 28592 25347
rect 28540 25304 28592 25313
rect 2504 25236 2556 25288
rect 8208 25236 8260 25288
rect 16396 25236 16448 25288
rect 20536 25236 20588 25288
rect 20904 25279 20956 25288
rect 20904 25245 20913 25279
rect 20913 25245 20947 25279
rect 20947 25245 20956 25279
rect 20904 25236 20956 25245
rect 22928 25236 22980 25288
rect 23572 25279 23624 25288
rect 23572 25245 23581 25279
rect 23581 25245 23615 25279
rect 23615 25245 23624 25279
rect 23572 25236 23624 25245
rect 24492 25236 24544 25288
rect 27160 25236 27212 25288
rect 27344 25236 27396 25288
rect 27804 25236 27856 25288
rect 29000 25236 29052 25288
rect 38292 25279 38344 25288
rect 3332 25168 3384 25220
rect 3700 25168 3752 25220
rect 2688 25143 2740 25152
rect 2688 25109 2697 25143
rect 2697 25109 2731 25143
rect 2731 25109 2740 25143
rect 2688 25100 2740 25109
rect 3424 25100 3476 25152
rect 9036 25168 9088 25220
rect 14832 25168 14884 25220
rect 28908 25168 28960 25220
rect 38292 25245 38301 25279
rect 38301 25245 38335 25279
rect 38335 25245 38344 25279
rect 38292 25236 38344 25245
rect 5448 25100 5500 25152
rect 10876 25143 10928 25152
rect 10876 25109 10885 25143
rect 10885 25109 10919 25143
rect 10919 25109 10928 25143
rect 10876 25100 10928 25109
rect 20996 25100 21048 25152
rect 24032 25143 24084 25152
rect 24032 25109 24041 25143
rect 24041 25109 24075 25143
rect 24075 25109 24084 25143
rect 24032 25100 24084 25109
rect 25320 25100 25372 25152
rect 27712 25143 27764 25152
rect 27712 25109 27721 25143
rect 27721 25109 27755 25143
rect 27755 25109 27764 25143
rect 27712 25100 27764 25109
rect 29828 25100 29880 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 19340 24896 19392 24948
rect 24032 24896 24084 24948
rect 17224 24871 17276 24880
rect 17224 24837 17233 24871
rect 17233 24837 17267 24871
rect 17267 24837 17276 24871
rect 17224 24828 17276 24837
rect 25320 24871 25372 24880
rect 25320 24837 25329 24871
rect 25329 24837 25363 24871
rect 25363 24837 25372 24871
rect 25320 24828 25372 24837
rect 7564 24760 7616 24812
rect 11704 24760 11756 24812
rect 16028 24760 16080 24812
rect 16120 24803 16172 24812
rect 16120 24769 16129 24803
rect 16129 24769 16163 24803
rect 16163 24769 16172 24803
rect 16120 24760 16172 24769
rect 20628 24760 20680 24812
rect 20996 24803 21048 24812
rect 20996 24769 21005 24803
rect 21005 24769 21039 24803
rect 21039 24769 21048 24803
rect 20996 24760 21048 24769
rect 22928 24760 22980 24812
rect 23480 24803 23532 24812
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 27988 24760 28040 24812
rect 28356 24760 28408 24812
rect 28632 24760 28684 24812
rect 2596 24692 2648 24744
rect 9772 24692 9824 24744
rect 13176 24692 13228 24744
rect 12992 24624 13044 24676
rect 15936 24692 15988 24744
rect 15660 24624 15712 24676
rect 17040 24624 17092 24676
rect 23388 24692 23440 24744
rect 23940 24692 23992 24744
rect 24032 24692 24084 24744
rect 29552 24692 29604 24744
rect 30472 24735 30524 24744
rect 30472 24701 30481 24735
rect 30481 24701 30515 24735
rect 30515 24701 30524 24735
rect 30472 24692 30524 24701
rect 23572 24624 23624 24676
rect 2780 24556 2832 24608
rect 3516 24599 3568 24608
rect 3516 24565 3525 24599
rect 3525 24565 3559 24599
rect 3559 24565 3568 24599
rect 3516 24556 3568 24565
rect 15936 24556 15988 24608
rect 20812 24599 20864 24608
rect 20812 24565 20821 24599
rect 20821 24565 20855 24599
rect 20855 24565 20864 24599
rect 20812 24556 20864 24565
rect 29920 24556 29972 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1768 24395 1820 24404
rect 1768 24361 1777 24395
rect 1777 24361 1811 24395
rect 1811 24361 1820 24395
rect 1768 24352 1820 24361
rect 4068 24395 4120 24404
rect 4068 24361 4077 24395
rect 4077 24361 4111 24395
rect 4111 24361 4120 24395
rect 4068 24352 4120 24361
rect 5908 24352 5960 24404
rect 13636 24352 13688 24404
rect 13728 24352 13780 24404
rect 15936 24352 15988 24404
rect 22284 24352 22336 24404
rect 29000 24395 29052 24404
rect 6644 24327 6696 24336
rect 6644 24293 6653 24327
rect 6653 24293 6687 24327
rect 6687 24293 6696 24327
rect 6644 24284 6696 24293
rect 1860 24216 1912 24268
rect 20352 24216 20404 24268
rect 20812 24259 20864 24268
rect 20812 24225 20821 24259
rect 20821 24225 20855 24259
rect 20855 24225 20864 24259
rect 20812 24216 20864 24225
rect 20904 24216 20956 24268
rect 21548 24216 21600 24268
rect 1952 24148 2004 24200
rect 2872 24148 2924 24200
rect 4068 24148 4120 24200
rect 7748 24148 7800 24200
rect 15292 24148 15344 24200
rect 16120 24148 16172 24200
rect 16396 24191 16448 24200
rect 16396 24157 16405 24191
rect 16405 24157 16439 24191
rect 16439 24157 16448 24191
rect 16396 24148 16448 24157
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 25412 24191 25464 24200
rect 17868 24080 17920 24132
rect 25412 24157 25421 24191
rect 25421 24157 25455 24191
rect 25455 24157 25464 24191
rect 25412 24148 25464 24157
rect 27160 24148 27212 24200
rect 5540 24012 5592 24064
rect 6184 24012 6236 24064
rect 10784 24012 10836 24064
rect 14556 24012 14608 24064
rect 15568 24012 15620 24064
rect 16120 24012 16172 24064
rect 18052 24012 18104 24064
rect 21364 24012 21416 24064
rect 22100 24123 22152 24132
rect 22100 24089 22109 24123
rect 22109 24089 22143 24123
rect 22143 24089 22152 24123
rect 22100 24080 22152 24089
rect 26332 24080 26384 24132
rect 29000 24361 29009 24395
rect 29009 24361 29043 24395
rect 29043 24361 29052 24395
rect 29000 24352 29052 24361
rect 33324 24284 33376 24336
rect 27528 24148 27580 24200
rect 22284 24012 22336 24064
rect 25136 24012 25188 24064
rect 28264 24055 28316 24064
rect 28264 24021 28273 24055
rect 28273 24021 28307 24055
rect 28307 24021 28316 24055
rect 28264 24012 28316 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 5908 23808 5960 23860
rect 13636 23808 13688 23860
rect 21180 23808 21232 23860
rect 21364 23851 21416 23860
rect 21364 23817 21373 23851
rect 21373 23817 21407 23851
rect 21407 23817 21416 23851
rect 21364 23808 21416 23817
rect 22100 23851 22152 23860
rect 22100 23817 22109 23851
rect 22109 23817 22143 23851
rect 22143 23817 22152 23851
rect 22100 23808 22152 23817
rect 5448 23740 5500 23792
rect 6828 23740 6880 23792
rect 10692 23740 10744 23792
rect 14924 23740 14976 23792
rect 27528 23808 27580 23860
rect 28356 23851 28408 23860
rect 28356 23817 28365 23851
rect 28365 23817 28399 23851
rect 28399 23817 28408 23851
rect 28356 23808 28408 23817
rect 7748 23715 7800 23724
rect 7748 23681 7757 23715
rect 7757 23681 7791 23715
rect 7791 23681 7800 23715
rect 7748 23672 7800 23681
rect 2780 23604 2832 23656
rect 3976 23604 4028 23656
rect 12348 23604 12400 23656
rect 13176 23604 13228 23656
rect 14832 23604 14884 23656
rect 3516 23536 3568 23588
rect 6736 23536 6788 23588
rect 10140 23536 10192 23588
rect 26608 23740 26660 23792
rect 27712 23740 27764 23792
rect 27988 23740 28040 23792
rect 29920 23783 29972 23792
rect 29920 23749 29929 23783
rect 29929 23749 29963 23783
rect 29963 23749 29972 23783
rect 29920 23740 29972 23749
rect 30472 23783 30524 23792
rect 30472 23749 30481 23783
rect 30481 23749 30515 23783
rect 30515 23749 30524 23783
rect 30472 23740 30524 23749
rect 15108 23672 15160 23724
rect 16396 23672 16448 23724
rect 18052 23715 18104 23724
rect 18052 23681 18061 23715
rect 18061 23681 18095 23715
rect 18095 23681 18104 23715
rect 18052 23672 18104 23681
rect 19984 23672 20036 23724
rect 20352 23715 20404 23724
rect 20352 23681 20361 23715
rect 20361 23681 20395 23715
rect 20395 23681 20404 23715
rect 20720 23715 20772 23724
rect 20352 23672 20404 23681
rect 20720 23681 20729 23715
rect 20729 23681 20763 23715
rect 20763 23681 20772 23715
rect 20720 23672 20772 23681
rect 22008 23715 22060 23724
rect 22008 23681 22017 23715
rect 22017 23681 22051 23715
rect 22051 23681 22060 23715
rect 22008 23672 22060 23681
rect 25136 23715 25188 23724
rect 25136 23681 25145 23715
rect 25145 23681 25179 23715
rect 25179 23681 25188 23715
rect 25136 23672 25188 23681
rect 26332 23715 26384 23724
rect 26332 23681 26341 23715
rect 26341 23681 26375 23715
rect 26375 23681 26384 23715
rect 28540 23715 28592 23724
rect 26332 23672 26384 23681
rect 28540 23681 28549 23715
rect 28549 23681 28583 23715
rect 28583 23681 28592 23715
rect 28540 23672 28592 23681
rect 38292 23715 38344 23724
rect 38292 23681 38301 23715
rect 38301 23681 38335 23715
rect 38335 23681 38344 23715
rect 38292 23672 38344 23681
rect 16764 23604 16816 23656
rect 16948 23604 17000 23656
rect 17868 23604 17920 23656
rect 18788 23647 18840 23656
rect 18788 23613 18797 23647
rect 18797 23613 18831 23647
rect 18831 23613 18840 23647
rect 18788 23604 18840 23613
rect 22284 23604 22336 23656
rect 23296 23647 23348 23656
rect 23296 23613 23305 23647
rect 23305 23613 23339 23647
rect 23339 23613 23348 23647
rect 23296 23604 23348 23613
rect 25228 23604 25280 23656
rect 29828 23647 29880 23656
rect 3700 23511 3752 23520
rect 3700 23477 3709 23511
rect 3709 23477 3743 23511
rect 3743 23477 3752 23511
rect 3700 23468 3752 23477
rect 5172 23468 5224 23520
rect 7840 23511 7892 23520
rect 7840 23477 7849 23511
rect 7849 23477 7883 23511
rect 7883 23477 7892 23511
rect 7840 23468 7892 23477
rect 10600 23468 10652 23520
rect 15016 23468 15068 23520
rect 21088 23536 21140 23588
rect 29828 23613 29837 23647
rect 29837 23613 29871 23647
rect 29871 23613 29880 23647
rect 29828 23604 29880 23613
rect 30104 23536 30156 23588
rect 15200 23468 15252 23520
rect 17868 23511 17920 23520
rect 17868 23477 17877 23511
rect 17877 23477 17911 23511
rect 17911 23477 17920 23511
rect 17868 23468 17920 23477
rect 18604 23468 18656 23520
rect 19708 23511 19760 23520
rect 19708 23477 19717 23511
rect 19717 23477 19751 23511
rect 19751 23477 19760 23511
rect 19708 23468 19760 23477
rect 24952 23511 25004 23520
rect 24952 23477 24961 23511
rect 24961 23477 24995 23511
rect 24995 23477 25004 23511
rect 24952 23468 25004 23477
rect 36452 23468 36504 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 5724 23307 5776 23316
rect 5724 23273 5733 23307
rect 5733 23273 5767 23307
rect 5767 23273 5776 23307
rect 5724 23264 5776 23273
rect 7380 23264 7432 23316
rect 11152 23239 11204 23248
rect 11152 23205 11161 23239
rect 11161 23205 11195 23239
rect 11195 23205 11204 23239
rect 11152 23196 11204 23205
rect 18788 23264 18840 23316
rect 26608 23307 26660 23316
rect 26608 23273 26617 23307
rect 26617 23273 26651 23307
rect 26651 23273 26660 23307
rect 26608 23264 26660 23273
rect 29828 23264 29880 23316
rect 4620 23128 4672 23180
rect 4988 23128 5040 23180
rect 1584 23103 1636 23112
rect 1584 23069 1593 23103
rect 1593 23069 1627 23103
rect 1627 23069 1636 23103
rect 1584 23060 1636 23069
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 13176 23128 13228 23180
rect 13268 23128 13320 23180
rect 19432 23196 19484 23248
rect 19800 23239 19852 23248
rect 19800 23205 19809 23239
rect 19809 23205 19843 23239
rect 19843 23205 19852 23239
rect 19800 23196 19852 23205
rect 20260 23196 20312 23248
rect 24768 23196 24820 23248
rect 14556 23060 14608 23112
rect 11796 23035 11848 23044
rect 1768 22967 1820 22976
rect 1768 22933 1777 22967
rect 1777 22933 1811 22967
rect 1811 22933 1820 22967
rect 1768 22924 1820 22933
rect 11796 23001 11805 23035
rect 11805 23001 11839 23035
rect 11839 23001 11848 23035
rect 11796 22992 11848 23001
rect 13820 22992 13872 23044
rect 15292 23060 15344 23112
rect 15660 22924 15712 22976
rect 16764 23171 16816 23180
rect 16764 23137 16773 23171
rect 16773 23137 16807 23171
rect 16807 23137 16816 23171
rect 16764 23128 16816 23137
rect 16488 23035 16540 23044
rect 16488 23001 16497 23035
rect 16497 23001 16531 23035
rect 16531 23001 16540 23035
rect 16488 22992 16540 23001
rect 17132 23060 17184 23112
rect 17960 23060 18012 23112
rect 18696 23060 18748 23112
rect 18236 22992 18288 23044
rect 19708 23128 19760 23180
rect 22192 23171 22244 23180
rect 22192 23137 22201 23171
rect 22201 23137 22235 23171
rect 22235 23137 22244 23171
rect 22192 23128 22244 23137
rect 23296 23171 23348 23180
rect 23296 23137 23305 23171
rect 23305 23137 23339 23171
rect 23339 23137 23348 23171
rect 23296 23128 23348 23137
rect 24952 23128 25004 23180
rect 19800 23060 19852 23112
rect 21364 23060 21416 23112
rect 20628 22992 20680 23044
rect 20812 22992 20864 23044
rect 22008 22992 22060 23044
rect 18696 22924 18748 22976
rect 19340 22967 19392 22976
rect 19340 22933 19349 22967
rect 19349 22933 19383 22967
rect 19383 22933 19392 22967
rect 19340 22924 19392 22933
rect 28264 23060 28316 23112
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 6460 22720 6512 22772
rect 2688 22652 2740 22704
rect 7380 22584 7432 22636
rect 7748 22584 7800 22636
rect 8208 22627 8260 22636
rect 8208 22593 8217 22627
rect 8217 22593 8251 22627
rect 8251 22593 8260 22627
rect 8208 22584 8260 22593
rect 9128 22652 9180 22704
rect 16488 22720 16540 22772
rect 17500 22695 17552 22704
rect 17500 22661 17509 22695
rect 17509 22661 17543 22695
rect 17543 22661 17552 22695
rect 17500 22652 17552 22661
rect 19984 22720 20036 22772
rect 21364 22763 21416 22772
rect 21364 22729 21373 22763
rect 21373 22729 21407 22763
rect 21407 22729 21416 22763
rect 21364 22720 21416 22729
rect 10600 22584 10652 22636
rect 15292 22584 15344 22636
rect 15568 22584 15620 22636
rect 20352 22652 20404 22704
rect 24768 22695 24820 22704
rect 24768 22661 24777 22695
rect 24777 22661 24811 22695
rect 24811 22661 24820 22695
rect 24768 22652 24820 22661
rect 27344 22695 27396 22704
rect 27344 22661 27353 22695
rect 27353 22661 27387 22695
rect 27387 22661 27396 22695
rect 27344 22652 27396 22661
rect 18696 22627 18748 22636
rect 2136 22516 2188 22568
rect 4620 22448 4672 22500
rect 18696 22593 18705 22627
rect 18705 22593 18739 22627
rect 18739 22593 18748 22627
rect 18696 22584 18748 22593
rect 20076 22584 20128 22636
rect 20628 22584 20680 22636
rect 26056 22627 26108 22636
rect 18144 22516 18196 22568
rect 26056 22593 26065 22627
rect 26065 22593 26099 22627
rect 26099 22593 26108 22627
rect 26056 22584 26108 22593
rect 25412 22516 25464 22568
rect 27620 22516 27672 22568
rect 27712 22559 27764 22568
rect 27712 22525 27721 22559
rect 27721 22525 27755 22559
rect 27755 22525 27764 22559
rect 28356 22559 28408 22568
rect 27712 22516 27764 22525
rect 28356 22525 28365 22559
rect 28365 22525 28399 22559
rect 28399 22525 28408 22559
rect 28356 22516 28408 22525
rect 12164 22448 12216 22500
rect 17776 22448 17828 22500
rect 7564 22380 7616 22432
rect 7748 22380 7800 22432
rect 9496 22380 9548 22432
rect 11796 22380 11848 22432
rect 18880 22423 18932 22432
rect 18880 22389 18889 22423
rect 18889 22389 18923 22423
rect 18923 22389 18932 22423
rect 18880 22380 18932 22389
rect 28540 22380 28592 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3700 22176 3752 22228
rect 2228 22040 2280 22092
rect 8300 22176 8352 22228
rect 9588 22176 9640 22228
rect 17776 22176 17828 22228
rect 18236 22176 18288 22228
rect 20260 22176 20312 22228
rect 26056 22219 26108 22228
rect 26056 22185 26065 22219
rect 26065 22185 26099 22219
rect 26099 22185 26108 22219
rect 26056 22176 26108 22185
rect 27344 22176 27396 22228
rect 8576 22083 8628 22092
rect 8576 22049 8585 22083
rect 8585 22049 8619 22083
rect 8619 22049 8628 22083
rect 8576 22040 8628 22049
rect 16028 22108 16080 22160
rect 20812 22108 20864 22160
rect 6552 22015 6604 22024
rect 6552 21981 6561 22015
rect 6561 21981 6595 22015
rect 6595 21981 6604 22015
rect 6552 21972 6604 21981
rect 9588 22015 9640 22024
rect 9588 21981 9597 22015
rect 9597 21981 9631 22015
rect 9631 21981 9640 22015
rect 9588 21972 9640 21981
rect 12900 22040 12952 22092
rect 13176 22040 13228 22092
rect 15936 22040 15988 22092
rect 17868 22040 17920 22092
rect 21272 22040 21324 22092
rect 28908 22151 28960 22160
rect 28908 22117 28917 22151
rect 28917 22117 28951 22151
rect 28951 22117 28960 22151
rect 28908 22108 28960 22117
rect 4620 21904 4672 21956
rect 7840 21904 7892 21956
rect 9496 21904 9548 21956
rect 11060 21904 11112 21956
rect 12532 21947 12584 21956
rect 12532 21913 12541 21947
rect 12541 21913 12575 21947
rect 12575 21913 12584 21947
rect 12532 21904 12584 21913
rect 9404 21836 9456 21888
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 11152 21836 11204 21888
rect 14464 21904 14516 21956
rect 14556 21904 14608 21956
rect 16396 21904 16448 21956
rect 19156 21972 19208 22024
rect 20168 21972 20220 22024
rect 20536 22015 20588 22024
rect 20536 21981 20545 22015
rect 20545 21981 20579 22015
rect 20579 21981 20588 22015
rect 20536 21972 20588 21981
rect 24124 22040 24176 22092
rect 28356 22083 28408 22092
rect 28356 22049 28365 22083
rect 28365 22049 28399 22083
rect 28399 22049 28408 22083
rect 28356 22040 28408 22049
rect 22376 21972 22428 22024
rect 24216 21972 24268 22024
rect 37280 22040 37332 22092
rect 15200 21836 15252 21888
rect 16672 21836 16724 21888
rect 17132 21836 17184 21888
rect 17408 21879 17460 21888
rect 17408 21845 17417 21879
rect 17417 21845 17451 21879
rect 17451 21845 17460 21879
rect 17408 21836 17460 21845
rect 18420 21836 18472 21888
rect 18604 21879 18656 21888
rect 18604 21845 18613 21879
rect 18613 21845 18647 21879
rect 18647 21845 18656 21879
rect 18604 21836 18656 21845
rect 23112 21904 23164 21956
rect 23204 21904 23256 21956
rect 20812 21836 20864 21888
rect 23572 21904 23624 21956
rect 30932 21972 30984 22024
rect 28448 21947 28500 21956
rect 28448 21913 28457 21947
rect 28457 21913 28491 21947
rect 28491 21913 28500 21947
rect 28448 21904 28500 21913
rect 30196 21879 30248 21888
rect 30196 21845 30205 21879
rect 30205 21845 30239 21879
rect 30239 21845 30248 21879
rect 30196 21836 30248 21845
rect 38200 21879 38252 21888
rect 38200 21845 38209 21879
rect 38209 21845 38243 21879
rect 38243 21845 38252 21879
rect 38200 21836 38252 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 6184 21632 6236 21684
rect 14556 21675 14608 21684
rect 4804 21564 4856 21616
rect 9404 21564 9456 21616
rect 12256 21564 12308 21616
rect 14556 21641 14565 21675
rect 14565 21641 14599 21675
rect 14599 21641 14608 21675
rect 14556 21632 14608 21641
rect 17500 21632 17552 21684
rect 20168 21675 20220 21684
rect 20168 21641 20177 21675
rect 20177 21641 20211 21675
rect 20211 21641 20220 21675
rect 20168 21632 20220 21641
rect 12532 21564 12584 21616
rect 17960 21564 18012 21616
rect 1768 21539 1820 21548
rect 1768 21505 1777 21539
rect 1777 21505 1811 21539
rect 1811 21505 1820 21539
rect 1768 21496 1820 21505
rect 13544 21496 13596 21548
rect 13820 21539 13872 21548
rect 13820 21505 13829 21539
rect 13829 21505 13863 21539
rect 13863 21505 13872 21539
rect 13820 21496 13872 21505
rect 14464 21539 14516 21548
rect 14464 21505 14473 21539
rect 14473 21505 14507 21539
rect 14507 21505 14516 21539
rect 14464 21496 14516 21505
rect 14832 21496 14884 21548
rect 17316 21496 17368 21548
rect 21916 21564 21968 21616
rect 23572 21632 23624 21684
rect 24216 21675 24268 21684
rect 24216 21641 24225 21675
rect 24225 21641 24259 21675
rect 24259 21641 24268 21675
rect 24216 21632 24268 21641
rect 29552 21675 29604 21684
rect 29552 21641 29561 21675
rect 29561 21641 29595 21675
rect 29595 21641 29604 21675
rect 29552 21632 29604 21641
rect 22192 21607 22244 21616
rect 20076 21539 20128 21548
rect 4620 21428 4672 21480
rect 6552 21471 6604 21480
rect 6552 21437 6561 21471
rect 6561 21437 6595 21471
rect 6595 21437 6604 21471
rect 6552 21428 6604 21437
rect 6276 21360 6328 21412
rect 9404 21428 9456 21480
rect 20076 21505 20085 21539
rect 20085 21505 20119 21539
rect 20119 21505 20128 21539
rect 20076 21496 20128 21505
rect 17868 21428 17920 21480
rect 20444 21428 20496 21480
rect 22192 21573 22201 21607
rect 22201 21573 22235 21607
rect 22235 21573 22244 21607
rect 22192 21564 22244 21573
rect 22836 21564 22888 21616
rect 17132 21360 17184 21412
rect 22376 21428 22428 21480
rect 2412 21292 2464 21344
rect 2780 21292 2832 21344
rect 7472 21292 7524 21344
rect 13912 21335 13964 21344
rect 13912 21301 13921 21335
rect 13921 21301 13955 21335
rect 13955 21301 13964 21335
rect 13912 21292 13964 21301
rect 14648 21292 14700 21344
rect 21088 21360 21140 21412
rect 27528 21496 27580 21548
rect 33048 21496 33100 21548
rect 19248 21292 19300 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6092 21088 6144 21140
rect 12164 21088 12216 21140
rect 14924 21088 14976 21140
rect 16396 21088 16448 21140
rect 21548 21088 21600 21140
rect 22836 21131 22888 21140
rect 22836 21097 22845 21131
rect 22845 21097 22879 21131
rect 22879 21097 22888 21131
rect 22836 21088 22888 21097
rect 28448 21088 28500 21140
rect 30932 21131 30984 21140
rect 30932 21097 30941 21131
rect 30941 21097 30975 21131
rect 30975 21097 30984 21131
rect 30932 21088 30984 21097
rect 2780 20995 2832 21004
rect 2780 20961 2789 20995
rect 2789 20961 2823 20995
rect 2823 20961 2832 20995
rect 3976 20995 4028 21004
rect 2780 20952 2832 20961
rect 3976 20961 3985 20995
rect 3985 20961 4019 20995
rect 4019 20961 4028 20995
rect 3976 20952 4028 20961
rect 4620 20952 4672 21004
rect 14096 20952 14148 21004
rect 17132 21020 17184 21072
rect 23020 21020 23072 21072
rect 29552 21020 29604 21072
rect 9496 20884 9548 20936
rect 15292 20884 15344 20936
rect 15476 20884 15528 20936
rect 18420 20952 18472 21004
rect 20720 20952 20772 21004
rect 16120 20927 16172 20936
rect 16120 20893 16129 20927
rect 16129 20893 16163 20927
rect 16163 20893 16172 20927
rect 16120 20884 16172 20893
rect 17684 20884 17736 20936
rect 19340 20884 19392 20936
rect 21456 20927 21508 20936
rect 21456 20893 21465 20927
rect 21465 20893 21499 20927
rect 21499 20893 21508 20927
rect 21456 20884 21508 20893
rect 3424 20859 3476 20868
rect 3424 20825 3433 20859
rect 3433 20825 3467 20859
rect 3467 20825 3476 20859
rect 3424 20816 3476 20825
rect 4712 20816 4764 20868
rect 9680 20816 9732 20868
rect 5632 20748 5684 20800
rect 7932 20748 7984 20800
rect 13452 20748 13504 20800
rect 16488 20748 16540 20800
rect 18512 20816 18564 20868
rect 18788 20816 18840 20868
rect 27988 20952 28040 21004
rect 23020 20927 23072 20936
rect 23020 20893 23029 20927
rect 23029 20893 23063 20927
rect 23063 20893 23072 20927
rect 23020 20884 23072 20893
rect 24768 20884 24820 20936
rect 27528 20884 27580 20936
rect 28080 20927 28132 20936
rect 28080 20893 28089 20927
rect 28089 20893 28123 20927
rect 28123 20893 28132 20927
rect 28080 20884 28132 20893
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 31116 20927 31168 20936
rect 31116 20893 31125 20927
rect 31125 20893 31159 20927
rect 31159 20893 31168 20927
rect 31116 20884 31168 20893
rect 18052 20748 18104 20800
rect 19340 20748 19392 20800
rect 23204 20748 23256 20800
rect 23572 20791 23624 20800
rect 23572 20757 23581 20791
rect 23581 20757 23615 20791
rect 23615 20757 23624 20791
rect 23572 20748 23624 20757
rect 27896 20748 27948 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1584 20544 1636 20596
rect 14740 20544 14792 20596
rect 7840 20476 7892 20528
rect 13452 20476 13504 20528
rect 1952 20451 2004 20460
rect 1952 20417 1961 20451
rect 1961 20417 1995 20451
rect 1995 20417 2004 20451
rect 1952 20408 2004 20417
rect 4620 20408 4672 20460
rect 14188 20408 14240 20460
rect 15200 20408 15252 20460
rect 16028 20544 16080 20596
rect 16304 20544 16356 20596
rect 20444 20587 20496 20596
rect 20444 20553 20453 20587
rect 20453 20553 20487 20587
rect 20487 20553 20496 20587
rect 20444 20544 20496 20553
rect 21456 20544 21508 20596
rect 28080 20544 28132 20596
rect 29920 20544 29972 20596
rect 31116 20587 31168 20596
rect 31116 20553 31125 20587
rect 31125 20553 31159 20587
rect 31159 20553 31168 20587
rect 31116 20544 31168 20553
rect 19340 20519 19392 20528
rect 19340 20485 19349 20519
rect 19349 20485 19383 20519
rect 19383 20485 19392 20519
rect 19340 20476 19392 20485
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 18236 20408 18288 20460
rect 9312 20383 9364 20392
rect 9312 20349 9321 20383
rect 9321 20349 9355 20383
rect 9355 20349 9364 20383
rect 9312 20340 9364 20349
rect 12900 20383 12952 20392
rect 12900 20349 12909 20383
rect 12909 20349 12943 20383
rect 12943 20349 12952 20383
rect 12900 20340 12952 20349
rect 3976 20204 4028 20256
rect 15568 20340 15620 20392
rect 15936 20340 15988 20392
rect 16948 20383 17000 20392
rect 16948 20349 16957 20383
rect 16957 20349 16991 20383
rect 16991 20349 17000 20383
rect 16948 20340 17000 20349
rect 15568 20247 15620 20256
rect 15568 20213 15577 20247
rect 15577 20213 15611 20247
rect 15611 20213 15620 20247
rect 15568 20204 15620 20213
rect 16948 20204 17000 20256
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 19984 20340 20036 20392
rect 21916 20408 21968 20460
rect 23572 20408 23624 20460
rect 27896 20451 27948 20460
rect 27896 20417 27905 20451
rect 27905 20417 27939 20451
rect 27939 20417 27948 20451
rect 27896 20408 27948 20417
rect 29460 20451 29512 20460
rect 29460 20417 29469 20451
rect 29469 20417 29503 20451
rect 29503 20417 29512 20451
rect 29460 20408 29512 20417
rect 30196 20408 30248 20460
rect 31024 20451 31076 20460
rect 31024 20417 31033 20451
rect 31033 20417 31067 20451
rect 31067 20417 31076 20451
rect 31024 20408 31076 20417
rect 36452 20408 36504 20460
rect 17408 20272 17460 20324
rect 22744 20340 22796 20392
rect 23112 20383 23164 20392
rect 23112 20349 23121 20383
rect 23121 20349 23155 20383
rect 23155 20349 23164 20383
rect 23112 20340 23164 20349
rect 30380 20340 30432 20392
rect 17960 20204 18012 20256
rect 22836 20204 22888 20256
rect 30472 20247 30524 20256
rect 30472 20213 30481 20247
rect 30481 20213 30515 20247
rect 30515 20213 30524 20247
rect 30472 20204 30524 20213
rect 31760 20204 31812 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2872 20000 2924 20052
rect 1768 19839 1820 19848
rect 1768 19805 1777 19839
rect 1777 19805 1811 19839
rect 1811 19805 1820 19839
rect 1768 19796 1820 19805
rect 2228 19796 2280 19848
rect 11060 20000 11112 20052
rect 13912 20000 13964 20052
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 17224 20000 17276 20052
rect 21916 20043 21968 20052
rect 21916 20009 21925 20043
rect 21925 20009 21959 20043
rect 21959 20009 21968 20043
rect 21916 20000 21968 20009
rect 23020 20000 23072 20052
rect 11428 19932 11480 19984
rect 15660 19932 15712 19984
rect 9496 19907 9548 19916
rect 9496 19873 9505 19907
rect 9505 19873 9539 19907
rect 9539 19873 9548 19907
rect 9496 19864 9548 19873
rect 14924 19864 14976 19916
rect 7932 19796 7984 19848
rect 11520 19796 11572 19848
rect 23112 19864 23164 19916
rect 28172 20000 28224 20052
rect 30380 20043 30432 20052
rect 30380 20009 30389 20043
rect 30389 20009 30423 20043
rect 30423 20009 30432 20043
rect 30380 20000 30432 20009
rect 33048 20000 33100 20052
rect 4620 19728 4672 19780
rect 6460 19771 6512 19780
rect 6460 19737 6469 19771
rect 6469 19737 6503 19771
rect 6503 19737 6512 19771
rect 6460 19728 6512 19737
rect 11152 19728 11204 19780
rect 14372 19728 14424 19780
rect 15016 19728 15068 19780
rect 17776 19796 17828 19848
rect 22560 19796 22612 19848
rect 22744 19839 22796 19848
rect 22744 19805 22753 19839
rect 22753 19805 22787 19839
rect 22787 19805 22796 19839
rect 22744 19796 22796 19805
rect 23296 19796 23348 19848
rect 25320 19796 25372 19848
rect 25872 19839 25924 19848
rect 25872 19805 25881 19839
rect 25881 19805 25915 19839
rect 25915 19805 25924 19839
rect 25872 19796 25924 19805
rect 28632 19864 28684 19916
rect 28908 19907 28960 19916
rect 28908 19873 28917 19907
rect 28917 19873 28951 19907
rect 28951 19873 28960 19907
rect 28908 19864 28960 19873
rect 30288 19839 30340 19848
rect 30288 19805 30297 19839
rect 30297 19805 30331 19839
rect 30331 19805 30340 19839
rect 30288 19796 30340 19805
rect 38292 19839 38344 19848
rect 38292 19805 38301 19839
rect 38301 19805 38335 19839
rect 38335 19805 38344 19839
rect 38292 19796 38344 19805
rect 28356 19771 28408 19780
rect 28356 19737 28365 19771
rect 28365 19737 28399 19771
rect 28399 19737 28408 19771
rect 28356 19728 28408 19737
rect 5540 19660 5592 19712
rect 5632 19660 5684 19712
rect 11796 19660 11848 19712
rect 22560 19703 22612 19712
rect 22560 19669 22569 19703
rect 22569 19669 22603 19703
rect 22603 19669 22612 19703
rect 22560 19660 22612 19669
rect 25412 19660 25464 19712
rect 26332 19703 26384 19712
rect 26332 19669 26341 19703
rect 26341 19669 26375 19703
rect 26375 19669 26384 19703
rect 26332 19660 26384 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3976 19499 4028 19508
rect 3976 19465 3985 19499
rect 3985 19465 4019 19499
rect 4019 19465 4028 19499
rect 3976 19456 4028 19465
rect 10784 19456 10836 19508
rect 11428 19388 11480 19440
rect 11796 19431 11848 19440
rect 11796 19397 11805 19431
rect 11805 19397 11839 19431
rect 11839 19397 11848 19431
rect 11796 19388 11848 19397
rect 13360 19388 13412 19440
rect 14096 19456 14148 19508
rect 19248 19456 19300 19508
rect 25320 19499 25372 19508
rect 25320 19465 25329 19499
rect 25329 19465 25363 19499
rect 25363 19465 25372 19499
rect 25320 19456 25372 19465
rect 17408 19388 17460 19440
rect 19340 19431 19392 19440
rect 19340 19397 19349 19431
rect 19349 19397 19383 19431
rect 19383 19397 19392 19431
rect 19340 19388 19392 19397
rect 27344 19431 27396 19440
rect 27344 19397 27353 19431
rect 27353 19397 27387 19431
rect 27387 19397 27396 19431
rect 27344 19388 27396 19397
rect 22560 19363 22612 19372
rect 22560 19329 22569 19363
rect 22569 19329 22603 19363
rect 22603 19329 22612 19363
rect 22560 19320 22612 19329
rect 25872 19320 25924 19372
rect 28448 19320 28500 19372
rect 28632 19320 28684 19372
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 2504 19295 2556 19304
rect 2504 19261 2513 19295
rect 2513 19261 2547 19295
rect 2547 19261 2556 19295
rect 2504 19252 2556 19261
rect 9312 19252 9364 19304
rect 12256 19295 12308 19304
rect 12256 19261 12265 19295
rect 12265 19261 12299 19295
rect 12299 19261 12308 19295
rect 12256 19252 12308 19261
rect 6736 19184 6788 19236
rect 12900 19252 12952 19304
rect 13912 19252 13964 19304
rect 16856 19295 16908 19304
rect 16856 19261 16865 19295
rect 16865 19261 16899 19295
rect 16899 19261 16908 19295
rect 16856 19252 16908 19261
rect 19432 19252 19484 19304
rect 20628 19295 20680 19304
rect 18144 19184 18196 19236
rect 8392 19116 8444 19168
rect 16672 19116 16724 19168
rect 19248 19116 19300 19168
rect 20628 19261 20637 19295
rect 20637 19261 20671 19295
rect 20671 19261 20680 19295
rect 20628 19252 20680 19261
rect 27252 19295 27304 19304
rect 27252 19261 27261 19295
rect 27261 19261 27295 19295
rect 27295 19261 27304 19295
rect 27252 19252 27304 19261
rect 27804 19227 27856 19236
rect 27804 19193 27813 19227
rect 27813 19193 27847 19227
rect 27847 19193 27856 19227
rect 27804 19184 27856 19193
rect 27896 19184 27948 19236
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 8300 18955 8352 18964
rect 2412 18751 2464 18760
rect 2412 18717 2421 18751
rect 2421 18717 2455 18751
rect 2455 18717 2464 18751
rect 2412 18708 2464 18717
rect 6092 18887 6144 18896
rect 6092 18853 6101 18887
rect 6101 18853 6135 18887
rect 6135 18853 6144 18887
rect 6092 18844 6144 18853
rect 4620 18776 4672 18828
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 9036 18912 9088 18964
rect 13360 18844 13412 18896
rect 13912 18776 13964 18828
rect 19340 18912 19392 18964
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 4896 18640 4948 18692
rect 6828 18683 6880 18692
rect 6828 18649 6837 18683
rect 6837 18649 6871 18683
rect 6871 18649 6880 18683
rect 6828 18640 6880 18649
rect 7564 18640 7616 18692
rect 10876 18640 10928 18692
rect 12348 18683 12400 18692
rect 12348 18649 12357 18683
rect 12357 18649 12391 18683
rect 12391 18649 12400 18683
rect 12348 18640 12400 18649
rect 15568 18640 15620 18692
rect 16856 18776 16908 18828
rect 19156 18776 19208 18828
rect 20168 18844 20220 18896
rect 24768 18844 24820 18896
rect 20628 18819 20680 18828
rect 20628 18785 20637 18819
rect 20637 18785 20671 18819
rect 20671 18785 20680 18819
rect 20628 18776 20680 18785
rect 19340 18708 19392 18760
rect 27344 18912 27396 18964
rect 27896 18912 27948 18964
rect 28356 18912 28408 18964
rect 30472 18912 30524 18964
rect 28448 18776 28500 18828
rect 27712 18751 27764 18760
rect 16488 18683 16540 18692
rect 11520 18572 11572 18624
rect 16488 18649 16497 18683
rect 16497 18649 16531 18683
rect 16531 18649 16540 18683
rect 16488 18640 16540 18649
rect 17040 18683 17092 18692
rect 17040 18649 17049 18683
rect 17049 18649 17083 18683
rect 17083 18649 17092 18683
rect 17040 18640 17092 18649
rect 15752 18572 15804 18624
rect 17960 18640 18012 18692
rect 19432 18640 19484 18692
rect 19984 18640 20036 18692
rect 25044 18640 25096 18692
rect 22652 18615 22704 18624
rect 22652 18581 22661 18615
rect 22661 18581 22695 18615
rect 22695 18581 22704 18615
rect 22652 18572 22704 18581
rect 24308 18572 24360 18624
rect 26056 18572 26108 18624
rect 27712 18717 27721 18751
rect 27721 18717 27755 18751
rect 27755 18717 27764 18751
rect 27712 18708 27764 18717
rect 28356 18751 28408 18760
rect 28356 18717 28365 18751
rect 28365 18717 28399 18751
rect 28399 18717 28408 18751
rect 28356 18708 28408 18717
rect 29460 18708 29512 18760
rect 29644 18708 29696 18760
rect 29828 18708 29880 18760
rect 38292 18751 38344 18760
rect 38292 18717 38301 18751
rect 38301 18717 38335 18751
rect 38335 18717 38344 18751
rect 38292 18708 38344 18717
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 3332 18368 3384 18420
rect 3884 18368 3936 18420
rect 6828 18368 6880 18420
rect 12348 18368 12400 18420
rect 20168 18368 20220 18420
rect 4068 18300 4120 18352
rect 4896 18300 4948 18352
rect 14924 18300 14976 18352
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 1584 18164 1636 18216
rect 2228 18164 2280 18216
rect 3792 18164 3844 18216
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 13176 18207 13228 18216
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 23848 18300 23900 18352
rect 16672 18232 16724 18284
rect 13176 18164 13228 18173
rect 9220 18096 9272 18148
rect 19156 18232 19208 18284
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 26240 18368 26292 18420
rect 26608 18368 26660 18420
rect 29644 18411 29696 18420
rect 29644 18377 29653 18411
rect 29653 18377 29687 18411
rect 29687 18377 29696 18411
rect 29644 18368 29696 18377
rect 24308 18343 24360 18352
rect 24308 18309 24317 18343
rect 24317 18309 24351 18343
rect 24351 18309 24360 18343
rect 24308 18300 24360 18309
rect 25504 18343 25556 18352
rect 25504 18309 25513 18343
rect 25513 18309 25547 18343
rect 25547 18309 25556 18343
rect 25504 18300 25556 18309
rect 26792 18232 26844 18284
rect 30288 18232 30340 18284
rect 2320 18028 2372 18080
rect 7288 18028 7340 18080
rect 14556 18028 14608 18080
rect 17224 18071 17276 18080
rect 17224 18037 17233 18071
rect 17233 18037 17267 18071
rect 17267 18037 17276 18071
rect 22560 18164 22612 18216
rect 24216 18207 24268 18216
rect 24216 18173 24225 18207
rect 24225 18173 24259 18207
rect 24259 18173 24268 18207
rect 24216 18164 24268 18173
rect 25412 18207 25464 18216
rect 25412 18173 25421 18207
rect 25421 18173 25455 18207
rect 25455 18173 25464 18207
rect 25412 18164 25464 18173
rect 30932 18207 30984 18216
rect 19340 18096 19392 18148
rect 20076 18096 20128 18148
rect 17224 18028 17276 18037
rect 20628 18028 20680 18080
rect 22468 18028 22520 18080
rect 30932 18173 30941 18207
rect 30941 18173 30975 18207
rect 30975 18173 30984 18207
rect 30932 18164 30984 18173
rect 31024 18096 31076 18148
rect 25044 18028 25096 18080
rect 29920 18028 29972 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 5080 17824 5132 17876
rect 10784 17824 10836 17876
rect 14924 17867 14976 17876
rect 14924 17833 14933 17867
rect 14933 17833 14967 17867
rect 14967 17833 14976 17867
rect 14924 17824 14976 17833
rect 18236 17824 18288 17876
rect 18880 17824 18932 17876
rect 22560 17824 22612 17876
rect 25504 17824 25556 17876
rect 29828 17824 29880 17876
rect 12440 17756 12492 17808
rect 4344 17731 4396 17740
rect 4344 17697 4353 17731
rect 4353 17697 4387 17731
rect 4387 17697 4396 17731
rect 4344 17688 4396 17697
rect 4620 17688 4672 17740
rect 5080 17688 5132 17740
rect 8944 17620 8996 17672
rect 14924 17688 14976 17740
rect 17224 17731 17276 17740
rect 15476 17620 15528 17672
rect 17224 17697 17233 17731
rect 17233 17697 17267 17731
rect 17267 17697 17276 17731
rect 17224 17688 17276 17697
rect 20812 17756 20864 17808
rect 22468 17688 22520 17740
rect 22652 17731 22704 17740
rect 22652 17697 22661 17731
rect 22661 17697 22695 17731
rect 22695 17697 22704 17731
rect 22652 17688 22704 17697
rect 26332 17756 26384 17808
rect 26424 17756 26476 17808
rect 26608 17688 26660 17740
rect 30932 17688 30984 17740
rect 17868 17620 17920 17672
rect 22008 17663 22060 17672
rect 22008 17629 22017 17663
rect 22017 17629 22051 17663
rect 22051 17629 22060 17663
rect 22008 17620 22060 17629
rect 25044 17663 25096 17672
rect 25044 17629 25053 17663
rect 25053 17629 25087 17663
rect 25087 17629 25096 17663
rect 25044 17620 25096 17629
rect 26332 17663 26384 17672
rect 6368 17595 6420 17604
rect 6368 17561 6377 17595
rect 6377 17561 6411 17595
rect 6411 17561 6420 17595
rect 6368 17552 6420 17561
rect 9404 17595 9456 17604
rect 9404 17561 9413 17595
rect 9413 17561 9447 17595
rect 9447 17561 9456 17595
rect 9404 17552 9456 17561
rect 18328 17595 18380 17604
rect 18328 17561 18337 17595
rect 18337 17561 18371 17595
rect 18371 17561 18380 17595
rect 18328 17552 18380 17561
rect 19340 17552 19392 17604
rect 20444 17595 20496 17604
rect 20444 17561 20453 17595
rect 20453 17561 20487 17595
rect 20487 17561 20496 17595
rect 20444 17552 20496 17561
rect 26332 17629 26341 17663
rect 26341 17629 26375 17663
rect 26375 17629 26384 17663
rect 26332 17620 26384 17629
rect 27896 17663 27948 17672
rect 27896 17629 27905 17663
rect 27905 17629 27939 17663
rect 27939 17629 27948 17663
rect 27896 17620 27948 17629
rect 29920 17663 29972 17672
rect 26240 17552 26292 17604
rect 27344 17552 27396 17604
rect 29920 17629 29929 17663
rect 29929 17629 29963 17663
rect 29963 17629 29972 17663
rect 29920 17620 29972 17629
rect 30564 17663 30616 17672
rect 30564 17629 30573 17663
rect 30573 17629 30607 17663
rect 30607 17629 30616 17663
rect 30564 17620 30616 17629
rect 30380 17552 30432 17604
rect 13636 17484 13688 17536
rect 15844 17527 15896 17536
rect 15844 17493 15853 17527
rect 15853 17493 15887 17527
rect 15887 17493 15896 17527
rect 15844 17484 15896 17493
rect 17960 17484 18012 17536
rect 20536 17484 20588 17536
rect 24216 17484 24268 17536
rect 29000 17527 29052 17536
rect 29000 17493 29009 17527
rect 29009 17493 29043 17527
rect 29043 17493 29052 17527
rect 29000 17484 29052 17493
rect 31024 17527 31076 17536
rect 31024 17493 31033 17527
rect 31033 17493 31067 17527
rect 31067 17493 31076 17527
rect 31024 17484 31076 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 9220 17280 9272 17332
rect 9312 17280 9364 17332
rect 7932 17212 7984 17264
rect 8668 17212 8720 17264
rect 13544 17255 13596 17264
rect 13544 17221 13553 17255
rect 13553 17221 13587 17255
rect 13587 17221 13596 17255
rect 13544 17212 13596 17221
rect 15844 17212 15896 17264
rect 18328 17280 18380 17332
rect 20444 17280 20496 17332
rect 17960 17212 18012 17264
rect 18972 17255 19024 17264
rect 18972 17221 18981 17255
rect 18981 17221 19015 17255
rect 19015 17221 19024 17255
rect 18972 17212 19024 17221
rect 25964 17255 26016 17264
rect 18420 17144 18472 17196
rect 25964 17221 25973 17255
rect 25973 17221 26007 17255
rect 26007 17221 26016 17255
rect 25964 17212 26016 17221
rect 26608 17212 26660 17264
rect 27896 17280 27948 17332
rect 30564 17280 30616 17332
rect 31024 17280 31076 17332
rect 31760 17212 31812 17264
rect 20628 17187 20680 17196
rect 4344 17076 4396 17128
rect 5172 17076 5224 17128
rect 8944 17076 8996 17128
rect 12900 17076 12952 17128
rect 13636 17076 13688 17128
rect 17592 17076 17644 17128
rect 20628 17153 20637 17187
rect 20637 17153 20671 17187
rect 20671 17153 20680 17187
rect 20628 17144 20680 17153
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 20996 17076 21048 17128
rect 27344 17144 27396 17196
rect 29000 17144 29052 17196
rect 30380 17144 30432 17196
rect 38292 17187 38344 17196
rect 38292 17153 38301 17187
rect 38301 17153 38335 17187
rect 38335 17153 38344 17187
rect 38292 17144 38344 17153
rect 14648 16940 14700 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 18512 17008 18564 17060
rect 26240 17076 26292 17128
rect 32404 17076 32456 17128
rect 24768 17008 24820 17060
rect 26516 17051 26568 17060
rect 26516 17017 26525 17051
rect 26525 17017 26559 17051
rect 26559 17017 26568 17051
rect 26516 17008 26568 17017
rect 22284 16940 22336 16992
rect 22468 16940 22520 16992
rect 35900 16940 35952 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 8392 16736 8444 16788
rect 8760 16736 8812 16788
rect 5172 16600 5224 16652
rect 11152 16600 11204 16652
rect 16488 16668 16540 16720
rect 16764 16668 16816 16720
rect 18972 16736 19024 16788
rect 20996 16779 21048 16788
rect 20996 16745 21005 16779
rect 21005 16745 21039 16779
rect 21039 16745 21048 16779
rect 20996 16736 21048 16745
rect 22284 16736 22336 16788
rect 23204 16736 23256 16788
rect 32404 16779 32456 16788
rect 32404 16745 32413 16779
rect 32413 16745 32447 16779
rect 32447 16745 32456 16779
rect 32404 16736 32456 16745
rect 21088 16668 21140 16720
rect 1768 16575 1820 16584
rect 1768 16541 1777 16575
rect 1777 16541 1811 16575
rect 1811 16541 1820 16575
rect 1768 16532 1820 16541
rect 8944 16532 8996 16584
rect 10324 16575 10376 16584
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 14832 16532 14884 16584
rect 15476 16600 15528 16652
rect 17500 16600 17552 16652
rect 18052 16532 18104 16584
rect 20996 16532 21048 16584
rect 25504 16532 25556 16584
rect 25872 16532 25924 16584
rect 27896 16600 27948 16652
rect 31024 16600 31076 16652
rect 1492 16396 1544 16448
rect 5448 16396 5500 16448
rect 13268 16464 13320 16516
rect 7564 16396 7616 16448
rect 15384 16439 15436 16448
rect 15384 16405 15393 16439
rect 15393 16405 15427 16439
rect 15427 16405 15436 16439
rect 15384 16396 15436 16405
rect 16396 16464 16448 16516
rect 23848 16464 23900 16516
rect 27344 16575 27396 16584
rect 27344 16541 27353 16575
rect 27353 16541 27387 16575
rect 27387 16541 27396 16575
rect 27344 16532 27396 16541
rect 30656 16575 30708 16584
rect 30656 16541 30665 16575
rect 30665 16541 30699 16575
rect 30699 16541 30708 16575
rect 30656 16532 30708 16541
rect 37096 16600 37148 16652
rect 19984 16396 20036 16448
rect 24768 16396 24820 16448
rect 26332 16396 26384 16448
rect 26608 16439 26660 16448
rect 26608 16405 26617 16439
rect 26617 16405 26651 16439
rect 26651 16405 26660 16439
rect 26608 16396 26660 16405
rect 31116 16439 31168 16448
rect 31116 16405 31125 16439
rect 31125 16405 31159 16439
rect 31159 16405 31168 16439
rect 31116 16396 31168 16405
rect 33600 16439 33652 16448
rect 33600 16405 33609 16439
rect 33609 16405 33643 16439
rect 33643 16405 33652 16439
rect 33600 16396 33652 16405
rect 35900 16396 35952 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 3976 16192 4028 16244
rect 15384 16192 15436 16244
rect 20996 16235 21048 16244
rect 11336 16124 11388 16176
rect 13268 16124 13320 16176
rect 17224 16124 17276 16176
rect 20996 16201 21005 16235
rect 21005 16201 21039 16235
rect 21039 16201 21048 16235
rect 20996 16192 21048 16201
rect 23112 16192 23164 16244
rect 24216 16192 24268 16244
rect 25504 16235 25556 16244
rect 25504 16201 25513 16235
rect 25513 16201 25547 16235
rect 25547 16201 25556 16235
rect 25504 16192 25556 16201
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 8944 16099 8996 16108
rect 8944 16065 8953 16099
rect 8953 16065 8987 16099
rect 8987 16065 8996 16099
rect 8944 16056 8996 16065
rect 14280 16056 14332 16108
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 20168 16099 20220 16108
rect 19248 16056 19300 16065
rect 20168 16065 20177 16099
rect 20177 16065 20211 16099
rect 20211 16065 20220 16099
rect 20168 16056 20220 16065
rect 20904 16056 20956 16108
rect 24768 16056 24820 16108
rect 3608 16031 3660 16040
rect 3608 15997 3617 16031
rect 3617 15997 3651 16031
rect 3651 15997 3660 16031
rect 3608 15988 3660 15997
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 10968 15988 11020 16040
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 14188 15988 14240 16040
rect 15108 15988 15160 16040
rect 17408 16031 17460 16040
rect 17408 15997 17417 16031
rect 17417 15997 17451 16031
rect 17451 15997 17460 16031
rect 17408 15988 17460 15997
rect 18696 15988 18748 16040
rect 22192 15988 22244 16040
rect 22744 16031 22796 16040
rect 22744 15997 22753 16031
rect 22753 15997 22787 16031
rect 22787 15997 22796 16031
rect 22744 15988 22796 15997
rect 23940 16031 23992 16040
rect 10600 15852 10652 15904
rect 18512 15920 18564 15972
rect 20444 15920 20496 15972
rect 23940 15997 23949 16031
rect 23949 15997 23983 16031
rect 23983 15997 23992 16031
rect 23940 15988 23992 15997
rect 24584 15988 24636 16040
rect 28448 16031 28500 16040
rect 28448 15997 28457 16031
rect 28457 15997 28491 16031
rect 28491 15997 28500 16031
rect 28448 15988 28500 15997
rect 28540 15988 28592 16040
rect 29552 16031 29604 16040
rect 29552 15997 29561 16031
rect 29561 15997 29595 16031
rect 29595 15997 29604 16031
rect 29552 15988 29604 15997
rect 29828 15988 29880 16040
rect 30104 15920 30156 15972
rect 28356 15852 28408 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3608 15648 3660 15700
rect 13176 15648 13228 15700
rect 14280 15648 14332 15700
rect 16396 15691 16448 15700
rect 16396 15657 16405 15691
rect 16405 15657 16439 15691
rect 16439 15657 16448 15691
rect 16396 15648 16448 15657
rect 17224 15691 17276 15700
rect 17224 15657 17233 15691
rect 17233 15657 17267 15691
rect 17267 15657 17276 15691
rect 17224 15648 17276 15657
rect 17592 15648 17644 15700
rect 22744 15691 22796 15700
rect 4068 15623 4120 15632
rect 4068 15589 4077 15623
rect 4077 15589 4111 15623
rect 4111 15589 4120 15623
rect 4068 15580 4120 15589
rect 10324 15512 10376 15564
rect 10968 15555 11020 15564
rect 10968 15521 10977 15555
rect 10977 15521 11011 15555
rect 11011 15521 11020 15555
rect 10968 15512 11020 15521
rect 4068 15444 4120 15496
rect 14832 15444 14884 15496
rect 15936 15487 15988 15496
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 18052 15487 18104 15496
rect 18052 15453 18061 15487
rect 18061 15453 18095 15487
rect 18095 15453 18104 15487
rect 18052 15444 18104 15453
rect 12808 15376 12860 15428
rect 12992 15419 13044 15428
rect 12992 15385 13001 15419
rect 13001 15385 13035 15419
rect 13035 15385 13044 15419
rect 18696 15555 18748 15564
rect 18696 15521 18705 15555
rect 18705 15521 18739 15555
rect 18739 15521 18748 15555
rect 18696 15512 18748 15521
rect 20260 15512 20312 15564
rect 22744 15657 22753 15691
rect 22753 15657 22787 15691
rect 22787 15657 22796 15691
rect 22744 15648 22796 15657
rect 23940 15691 23992 15700
rect 23940 15657 23949 15691
rect 23949 15657 23983 15691
rect 23983 15657 23992 15691
rect 23940 15648 23992 15657
rect 25228 15691 25280 15700
rect 25228 15657 25237 15691
rect 25237 15657 25271 15691
rect 25271 15657 25280 15691
rect 25228 15648 25280 15657
rect 28540 15648 28592 15700
rect 29828 15691 29880 15700
rect 29828 15657 29837 15691
rect 29837 15657 29871 15691
rect 29871 15657 29880 15691
rect 29828 15648 29880 15657
rect 30656 15648 30708 15700
rect 25412 15580 25464 15632
rect 24584 15555 24636 15564
rect 21364 15444 21416 15496
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 26424 15555 26476 15564
rect 26424 15521 26433 15555
rect 26433 15521 26467 15555
rect 26467 15521 26476 15555
rect 26424 15512 26476 15521
rect 28448 15555 28500 15564
rect 28448 15521 28457 15555
rect 28457 15521 28491 15555
rect 28491 15521 28500 15555
rect 28448 15512 28500 15521
rect 22652 15487 22704 15496
rect 22652 15453 22661 15487
rect 22661 15453 22695 15487
rect 22695 15453 22704 15487
rect 22652 15444 22704 15453
rect 23848 15487 23900 15496
rect 23848 15453 23857 15487
rect 23857 15453 23891 15487
rect 23891 15453 23900 15487
rect 23848 15444 23900 15453
rect 25872 15444 25924 15496
rect 26608 15487 26660 15496
rect 26608 15453 26617 15487
rect 26617 15453 26651 15487
rect 26651 15453 26660 15487
rect 26608 15444 26660 15453
rect 27988 15487 28040 15496
rect 27988 15453 27997 15487
rect 27997 15453 28031 15487
rect 28031 15453 28040 15487
rect 27988 15444 28040 15453
rect 30564 15487 30616 15496
rect 30564 15453 30573 15487
rect 30573 15453 30607 15487
rect 30607 15453 30616 15487
rect 30564 15444 30616 15453
rect 31116 15580 31168 15632
rect 32404 15444 32456 15496
rect 12992 15376 13044 15385
rect 15384 15308 15436 15360
rect 21272 15376 21324 15428
rect 22928 15376 22980 15428
rect 28540 15376 28592 15428
rect 20996 15308 21048 15360
rect 28080 15308 28132 15360
rect 38200 15351 38252 15360
rect 38200 15317 38209 15351
rect 38209 15317 38243 15351
rect 38243 15317 38252 15351
rect 38200 15308 38252 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 10508 15104 10560 15156
rect 4896 15036 4948 15088
rect 5080 15079 5132 15088
rect 5080 15045 5089 15079
rect 5089 15045 5123 15079
rect 5123 15045 5132 15079
rect 5080 15036 5132 15045
rect 12164 15036 12216 15088
rect 1584 14968 1636 15020
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 4068 14968 4120 15020
rect 16580 15036 16632 15088
rect 17500 15104 17552 15156
rect 20168 15104 20220 15156
rect 20996 15147 21048 15156
rect 20996 15113 21005 15147
rect 21005 15113 21039 15147
rect 21039 15113 21048 15147
rect 20996 15104 21048 15113
rect 25228 15104 25280 15156
rect 25872 15147 25924 15156
rect 25872 15113 25881 15147
rect 25881 15113 25915 15147
rect 25915 15113 25924 15147
rect 25872 15104 25924 15113
rect 26608 15104 26660 15156
rect 27988 15104 28040 15156
rect 30564 15104 30616 15156
rect 18052 15036 18104 15088
rect 22008 15036 22060 15088
rect 24400 15036 24452 15088
rect 24768 15036 24820 15088
rect 20076 15011 20128 15020
rect 2136 14943 2188 14952
rect 2136 14909 2145 14943
rect 2145 14909 2179 14943
rect 2179 14909 2188 14943
rect 2136 14900 2188 14909
rect 5172 14900 5224 14952
rect 7748 14943 7800 14952
rect 7748 14909 7757 14943
rect 7757 14909 7791 14943
rect 7791 14909 7800 14943
rect 9496 14943 9548 14952
rect 7748 14900 7800 14909
rect 9496 14909 9505 14943
rect 9505 14909 9539 14943
rect 9539 14909 9548 14943
rect 9496 14900 9548 14909
rect 12900 14900 12952 14952
rect 14004 14943 14056 14952
rect 14004 14909 14013 14943
rect 14013 14909 14047 14943
rect 14047 14909 14056 14943
rect 14004 14900 14056 14909
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 12624 14832 12676 14884
rect 9680 14764 9732 14816
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 17960 14900 18012 14952
rect 21180 14968 21232 15020
rect 25596 14968 25648 15020
rect 27068 14968 27120 15020
rect 28540 15011 28592 15020
rect 28540 14977 28549 15011
rect 28549 14977 28583 15011
rect 28583 14977 28592 15011
rect 28540 14968 28592 14977
rect 15108 14832 15160 14884
rect 24676 14900 24728 14952
rect 21548 14832 21600 14884
rect 24584 14832 24636 14884
rect 26332 14900 26384 14952
rect 27528 14832 27580 14884
rect 22836 14764 22888 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4712 14560 4764 14612
rect 7748 14560 7800 14612
rect 11152 14603 11204 14612
rect 11152 14569 11161 14603
rect 11161 14569 11195 14603
rect 11195 14569 11204 14603
rect 11152 14560 11204 14569
rect 11336 14560 11388 14612
rect 21364 14603 21416 14612
rect 21364 14569 21373 14603
rect 21373 14569 21407 14603
rect 21407 14569 21416 14603
rect 21364 14560 21416 14569
rect 4804 14492 4856 14544
rect 2504 14424 2556 14476
rect 5172 14424 5224 14476
rect 3332 14356 3384 14408
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 8944 14424 8996 14476
rect 9404 14467 9456 14476
rect 9404 14433 9413 14467
rect 9413 14433 9447 14467
rect 9447 14433 9456 14467
rect 9404 14424 9456 14433
rect 10968 14492 11020 14544
rect 16764 14492 16816 14544
rect 25596 14535 25648 14544
rect 15016 14424 15068 14476
rect 15476 14424 15528 14476
rect 16948 14424 17000 14476
rect 20904 14424 20956 14476
rect 11612 14399 11664 14408
rect 11612 14365 11621 14399
rect 11621 14365 11655 14399
rect 11655 14365 11664 14399
rect 11612 14356 11664 14365
rect 2136 14220 2188 14272
rect 5264 14288 5316 14340
rect 9680 14331 9732 14340
rect 9680 14297 9689 14331
rect 9689 14297 9723 14331
rect 9723 14297 9732 14331
rect 9680 14288 9732 14297
rect 11428 14288 11480 14340
rect 5540 14220 5592 14272
rect 9220 14220 9272 14272
rect 10324 14220 10376 14272
rect 14464 14356 14516 14408
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 16304 14399 16356 14408
rect 13820 14288 13872 14340
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 18144 14356 18196 14408
rect 20812 14356 20864 14408
rect 25596 14501 25605 14535
rect 25605 14501 25639 14535
rect 25639 14501 25648 14535
rect 25596 14492 25648 14501
rect 26332 14603 26384 14612
rect 26332 14569 26341 14603
rect 26341 14569 26375 14603
rect 26375 14569 26384 14603
rect 28632 14603 28684 14612
rect 26332 14560 26384 14569
rect 28632 14569 28641 14603
rect 28641 14569 28675 14603
rect 28675 14569 28684 14603
rect 28632 14560 28684 14569
rect 23848 14424 23900 14476
rect 22836 14399 22888 14408
rect 22836 14365 22845 14399
rect 22845 14365 22879 14399
rect 22879 14365 22888 14399
rect 22836 14356 22888 14365
rect 24584 14356 24636 14408
rect 29920 14424 29972 14476
rect 27712 14356 27764 14408
rect 28264 14356 28316 14408
rect 16672 14288 16724 14340
rect 14832 14220 14884 14272
rect 18144 14220 18196 14272
rect 18880 14220 18932 14272
rect 20536 14288 20588 14340
rect 26332 14288 26384 14340
rect 26792 14288 26844 14340
rect 28448 14220 28500 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 9496 14016 9548 14068
rect 20536 14016 20588 14068
rect 22744 14016 22796 14068
rect 4896 13948 4948 14000
rect 1584 13880 1636 13932
rect 2504 13880 2556 13932
rect 4068 13812 4120 13864
rect 9496 13880 9548 13932
rect 10324 13948 10376 14000
rect 16764 13948 16816 14000
rect 17224 13991 17276 14000
rect 17224 13957 17233 13991
rect 17233 13957 17267 13991
rect 17267 13957 17276 13991
rect 17224 13948 17276 13957
rect 18880 13991 18932 14000
rect 18880 13957 18889 13991
rect 18889 13957 18923 13991
rect 18923 13957 18932 13991
rect 18880 13948 18932 13957
rect 18972 13991 19024 14000
rect 18972 13957 18981 13991
rect 18981 13957 19015 13991
rect 19015 13957 19024 13991
rect 18972 13948 19024 13957
rect 21272 13948 21324 14000
rect 23480 13991 23532 14000
rect 23480 13957 23489 13991
rect 23489 13957 23523 13991
rect 23523 13957 23532 13991
rect 23480 13948 23532 13957
rect 24952 14016 25004 14068
rect 28264 14059 28316 14068
rect 15108 13880 15160 13932
rect 15752 13880 15804 13932
rect 16304 13880 16356 13932
rect 20904 13880 20956 13932
rect 23020 13880 23072 13932
rect 14004 13812 14056 13864
rect 14740 13812 14792 13864
rect 16488 13812 16540 13864
rect 17592 13855 17644 13864
rect 17592 13821 17601 13855
rect 17601 13821 17635 13855
rect 17635 13821 17644 13855
rect 17592 13812 17644 13821
rect 18236 13812 18288 13864
rect 19340 13855 19392 13864
rect 19340 13821 19349 13855
rect 19349 13821 19383 13855
rect 19383 13821 19392 13855
rect 19340 13812 19392 13821
rect 19984 13855 20036 13864
rect 19984 13821 19993 13855
rect 19993 13821 20027 13855
rect 20027 13821 20036 13855
rect 19984 13812 20036 13821
rect 22192 13855 22244 13864
rect 22192 13821 22201 13855
rect 22201 13821 22235 13855
rect 22235 13821 22244 13855
rect 22192 13812 22244 13821
rect 23388 13855 23440 13864
rect 23388 13821 23397 13855
rect 23397 13821 23431 13855
rect 23431 13821 23440 13855
rect 23388 13812 23440 13821
rect 24676 13923 24728 13932
rect 24676 13889 24685 13923
rect 24685 13889 24719 13923
rect 24719 13889 24728 13923
rect 24676 13880 24728 13889
rect 26332 13880 26384 13932
rect 28264 14025 28273 14059
rect 28273 14025 28307 14059
rect 28307 14025 28316 14059
rect 28264 14016 28316 14025
rect 37096 14016 37148 14068
rect 28448 13923 28500 13932
rect 28448 13889 28457 13923
rect 28457 13889 28491 13923
rect 28491 13889 28500 13923
rect 28448 13880 28500 13889
rect 38292 13923 38344 13932
rect 38292 13889 38301 13923
rect 38301 13889 38335 13923
rect 38335 13889 38344 13923
rect 38292 13880 38344 13889
rect 26976 13812 27028 13864
rect 23848 13744 23900 13796
rect 27160 13719 27212 13728
rect 27160 13685 27169 13719
rect 27169 13685 27203 13719
rect 27203 13685 27212 13719
rect 27160 13676 27212 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 11520 13515 11572 13524
rect 11520 13481 11529 13515
rect 11529 13481 11563 13515
rect 11563 13481 11572 13515
rect 11520 13472 11572 13481
rect 12808 13472 12860 13524
rect 17224 13472 17276 13524
rect 17960 13515 18012 13524
rect 17960 13481 17969 13515
rect 17969 13481 18003 13515
rect 18003 13481 18012 13515
rect 17960 13472 18012 13481
rect 23480 13472 23532 13524
rect 29920 13515 29972 13524
rect 29920 13481 29929 13515
rect 29929 13481 29963 13515
rect 29963 13481 29972 13515
rect 29920 13472 29972 13481
rect 14004 13404 14056 13456
rect 27804 13404 27856 13456
rect 30840 13447 30892 13456
rect 9404 13336 9456 13388
rect 9772 13379 9824 13388
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 15568 13336 15620 13388
rect 19984 13336 20036 13388
rect 23388 13379 23440 13388
rect 23388 13345 23397 13379
rect 23397 13345 23431 13379
rect 23431 13345 23440 13379
rect 23388 13336 23440 13345
rect 27160 13336 27212 13388
rect 2688 13268 2740 13320
rect 13452 13268 13504 13320
rect 15016 13311 15068 13320
rect 15016 13277 15025 13311
rect 15025 13277 15059 13311
rect 15059 13277 15068 13311
rect 15016 13268 15068 13277
rect 15660 13268 15712 13320
rect 18144 13311 18196 13320
rect 18144 13277 18153 13311
rect 18153 13277 18187 13311
rect 18187 13277 18196 13311
rect 18144 13268 18196 13277
rect 21732 13311 21784 13320
rect 10508 13200 10560 13252
rect 11428 13200 11480 13252
rect 14464 13200 14516 13252
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 24952 13311 25004 13320
rect 24952 13277 24961 13311
rect 24961 13277 24995 13311
rect 24995 13277 25004 13311
rect 24952 13268 25004 13277
rect 26240 13268 26292 13320
rect 26608 13268 26660 13320
rect 30840 13413 30849 13447
rect 30849 13413 30883 13447
rect 30883 13413 30892 13447
rect 30840 13404 30892 13413
rect 30472 13379 30524 13388
rect 30472 13345 30481 13379
rect 30481 13345 30515 13379
rect 30515 13345 30524 13379
rect 30472 13336 30524 13345
rect 36912 13336 36964 13388
rect 23112 13200 23164 13252
rect 1768 13175 1820 13184
rect 1768 13141 1777 13175
rect 1777 13141 1811 13175
rect 1811 13141 1820 13175
rect 1768 13132 1820 13141
rect 13360 13132 13412 13184
rect 14556 13132 14608 13184
rect 15200 13132 15252 13184
rect 20812 13132 20864 13184
rect 20904 13132 20956 13184
rect 28080 13132 28132 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 7564 12928 7616 12980
rect 12348 12928 12400 12980
rect 18972 12928 19024 12980
rect 3240 12860 3292 12912
rect 10968 12860 11020 12912
rect 13360 12903 13412 12912
rect 13360 12869 13369 12903
rect 13369 12869 13403 12903
rect 13403 12869 13412 12903
rect 13360 12860 13412 12869
rect 14740 12860 14792 12912
rect 16028 12903 16080 12912
rect 16028 12869 16037 12903
rect 16037 12869 16071 12903
rect 16071 12869 16080 12903
rect 16028 12860 16080 12869
rect 18604 12860 18656 12912
rect 20904 12903 20956 12912
rect 20904 12869 20913 12903
rect 20913 12869 20947 12903
rect 20947 12869 20956 12903
rect 20904 12860 20956 12869
rect 30840 12928 30892 12980
rect 24860 12860 24912 12912
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 11612 12792 11664 12844
rect 15292 12792 15344 12844
rect 15752 12835 15804 12844
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 15752 12792 15804 12801
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 23204 12835 23256 12844
rect 23204 12801 23213 12835
rect 23213 12801 23247 12835
rect 23247 12801 23256 12835
rect 23204 12792 23256 12801
rect 24400 12835 24452 12844
rect 24400 12801 24409 12835
rect 24409 12801 24443 12835
rect 24443 12801 24452 12835
rect 24400 12792 24452 12801
rect 6276 12724 6328 12776
rect 6828 12724 6880 12776
rect 8576 12588 8628 12640
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 12900 12724 12952 12776
rect 13452 12724 13504 12776
rect 14556 12724 14608 12776
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 17592 12767 17644 12776
rect 17592 12733 17601 12767
rect 17601 12733 17635 12767
rect 17635 12733 17644 12767
rect 17592 12724 17644 12733
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 21180 12767 21232 12776
rect 21180 12733 21189 12767
rect 21189 12733 21223 12767
rect 21223 12733 21232 12767
rect 21180 12724 21232 12733
rect 22376 12767 22428 12776
rect 22376 12733 22385 12767
rect 22385 12733 22419 12767
rect 22419 12733 22428 12767
rect 22376 12724 22428 12733
rect 16028 12656 16080 12708
rect 16948 12656 17000 12708
rect 23848 12656 23900 12708
rect 25780 12792 25832 12844
rect 26332 12835 26384 12844
rect 26332 12801 26341 12835
rect 26341 12801 26375 12835
rect 26375 12801 26384 12835
rect 26332 12792 26384 12801
rect 26792 12792 26844 12844
rect 27804 12835 27856 12844
rect 27804 12801 27813 12835
rect 27813 12801 27847 12835
rect 27847 12801 27856 12835
rect 27804 12792 27856 12801
rect 28080 12724 28132 12776
rect 14648 12588 14700 12640
rect 24952 12588 25004 12640
rect 27252 12631 27304 12640
rect 27252 12597 27261 12631
rect 27261 12597 27295 12631
rect 27295 12597 27304 12631
rect 27252 12588 27304 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3240 12427 3292 12436
rect 3240 12393 3249 12427
rect 3249 12393 3283 12427
rect 3283 12393 3292 12427
rect 3240 12384 3292 12393
rect 12164 12384 12216 12436
rect 16212 12384 16264 12436
rect 16580 12427 16632 12436
rect 16580 12393 16589 12427
rect 16589 12393 16623 12427
rect 16623 12393 16632 12427
rect 16580 12384 16632 12393
rect 18880 12384 18932 12436
rect 20812 12427 20864 12436
rect 20812 12393 20821 12427
rect 20821 12393 20855 12427
rect 20855 12393 20864 12427
rect 20812 12384 20864 12393
rect 21732 12384 21784 12436
rect 12624 12316 12676 12368
rect 6368 12291 6420 12300
rect 6368 12257 6377 12291
rect 6377 12257 6411 12291
rect 6411 12257 6420 12291
rect 6368 12248 6420 12257
rect 13636 12248 13688 12300
rect 15292 12248 15344 12300
rect 3332 12180 3384 12232
rect 5632 12180 5684 12232
rect 7932 12180 7984 12232
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 13452 12180 13504 12232
rect 13820 12180 13872 12232
rect 9312 12112 9364 12164
rect 14556 12155 14608 12164
rect 14556 12121 14565 12155
rect 14565 12121 14599 12155
rect 14599 12121 14608 12155
rect 14556 12112 14608 12121
rect 15200 12112 15252 12164
rect 7840 12087 7892 12096
rect 7840 12053 7849 12087
rect 7849 12053 7883 12087
rect 7883 12053 7892 12087
rect 7840 12044 7892 12053
rect 12808 12044 12860 12096
rect 14924 12044 14976 12096
rect 15292 12044 15344 12096
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 16488 12223 16540 12232
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 16488 12180 16540 12189
rect 17592 12316 17644 12368
rect 27344 12316 27396 12368
rect 18420 12223 18472 12232
rect 18420 12189 18429 12223
rect 18429 12189 18463 12223
rect 18463 12189 18472 12223
rect 18420 12180 18472 12189
rect 20444 12180 20496 12232
rect 21364 12223 21416 12232
rect 21364 12189 21373 12223
rect 21373 12189 21407 12223
rect 21407 12189 21416 12223
rect 21364 12180 21416 12189
rect 21640 12112 21692 12164
rect 24400 12180 24452 12232
rect 26056 12180 26108 12232
rect 30840 12180 30892 12232
rect 18144 12044 18196 12096
rect 22376 12044 22428 12096
rect 23204 12044 23256 12096
rect 23572 12044 23624 12096
rect 26148 12044 26200 12096
rect 32496 12044 32548 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 5540 11840 5592 11892
rect 5816 11840 5868 11892
rect 6736 11772 6788 11824
rect 10692 11840 10744 11892
rect 12900 11840 12952 11892
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 2504 11704 2556 11756
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 6828 11704 6880 11756
rect 6920 11704 6972 11756
rect 14464 11772 14516 11824
rect 7380 11636 7432 11688
rect 9588 11636 9640 11688
rect 13820 11704 13872 11756
rect 15016 11704 15068 11756
rect 15660 11704 15712 11756
rect 16488 11772 16540 11824
rect 18144 11840 18196 11892
rect 18420 11840 18472 11892
rect 27068 11840 27120 11892
rect 28080 11840 28132 11892
rect 32404 11840 32456 11892
rect 18236 11772 18288 11824
rect 18972 11815 19024 11824
rect 18972 11781 18981 11815
rect 18981 11781 19015 11815
rect 19015 11781 19024 11815
rect 18972 11772 19024 11781
rect 19984 11772 20036 11824
rect 25964 11772 26016 11824
rect 12532 11636 12584 11688
rect 17592 11704 17644 11756
rect 20260 11704 20312 11756
rect 23204 11747 23256 11756
rect 23204 11713 23213 11747
rect 23213 11713 23247 11747
rect 23247 11713 23256 11747
rect 23204 11704 23256 11713
rect 17500 11636 17552 11688
rect 17868 11636 17920 11688
rect 6368 11500 6420 11552
rect 6828 11500 6880 11552
rect 11612 11500 11664 11552
rect 11796 11543 11848 11552
rect 11796 11509 11805 11543
rect 11805 11509 11839 11543
rect 11839 11509 11848 11543
rect 11796 11500 11848 11509
rect 14556 11568 14608 11620
rect 21364 11636 21416 11688
rect 23388 11679 23440 11688
rect 23388 11645 23397 11679
rect 23397 11645 23431 11679
rect 23431 11645 23440 11679
rect 23388 11636 23440 11645
rect 25780 11679 25832 11688
rect 18972 11568 19024 11620
rect 15292 11500 15344 11552
rect 15384 11500 15436 11552
rect 16028 11500 16080 11552
rect 22652 11500 22704 11552
rect 23020 11568 23072 11620
rect 25228 11568 25280 11620
rect 25780 11645 25789 11679
rect 25789 11645 25823 11679
rect 25823 11645 25832 11679
rect 27712 11772 27764 11824
rect 27252 11704 27304 11756
rect 32496 11747 32548 11756
rect 32496 11713 32505 11747
rect 32505 11713 32539 11747
rect 32539 11713 32548 11747
rect 32496 11704 32548 11713
rect 38292 11747 38344 11756
rect 38292 11713 38301 11747
rect 38301 11713 38335 11747
rect 38335 11713 38344 11747
rect 38292 11704 38344 11713
rect 27160 11679 27212 11688
rect 25780 11636 25832 11645
rect 27160 11645 27169 11679
rect 27169 11645 27203 11679
rect 27203 11645 27212 11679
rect 27160 11636 27212 11645
rect 31760 11636 31812 11688
rect 25872 11568 25924 11620
rect 25044 11500 25096 11552
rect 34060 11500 34112 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 4068 11296 4120 11348
rect 9220 11228 9272 11280
rect 11612 11228 11664 11280
rect 14096 11228 14148 11280
rect 15108 11271 15160 11280
rect 15108 11237 15117 11271
rect 15117 11237 15151 11271
rect 15151 11237 15160 11271
rect 15108 11228 15160 11237
rect 1676 11160 1728 11212
rect 3976 11160 4028 11212
rect 5632 11160 5684 11212
rect 13728 11160 13780 11212
rect 18420 11296 18472 11348
rect 18604 11339 18656 11348
rect 18604 11305 18613 11339
rect 18613 11305 18647 11339
rect 18647 11305 18656 11339
rect 18604 11296 18656 11305
rect 23388 11339 23440 11348
rect 23388 11305 23397 11339
rect 23397 11305 23431 11339
rect 23431 11305 23440 11339
rect 23388 11296 23440 11305
rect 25228 11339 25280 11348
rect 25228 11305 25237 11339
rect 25237 11305 25271 11339
rect 25271 11305 25280 11339
rect 25228 11296 25280 11305
rect 25964 11339 26016 11348
rect 25964 11305 25973 11339
rect 25973 11305 26007 11339
rect 26007 11305 26016 11339
rect 25964 11296 26016 11305
rect 27528 11296 27580 11348
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 9772 11092 9824 11144
rect 11796 11092 11848 11144
rect 16672 11160 16724 11212
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 17684 11160 17736 11212
rect 25780 11228 25832 11280
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15660 11135 15712 11144
rect 15016 11092 15068 11101
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 15844 11092 15896 11144
rect 16488 11092 16540 11144
rect 24952 11160 25004 11212
rect 26976 11160 27028 11212
rect 19432 11092 19484 11144
rect 21640 11135 21692 11144
rect 21640 11101 21649 11135
rect 21649 11101 21683 11135
rect 21683 11101 21692 11135
rect 21640 11092 21692 11101
rect 22652 11092 22704 11144
rect 23572 11135 23624 11144
rect 5540 11024 5592 11076
rect 5724 11024 5776 11076
rect 12992 11024 13044 11076
rect 17592 11067 17644 11076
rect 17592 11033 17601 11067
rect 17601 11033 17635 11067
rect 17635 11033 17644 11067
rect 17592 11024 17644 11033
rect 17868 11024 17920 11076
rect 21180 11067 21232 11076
rect 11520 10956 11572 11008
rect 19340 10956 19392 11008
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 26148 11135 26200 11144
rect 24768 11024 24820 11076
rect 26148 11101 26157 11135
rect 26157 11101 26191 11135
rect 26191 11101 26200 11135
rect 26148 11092 26200 11101
rect 29736 11092 29788 11144
rect 26700 11024 26752 11076
rect 22836 10999 22888 11008
rect 22836 10965 22845 10999
rect 22845 10965 22879 10999
rect 22879 10965 22888 10999
rect 22836 10956 22888 10965
rect 31392 10999 31444 11008
rect 31392 10965 31401 10999
rect 31401 10965 31435 10999
rect 31435 10965 31444 10999
rect 31392 10956 31444 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 8760 10795 8812 10804
rect 8760 10761 8769 10795
rect 8769 10761 8803 10795
rect 8803 10761 8812 10795
rect 8760 10752 8812 10761
rect 9404 10752 9456 10804
rect 15016 10752 15068 10804
rect 17684 10752 17736 10804
rect 18236 10752 18288 10804
rect 36912 10752 36964 10804
rect 7564 10684 7616 10736
rect 14004 10684 14056 10736
rect 16212 10684 16264 10736
rect 16488 10684 16540 10736
rect 19340 10727 19392 10736
rect 19340 10693 19349 10727
rect 19349 10693 19383 10727
rect 19383 10693 19392 10727
rect 19340 10684 19392 10693
rect 20260 10684 20312 10736
rect 4620 10616 4672 10668
rect 5632 10616 5684 10668
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 15752 10616 15804 10668
rect 17500 10616 17552 10668
rect 22836 10616 22888 10668
rect 26056 10684 26108 10736
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 11428 10548 11480 10600
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 14832 10548 14884 10600
rect 16580 10480 16632 10532
rect 17408 10480 17460 10532
rect 22744 10548 22796 10600
rect 24768 10616 24820 10668
rect 24952 10548 25004 10600
rect 25688 10548 25740 10600
rect 27620 10616 27672 10668
rect 38292 10659 38344 10668
rect 38292 10625 38301 10659
rect 38301 10625 38335 10659
rect 38335 10625 38344 10659
rect 38292 10616 38344 10625
rect 32312 10548 32364 10600
rect 25872 10480 25924 10532
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 9680 10412 9732 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 23572 10455 23624 10464
rect 23572 10421 23581 10455
rect 23581 10421 23615 10455
rect 23615 10421 23624 10455
rect 23572 10412 23624 10421
rect 24032 10455 24084 10464
rect 24032 10421 24041 10455
rect 24041 10421 24075 10455
rect 24075 10421 24084 10455
rect 24032 10412 24084 10421
rect 24860 10412 24912 10464
rect 25320 10455 25372 10464
rect 25320 10421 25329 10455
rect 25329 10421 25363 10455
rect 25363 10421 25372 10455
rect 25320 10412 25372 10421
rect 33140 10412 33192 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 3884 10208 3936 10260
rect 4988 10140 5040 10192
rect 1584 10115 1636 10124
rect 1584 10081 1593 10115
rect 1593 10081 1627 10115
rect 1627 10081 1636 10115
rect 1584 10072 1636 10081
rect 2504 10072 2556 10124
rect 8576 10208 8628 10260
rect 15476 10208 15528 10260
rect 17592 10208 17644 10260
rect 19432 10208 19484 10260
rect 23112 10251 23164 10260
rect 23112 10217 23121 10251
rect 23121 10217 23155 10251
rect 23155 10217 23164 10251
rect 23112 10208 23164 10217
rect 11520 10140 11572 10192
rect 3148 9936 3200 9988
rect 12348 10072 12400 10124
rect 15016 10072 15068 10124
rect 3332 10004 3384 10056
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 9772 10004 9824 10056
rect 11428 10004 11480 10056
rect 17960 10047 18012 10056
rect 5632 9936 5684 9988
rect 6276 9936 6328 9988
rect 10140 9979 10192 9988
rect 10140 9945 10149 9979
rect 10149 9945 10183 9979
rect 10183 9945 10192 9979
rect 10140 9936 10192 9945
rect 13268 9936 13320 9988
rect 16212 9936 16264 9988
rect 17960 10013 17969 10047
rect 17969 10013 18003 10047
rect 18003 10013 18012 10047
rect 17960 10004 18012 10013
rect 20076 10115 20128 10124
rect 20076 10081 20085 10115
rect 20085 10081 20119 10115
rect 20119 10081 20128 10115
rect 20076 10072 20128 10081
rect 20444 10072 20496 10124
rect 24860 10115 24912 10124
rect 24860 10081 24869 10115
rect 24869 10081 24903 10115
rect 24903 10081 24912 10115
rect 24860 10072 24912 10081
rect 26516 10115 26568 10124
rect 26516 10081 26525 10115
rect 26525 10081 26559 10115
rect 26559 10081 26568 10115
rect 26516 10072 26568 10081
rect 19248 10004 19300 10056
rect 20812 10004 20864 10056
rect 21916 10047 21968 10056
rect 18328 9936 18380 9988
rect 21916 10013 21925 10047
rect 21925 10013 21959 10047
rect 21959 10013 21968 10047
rect 21916 10004 21968 10013
rect 24032 10004 24084 10056
rect 24676 10047 24728 10056
rect 24676 10013 24685 10047
rect 24685 10013 24719 10047
rect 24719 10013 24728 10047
rect 24676 10004 24728 10013
rect 31392 10047 31444 10056
rect 31392 10013 31401 10047
rect 31401 10013 31435 10047
rect 31435 10013 31444 10047
rect 31392 10004 31444 10013
rect 33140 10047 33192 10056
rect 33140 10013 33149 10047
rect 33149 10013 33183 10047
rect 33183 10013 33192 10047
rect 33140 10004 33192 10013
rect 25872 9979 25924 9988
rect 25872 9945 25881 9979
rect 25881 9945 25915 9979
rect 25915 9945 25924 9979
rect 25872 9936 25924 9945
rect 26240 9936 26292 9988
rect 6368 9868 6420 9920
rect 11980 9868 12032 9920
rect 13728 9868 13780 9920
rect 17500 9868 17552 9920
rect 20260 9868 20312 9920
rect 22376 9911 22428 9920
rect 22376 9877 22385 9911
rect 22385 9877 22419 9911
rect 22419 9877 22428 9911
rect 22376 9868 22428 9877
rect 25504 9868 25556 9920
rect 32864 9868 32916 9920
rect 38016 9868 38068 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 3792 9596 3844 9648
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 6000 9528 6052 9580
rect 6368 9664 6420 9716
rect 9680 9664 9732 9716
rect 9772 9664 9824 9716
rect 9036 9596 9088 9648
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 6460 9460 6512 9512
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 8392 9460 8444 9512
rect 10784 9596 10836 9648
rect 12532 9596 12584 9648
rect 14924 9596 14976 9648
rect 15752 9596 15804 9648
rect 16672 9596 16724 9648
rect 6920 9324 6972 9376
rect 13820 9528 13872 9580
rect 15936 9528 15988 9580
rect 16948 9528 17000 9580
rect 11980 9503 12032 9512
rect 10048 9324 10100 9376
rect 11520 9324 11572 9376
rect 11980 9469 11989 9503
rect 11989 9469 12023 9503
rect 12023 9469 12032 9503
rect 11980 9460 12032 9469
rect 13728 9503 13780 9512
rect 13728 9469 13737 9503
rect 13737 9469 13771 9503
rect 13771 9469 13780 9503
rect 13728 9460 13780 9469
rect 13176 9324 13228 9376
rect 17408 9596 17460 9648
rect 23572 9664 23624 9716
rect 24768 9664 24820 9716
rect 26240 9664 26292 9716
rect 18236 9596 18288 9648
rect 19340 9596 19392 9648
rect 19984 9596 20036 9648
rect 17224 9503 17276 9512
rect 17224 9469 17233 9503
rect 17233 9469 17267 9503
rect 17267 9469 17276 9503
rect 17224 9460 17276 9469
rect 17316 9460 17368 9512
rect 18972 9503 19024 9512
rect 18972 9469 18981 9503
rect 18981 9469 19015 9503
rect 19015 9469 19024 9503
rect 18972 9460 19024 9469
rect 19248 9528 19300 9580
rect 23020 9528 23072 9580
rect 25504 9596 25556 9648
rect 29552 9596 29604 9648
rect 25320 9571 25372 9580
rect 25320 9537 25329 9571
rect 25329 9537 25363 9571
rect 25363 9537 25372 9571
rect 25320 9528 25372 9537
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 20720 9460 20772 9512
rect 23204 9460 23256 9512
rect 15568 9392 15620 9444
rect 20536 9392 20588 9444
rect 27896 9528 27948 9580
rect 33048 9528 33100 9580
rect 15844 9324 15896 9376
rect 16028 9324 16080 9376
rect 16764 9324 16816 9376
rect 17776 9324 17828 9376
rect 18052 9324 18104 9376
rect 20720 9324 20772 9376
rect 20996 9367 21048 9376
rect 20996 9333 21005 9367
rect 21005 9333 21039 9367
rect 21039 9333 21048 9367
rect 20996 9324 21048 9333
rect 22100 9367 22152 9376
rect 22100 9333 22109 9367
rect 22109 9333 22143 9367
rect 22143 9333 22152 9367
rect 22100 9324 22152 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4620 9120 4672 9172
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 6736 9163 6788 9172
rect 6736 9129 6745 9163
rect 6745 9129 6779 9163
rect 6779 9129 6788 9163
rect 6736 9120 6788 9129
rect 6828 9120 6880 9172
rect 1860 9052 1912 9104
rect 11796 9052 11848 9104
rect 8392 8984 8444 9036
rect 15108 9052 15160 9104
rect 15292 9095 15344 9104
rect 15292 9061 15301 9095
rect 15301 9061 15335 9095
rect 15335 9061 15344 9095
rect 15292 9052 15344 9061
rect 15384 9052 15436 9104
rect 16396 9052 16448 9104
rect 17960 9120 18012 9172
rect 18236 9120 18288 9172
rect 16948 9052 17000 9104
rect 17040 9052 17092 9104
rect 24952 9120 25004 9172
rect 25044 9120 25096 9172
rect 14096 8984 14148 9036
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 6828 8916 6880 8968
rect 15108 8916 15160 8968
rect 15752 8916 15804 8968
rect 16028 8984 16080 9036
rect 18972 8984 19024 9036
rect 22008 8984 22060 9036
rect 23204 9027 23256 9036
rect 23204 8993 23213 9027
rect 23213 8993 23247 9027
rect 23247 8993 23256 9027
rect 23204 8984 23256 8993
rect 16672 8916 16724 8968
rect 17500 8916 17552 8968
rect 17684 8916 17736 8968
rect 3976 8848 4028 8900
rect 7564 8848 7616 8900
rect 8208 8848 8260 8900
rect 15936 8848 15988 8900
rect 6000 8780 6052 8832
rect 11520 8780 11572 8832
rect 11980 8780 12032 8832
rect 16488 8780 16540 8832
rect 16948 8780 17000 8832
rect 19432 8780 19484 8832
rect 20260 8823 20312 8832
rect 20260 8789 20269 8823
rect 20269 8789 20303 8823
rect 20303 8789 20312 8823
rect 20260 8780 20312 8789
rect 20812 8959 20864 8968
rect 20812 8925 20821 8959
rect 20821 8925 20855 8959
rect 20855 8925 20864 8959
rect 20812 8916 20864 8925
rect 20996 8848 21048 8900
rect 22100 8891 22152 8900
rect 22100 8857 22109 8891
rect 22109 8857 22143 8891
rect 22143 8857 22152 8891
rect 22100 8848 22152 8857
rect 23572 8848 23624 8900
rect 24768 8984 24820 9036
rect 24952 8916 25004 8968
rect 26148 8959 26200 8968
rect 26148 8925 26157 8959
rect 26157 8925 26191 8959
rect 26191 8925 26200 8959
rect 26148 8916 26200 8925
rect 32864 8916 32916 8968
rect 28724 8848 28776 8900
rect 22836 8780 22888 8832
rect 25228 8823 25280 8832
rect 25228 8789 25237 8823
rect 25237 8789 25271 8823
rect 25271 8789 25280 8823
rect 25228 8780 25280 8789
rect 30288 8780 30340 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 6644 8576 6696 8628
rect 21916 8576 21968 8628
rect 23572 8619 23624 8628
rect 23572 8585 23581 8619
rect 23581 8585 23615 8619
rect 23615 8585 23624 8619
rect 23572 8576 23624 8585
rect 8208 8508 8260 8560
rect 9588 8508 9640 8560
rect 6828 8440 6880 8492
rect 8300 8483 8352 8492
rect 8300 8449 8309 8483
rect 8309 8449 8343 8483
rect 8343 8449 8352 8483
rect 8300 8440 8352 8449
rect 9404 8440 9456 8492
rect 13820 8508 13872 8560
rect 3332 8372 3384 8424
rect 10140 8372 10192 8424
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 13636 8372 13688 8424
rect 17500 8508 17552 8560
rect 17684 8508 17736 8560
rect 22376 8508 22428 8560
rect 22836 8508 22888 8560
rect 27896 8508 27948 8560
rect 15476 8483 15528 8492
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15476 8440 15528 8449
rect 16028 8440 16080 8492
rect 16764 8440 16816 8492
rect 23020 8483 23072 8492
rect 17500 8415 17552 8424
rect 1768 8347 1820 8356
rect 1768 8313 1777 8347
rect 1777 8313 1811 8347
rect 1811 8313 1820 8347
rect 1768 8304 1820 8313
rect 3148 8304 3200 8356
rect 6644 8304 6696 8356
rect 17500 8381 17509 8415
rect 17509 8381 17543 8415
rect 17543 8381 17552 8415
rect 17500 8372 17552 8381
rect 23020 8449 23029 8483
rect 23029 8449 23063 8483
rect 23063 8449 23072 8483
rect 23020 8440 23072 8449
rect 25228 8440 25280 8492
rect 25136 8415 25188 8424
rect 15752 8304 15804 8356
rect 25136 8381 25145 8415
rect 25145 8381 25179 8415
rect 25179 8381 25188 8415
rect 25136 8372 25188 8381
rect 25504 8347 25556 8356
rect 25504 8313 25513 8347
rect 25513 8313 25547 8347
rect 25547 8313 25556 8347
rect 25504 8304 25556 8313
rect 16028 8236 16080 8288
rect 16396 8236 16448 8288
rect 16488 8236 16540 8288
rect 16672 8236 16724 8288
rect 17684 8236 17736 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 8668 8032 8720 8084
rect 9036 8032 9088 8084
rect 13176 8075 13228 8084
rect 13176 8041 13185 8075
rect 13185 8041 13219 8075
rect 13219 8041 13228 8075
rect 13176 8032 13228 8041
rect 14648 8032 14700 8084
rect 16672 8032 16724 8084
rect 3792 7964 3844 8016
rect 16948 7964 17000 8016
rect 5816 7896 5868 7948
rect 5356 7828 5408 7880
rect 9772 7828 9824 7880
rect 17776 7896 17828 7948
rect 12624 7828 12676 7880
rect 17040 7828 17092 7880
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 24676 8032 24728 8084
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 25136 7939 25188 7948
rect 25136 7905 25145 7939
rect 25145 7905 25179 7939
rect 25179 7905 25188 7939
rect 25136 7896 25188 7905
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 27896 7828 27948 7880
rect 28724 7871 28776 7880
rect 28724 7837 28733 7871
rect 28733 7837 28767 7871
rect 28767 7837 28776 7871
rect 28724 7828 28776 7837
rect 14464 7803 14516 7812
rect 14464 7769 14473 7803
rect 14473 7769 14507 7803
rect 14507 7769 14516 7803
rect 14464 7760 14516 7769
rect 15108 7803 15160 7812
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 13084 7692 13136 7744
rect 15108 7769 15117 7803
rect 15117 7769 15151 7803
rect 15151 7769 15160 7803
rect 15108 7760 15160 7769
rect 15476 7692 15528 7744
rect 16672 7760 16724 7812
rect 23480 7760 23532 7812
rect 31668 7692 31720 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 12992 7531 13044 7540
rect 12992 7497 13001 7531
rect 13001 7497 13035 7531
rect 13035 7497 13044 7531
rect 12992 7488 13044 7497
rect 14464 7531 14516 7540
rect 14464 7497 14473 7531
rect 14473 7497 14507 7531
rect 14507 7497 14516 7531
rect 14464 7488 14516 7497
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 3424 7352 3476 7404
rect 9864 7420 9916 7472
rect 10324 7420 10376 7472
rect 19340 7488 19392 7540
rect 22008 7531 22060 7540
rect 22008 7497 22017 7531
rect 22017 7497 22051 7531
rect 22051 7497 22060 7531
rect 22008 7488 22060 7497
rect 22192 7488 22244 7540
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 12624 7352 12676 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 13084 7352 13136 7404
rect 20352 7420 20404 7472
rect 16764 7352 16816 7404
rect 17040 7352 17092 7404
rect 22836 7395 22888 7404
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 11980 7284 12032 7336
rect 10784 7216 10836 7268
rect 17316 7284 17368 7336
rect 20628 7284 20680 7336
rect 17408 7216 17460 7268
rect 19340 7216 19392 7268
rect 22836 7361 22845 7395
rect 22845 7361 22879 7395
rect 22879 7361 22888 7395
rect 22836 7352 22888 7361
rect 23388 7395 23440 7404
rect 23388 7361 23397 7395
rect 23397 7361 23431 7395
rect 23431 7361 23440 7395
rect 23388 7352 23440 7361
rect 34060 7352 34112 7404
rect 24032 7327 24084 7336
rect 24032 7293 24041 7327
rect 24041 7293 24075 7327
rect 24075 7293 24084 7327
rect 24032 7284 24084 7293
rect 4620 7148 4672 7200
rect 5540 7148 5592 7200
rect 16304 7148 16356 7200
rect 17868 7148 17920 7200
rect 24400 7191 24452 7200
rect 24400 7157 24409 7191
rect 24409 7157 24443 7191
rect 24443 7157 24452 7191
rect 24400 7148 24452 7157
rect 38200 7191 38252 7200
rect 38200 7157 38209 7191
rect 38209 7157 38243 7191
rect 38243 7157 38252 7191
rect 38200 7148 38252 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 6000 6987 6052 6996
rect 6000 6953 6009 6987
rect 6009 6953 6043 6987
rect 6043 6953 6052 6987
rect 6000 6944 6052 6953
rect 7196 6944 7248 6996
rect 7840 6944 7892 6996
rect 15476 6987 15528 6996
rect 9220 6851 9272 6860
rect 9220 6817 9229 6851
rect 9229 6817 9263 6851
rect 9263 6817 9272 6851
rect 9220 6808 9272 6817
rect 10968 6876 11020 6928
rect 15476 6953 15485 6987
rect 15485 6953 15519 6987
rect 15519 6953 15528 6987
rect 15476 6944 15528 6953
rect 16948 6944 17000 6996
rect 19248 6944 19300 6996
rect 17040 6876 17092 6928
rect 20628 6876 20680 6928
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 11612 6808 11664 6860
rect 17500 6808 17552 6860
rect 19524 6851 19576 6860
rect 19524 6817 19533 6851
rect 19533 6817 19567 6851
rect 19567 6817 19576 6851
rect 19524 6808 19576 6817
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 12256 6740 12308 6792
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 16120 6740 16172 6792
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 5632 6672 5684 6724
rect 2688 6647 2740 6656
rect 2688 6613 2697 6647
rect 2697 6613 2731 6647
rect 2731 6613 2740 6647
rect 2688 6604 2740 6613
rect 5816 6604 5868 6656
rect 6460 6604 6512 6656
rect 7196 6647 7248 6656
rect 7196 6613 7205 6647
rect 7205 6613 7239 6647
rect 7239 6613 7248 6647
rect 7196 6604 7248 6613
rect 7380 6604 7432 6656
rect 7932 6604 7984 6656
rect 13544 6672 13596 6724
rect 17776 6715 17828 6724
rect 12164 6604 12216 6656
rect 14556 6604 14608 6656
rect 16764 6604 16816 6656
rect 17776 6681 17785 6715
rect 17785 6681 17819 6715
rect 17819 6681 17828 6715
rect 17776 6672 17828 6681
rect 17868 6715 17920 6724
rect 17868 6681 17877 6715
rect 17877 6681 17911 6715
rect 17911 6681 17920 6715
rect 17868 6672 17920 6681
rect 18052 6672 18104 6724
rect 19064 6604 19116 6656
rect 20536 6740 20588 6792
rect 19524 6672 19576 6724
rect 23388 6740 23440 6792
rect 23480 6740 23532 6792
rect 27528 6740 27580 6792
rect 29828 6672 29880 6724
rect 22284 6604 22336 6656
rect 23480 6604 23532 6656
rect 23756 6647 23808 6656
rect 23756 6613 23765 6647
rect 23765 6613 23799 6647
rect 23799 6613 23808 6647
rect 23756 6604 23808 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 6736 6443 6788 6452
rect 6736 6409 6745 6443
rect 6745 6409 6779 6443
rect 6779 6409 6788 6443
rect 6736 6400 6788 6409
rect 5540 6332 5592 6384
rect 10784 6400 10836 6452
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 15660 6400 15712 6452
rect 16948 6400 17000 6452
rect 19432 6400 19484 6452
rect 20352 6443 20404 6452
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 7748 6332 7800 6384
rect 7840 6332 7892 6384
rect 9772 6332 9824 6384
rect 13268 6332 13320 6384
rect 15752 6375 15804 6384
rect 15752 6341 15761 6375
rect 15761 6341 15795 6375
rect 15795 6341 15804 6375
rect 15752 6332 15804 6341
rect 20352 6409 20361 6443
rect 20361 6409 20395 6443
rect 20395 6409 20404 6443
rect 20352 6400 20404 6409
rect 23388 6443 23440 6452
rect 23388 6409 23397 6443
rect 23397 6409 23431 6443
rect 23431 6409 23440 6443
rect 23388 6400 23440 6409
rect 24032 6400 24084 6452
rect 7196 6264 7248 6316
rect 10140 6264 10192 6316
rect 12164 6264 12216 6316
rect 14924 6307 14976 6316
rect 14924 6273 14933 6307
rect 14933 6273 14967 6307
rect 14967 6273 14976 6307
rect 14924 6264 14976 6273
rect 16396 6264 16448 6316
rect 17132 6264 17184 6316
rect 18972 6264 19024 6316
rect 19064 6264 19116 6316
rect 23480 6332 23532 6384
rect 24400 6332 24452 6384
rect 23756 6264 23808 6316
rect 27160 6264 27212 6316
rect 1768 6171 1820 6180
rect 1768 6137 1777 6171
rect 1777 6137 1811 6171
rect 1811 6137 1820 6171
rect 1768 6128 1820 6137
rect 5816 6196 5868 6248
rect 12072 6196 12124 6248
rect 12440 6196 12492 6248
rect 13728 6196 13780 6248
rect 17408 6196 17460 6248
rect 20076 6196 20128 6248
rect 7196 6128 7248 6180
rect 11612 6128 11664 6180
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 2412 6060 2464 6069
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 7748 6060 7800 6112
rect 15108 6128 15160 6180
rect 17776 6128 17828 6180
rect 26516 6128 26568 6180
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 14464 6060 14516 6112
rect 18880 6060 18932 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 6276 5856 6328 5908
rect 7840 5899 7892 5908
rect 7840 5865 7849 5899
rect 7849 5865 7883 5899
rect 7883 5865 7892 5899
rect 7840 5856 7892 5865
rect 7932 5856 7984 5908
rect 12256 5899 12308 5908
rect 2412 5788 2464 5840
rect 7196 5788 7248 5840
rect 11704 5788 11756 5840
rect 12256 5865 12265 5899
rect 12265 5865 12299 5899
rect 12299 5865 12308 5899
rect 12256 5856 12308 5865
rect 12348 5856 12400 5908
rect 17408 5856 17460 5908
rect 12440 5788 12492 5840
rect 13544 5831 13596 5840
rect 4620 5652 4672 5704
rect 8300 5720 8352 5772
rect 2780 5584 2832 5636
rect 8484 5652 8536 5704
rect 13544 5797 13553 5831
rect 13553 5797 13587 5831
rect 13587 5797 13596 5831
rect 13544 5788 13596 5797
rect 14188 5720 14240 5772
rect 19340 5788 19392 5840
rect 26608 5856 26660 5908
rect 29828 5899 29880 5908
rect 29828 5865 29837 5899
rect 29837 5865 29871 5899
rect 29871 5865 29880 5899
rect 29828 5856 29880 5865
rect 23480 5788 23532 5840
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 14464 5720 14516 5729
rect 14556 5720 14608 5772
rect 20996 5720 21048 5772
rect 26332 5720 26384 5772
rect 12532 5584 12584 5636
rect 12808 5584 12860 5636
rect 14924 5652 14976 5704
rect 16856 5652 16908 5704
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 36728 5652 36780 5704
rect 37188 5652 37240 5704
rect 16580 5627 16632 5636
rect 16580 5593 16589 5627
rect 16589 5593 16623 5627
rect 16623 5593 16632 5627
rect 16580 5584 16632 5593
rect 2872 5516 2924 5568
rect 11520 5516 11572 5568
rect 20076 5516 20128 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 6460 5176 6512 5228
rect 17868 5312 17920 5364
rect 7380 5287 7432 5296
rect 7380 5253 7389 5287
rect 7389 5253 7423 5287
rect 7423 5253 7432 5287
rect 7380 5244 7432 5253
rect 12900 5244 12952 5296
rect 30288 5244 30340 5296
rect 10140 5219 10192 5228
rect 10140 5185 10149 5219
rect 10149 5185 10183 5219
rect 10183 5185 10192 5219
rect 10140 5176 10192 5185
rect 12348 5176 12400 5228
rect 7288 5151 7340 5160
rect 7288 5117 7297 5151
rect 7297 5117 7331 5151
rect 7331 5117 7340 5151
rect 7288 5108 7340 5117
rect 11980 5108 12032 5160
rect 18420 5176 18472 5228
rect 31668 5219 31720 5228
rect 31668 5185 31677 5219
rect 31677 5185 31711 5219
rect 31711 5185 31720 5219
rect 31668 5176 31720 5185
rect 33692 5040 33744 5092
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 6644 5015 6696 5024
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 14280 4972 14332 5024
rect 34060 4972 34112 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 13728 4564 13780 4616
rect 35624 4564 35676 4616
rect 11152 4471 11204 4480
rect 11152 4437 11161 4471
rect 11161 4437 11195 4471
rect 11195 4437 11204 4471
rect 11152 4428 11204 4437
rect 11888 4471 11940 4480
rect 11888 4437 11897 4471
rect 11897 4437 11931 4471
rect 11931 4437 11940 4471
rect 11888 4428 11940 4437
rect 18328 4428 18380 4480
rect 27804 4471 27856 4480
rect 27804 4437 27813 4471
rect 27813 4437 27847 4471
rect 27847 4437 27856 4471
rect 27804 4428 27856 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 12348 4267 12400 4276
rect 12348 4233 12357 4267
rect 12357 4233 12391 4267
rect 12391 4233 12400 4267
rect 12348 4224 12400 4233
rect 11152 4088 11204 4140
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 16856 4088 16908 4140
rect 16948 3952 17000 4004
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2780 3680 2832 3732
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 6644 3519 6696 3528
rect 6644 3485 6653 3519
rect 6653 3485 6687 3519
rect 6687 3485 6696 3519
rect 6644 3476 6696 3485
rect 17592 3476 17644 3528
rect 38016 3519 38068 3528
rect 38016 3485 38025 3519
rect 38025 3485 38059 3519
rect 38059 3485 38068 3519
rect 38016 3476 38068 3485
rect 21180 3408 21232 3460
rect 6552 3340 6604 3392
rect 11060 3340 11112 3392
rect 18604 3340 18656 3392
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 7288 3136 7340 3188
rect 16672 3136 16724 3188
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 17592 3179 17644 3188
rect 17592 3145 17601 3179
rect 17601 3145 17635 3179
rect 17635 3145 17644 3179
rect 17592 3136 17644 3145
rect 36728 3179 36780 3188
rect 36728 3145 36737 3179
rect 36737 3145 36771 3179
rect 36771 3145 36780 3179
rect 36728 3136 36780 3145
rect 2872 3068 2924 3120
rect 2780 3000 2832 3052
rect 11796 3068 11848 3120
rect 18328 3111 18380 3120
rect 18328 3077 18337 3111
rect 18337 3077 18371 3111
rect 18371 3077 18380 3111
rect 18328 3068 18380 3077
rect 34060 3068 34112 3120
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11152 3000 11204 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17224 3000 17276 3052
rect 36912 3043 36964 3052
rect 36912 3009 36921 3043
rect 36921 3009 36955 3043
rect 36955 3009 36964 3043
rect 36912 3000 36964 3009
rect 27804 2932 27856 2984
rect 8300 2864 8352 2916
rect 11980 2864 12032 2916
rect 20 2796 72 2848
rect 9128 2796 9180 2848
rect 38200 2839 38252 2848
rect 38200 2805 38209 2839
rect 38209 2805 38243 2839
rect 38243 2805 38252 2839
rect 38200 2796 38252 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4712 2592 4764 2644
rect 11152 2592 11204 2644
rect 17132 2592 17184 2644
rect 21272 2592 21324 2644
rect 23848 2592 23900 2644
rect 27160 2635 27212 2644
rect 27160 2601 27169 2635
rect 27169 2601 27203 2635
rect 27203 2601 27212 2635
rect 27160 2592 27212 2601
rect 27528 2592 27580 2644
rect 29736 2635 29788 2644
rect 29736 2601 29745 2635
rect 29745 2601 29779 2635
rect 29779 2601 29788 2635
rect 29736 2592 29788 2601
rect 32312 2635 32364 2644
rect 32312 2601 32321 2635
rect 32321 2601 32355 2635
rect 32355 2601 32364 2635
rect 32312 2592 32364 2601
rect 33048 2592 33100 2644
rect 35624 2592 35676 2644
rect 4804 2524 4856 2576
rect 10140 2524 10192 2576
rect 27896 2524 27948 2576
rect 2596 2388 2648 2440
rect 7104 2456 7156 2508
rect 33692 2456 33744 2508
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 8300 2388 8352 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 10324 2388 10376 2440
rect 12256 2388 12308 2440
rect 14280 2431 14332 2440
rect 14280 2397 14289 2431
rect 14289 2397 14323 2431
rect 14323 2397 14332 2431
rect 14280 2388 14332 2397
rect 15476 2388 15528 2440
rect 16764 2388 16816 2440
rect 18604 2431 18656 2440
rect 18604 2397 18613 2431
rect 18613 2397 18647 2431
rect 18647 2397 18656 2431
rect 18604 2388 18656 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 21272 2388 21324 2440
rect 22284 2388 22336 2440
rect 24492 2388 24544 2440
rect 26424 2388 26476 2440
rect 27712 2388 27764 2440
rect 29000 2388 29052 2440
rect 30932 2388 30984 2440
rect 32220 2388 32272 2440
rect 34152 2388 34204 2440
rect 35440 2388 35492 2440
rect 26148 2320 26200 2372
rect 1308 2252 1360 2304
rect 4528 2252 4580 2304
rect 5816 2252 5868 2304
rect 7748 2252 7800 2304
rect 9036 2252 9088 2304
rect 13544 2252 13596 2304
rect 16764 2252 16816 2304
rect 18696 2252 18748 2304
rect 19984 2252 20036 2304
rect 23204 2252 23256 2304
rect 38660 2320 38712 2372
rect 37372 2252 37424 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 2778 39536 2834 39545
rect 2778 39471 2834 39480
rect 676 36922 704 39200
rect 1964 37262 1992 39200
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 664 36916 716 36922
rect 664 36858 716 36864
rect 1596 34746 1624 37198
rect 2792 37194 2820 39471
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 20626 39200 20682 39800
rect 22558 39200 22614 39800
rect 23846 39200 23902 39800
rect 25778 39200 25834 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 31574 39200 31630 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 3146 37496 3202 37505
rect 3146 37431 3202 37440
rect 3160 37262 3188 37431
rect 3148 37256 3200 37262
rect 3896 37244 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5184 37262 5212 39200
rect 7116 37262 7144 39200
rect 8404 37262 8432 39200
rect 10336 37262 10364 39200
rect 11624 37262 11652 39200
rect 4160 37256 4212 37262
rect 3896 37216 4160 37244
rect 3148 37198 3200 37204
rect 4160 37198 4212 37204
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 10324 37256 10376 37262
rect 10324 37198 10376 37204
rect 11612 37256 11664 37262
rect 11612 37198 11664 37204
rect 11980 37256 12032 37262
rect 11980 37198 12032 37204
rect 2780 37188 2832 37194
rect 2780 37130 2832 37136
rect 6828 37188 6880 37194
rect 6828 37130 6880 37136
rect 2320 37120 2372 37126
rect 2320 37062 2372 37068
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 1768 36168 1820 36174
rect 1766 36136 1768 36145
rect 1820 36136 1822 36145
rect 1766 36071 1822 36080
rect 1584 34740 1636 34746
rect 1584 34682 1636 34688
rect 1952 34604 2004 34610
rect 1952 34546 2004 34552
rect 1766 34096 1822 34105
rect 1766 34031 1822 34040
rect 1780 33998 1808 34031
rect 1768 33992 1820 33998
rect 1768 33934 1820 33940
rect 1676 33856 1728 33862
rect 1676 33798 1728 33804
rect 1492 32428 1544 32434
rect 1492 32370 1544 32376
rect 1504 16454 1532 32370
rect 1584 30048 1636 30054
rect 1584 29990 1636 29996
rect 1596 28082 1624 29990
rect 1584 28076 1636 28082
rect 1584 28018 1636 28024
rect 1688 26994 1716 33798
rect 1964 33658 1992 34546
rect 1952 33652 2004 33658
rect 1952 33594 2004 33600
rect 2136 33516 2188 33522
rect 2136 33458 2188 33464
rect 1768 32904 1820 32910
rect 1768 32846 1820 32852
rect 1780 32745 1808 32846
rect 1860 32768 1912 32774
rect 1766 32736 1822 32745
rect 1860 32710 1912 32716
rect 1766 32671 1822 32680
rect 1766 30696 1822 30705
rect 1766 30631 1822 30640
rect 1780 30258 1808 30631
rect 1768 30252 1820 30258
rect 1768 30194 1820 30200
rect 1872 29646 1900 32710
rect 1952 32224 2004 32230
rect 1952 32166 2004 32172
rect 1964 31793 1992 32166
rect 1950 31784 2006 31793
rect 1950 31719 2006 31728
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 1964 30938 1992 31282
rect 1952 30932 2004 30938
rect 1952 30874 2004 30880
rect 1860 29640 1912 29646
rect 2148 29594 2176 33458
rect 2228 33312 2280 33318
rect 2228 33254 2280 33260
rect 1860 29582 1912 29588
rect 1964 29566 2176 29594
rect 1766 29336 1822 29345
rect 1766 29271 1822 29280
rect 1780 29170 1808 29271
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1964 29050 1992 29566
rect 2136 29504 2188 29510
rect 2136 29446 2188 29452
rect 1872 29022 1992 29050
rect 1766 27976 1822 27985
rect 1766 27911 1822 27920
rect 1780 27470 1808 27911
rect 1768 27464 1820 27470
rect 1768 27406 1820 27412
rect 1676 26988 1728 26994
rect 1676 26930 1728 26936
rect 1872 26874 1900 29022
rect 1952 28960 2004 28966
rect 1952 28902 2004 28908
rect 1964 28558 1992 28902
rect 1952 28552 2004 28558
rect 1952 28494 2004 28500
rect 1952 28416 2004 28422
rect 1952 28358 2004 28364
rect 1688 26846 1900 26874
rect 1584 23112 1636 23118
rect 1584 23054 1636 23060
rect 1596 20602 1624 23054
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1584 18216 1636 18222
rect 1584 18158 1636 18164
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1596 16114 1624 18158
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1596 15026 1624 16050
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1596 14385 1624 14962
rect 1582 14376 1638 14385
rect 1582 14311 1638 14320
rect 1596 13938 1624 14311
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1688 11218 1716 26846
rect 1860 26784 1912 26790
rect 1860 26726 1912 26732
rect 1872 26450 1900 26726
rect 1860 26444 1912 26450
rect 1860 26386 1912 26392
rect 1860 25832 1912 25838
rect 1860 25774 1912 25780
rect 1766 24576 1822 24585
rect 1766 24511 1822 24520
rect 1780 24410 1808 24511
rect 1768 24404 1820 24410
rect 1768 24346 1820 24352
rect 1872 24274 1900 25774
rect 1860 24268 1912 24274
rect 1860 24210 1912 24216
rect 1964 24206 1992 28358
rect 1952 24200 2004 24206
rect 1952 24142 2004 24148
rect 1768 22976 1820 22982
rect 1768 22918 1820 22924
rect 1780 22545 1808 22918
rect 2148 22574 2176 29446
rect 2240 25838 2268 33254
rect 2332 29170 2360 37062
rect 2872 36780 2924 36786
rect 2872 36722 2924 36728
rect 2884 33114 2912 36722
rect 3516 36032 3568 36038
rect 3516 35974 3568 35980
rect 3056 33448 3108 33454
rect 3056 33390 3108 33396
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2872 31952 2924 31958
rect 2872 31894 2924 31900
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2504 31136 2556 31142
rect 2504 31078 2556 31084
rect 2412 30592 2464 30598
rect 2412 30534 2464 30540
rect 2320 29164 2372 29170
rect 2320 29106 2372 29112
rect 2424 25906 2452 30534
rect 2516 26450 2544 31078
rect 2792 30734 2820 31758
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 2596 30252 2648 30258
rect 2596 30194 2648 30200
rect 2608 29102 2636 30194
rect 2780 30116 2832 30122
rect 2780 30058 2832 30064
rect 2792 29714 2820 30058
rect 2780 29708 2832 29714
rect 2780 29650 2832 29656
rect 2884 29578 2912 31894
rect 3068 29714 3096 33390
rect 3148 30592 3200 30598
rect 3148 30534 3200 30540
rect 3056 29708 3108 29714
rect 3056 29650 3108 29656
rect 2872 29572 2924 29578
rect 2872 29514 2924 29520
rect 2596 29096 2648 29102
rect 2596 29038 2648 29044
rect 2504 26444 2556 26450
rect 2504 26386 2556 26392
rect 2412 25900 2464 25906
rect 2412 25842 2464 25848
rect 2228 25832 2280 25838
rect 2228 25774 2280 25780
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2136 22568 2188 22574
rect 1766 22536 1822 22545
rect 2136 22510 2188 22516
rect 1766 22471 1822 22480
rect 2228 22092 2280 22098
rect 2228 22034 2280 22040
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1780 21185 1808 21490
rect 1766 21176 1822 21185
rect 1766 21111 1822 21120
rect 1950 20496 2006 20505
rect 1950 20431 1952 20440
rect 2004 20431 2006 20440
rect 1952 20402 2004 20408
rect 2240 19854 2268 22034
rect 2412 21344 2464 21350
rect 2412 21286 2464 21292
rect 1768 19848 1820 19854
rect 1766 19816 1768 19825
rect 2228 19848 2280 19854
rect 1820 19816 1822 19825
rect 2228 19790 2280 19796
rect 1766 19751 1822 19760
rect 2240 19310 2268 19790
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17785 1808 18226
rect 2240 18222 2268 19246
rect 2424 18766 2452 21286
rect 2516 19310 2544 25230
rect 2608 24750 2636 29038
rect 3068 28218 3096 29650
rect 3056 28212 3108 28218
rect 3056 28154 3108 28160
rect 3160 28150 3188 30534
rect 3528 28626 3556 35974
rect 3700 31680 3752 31686
rect 3700 31622 3752 31628
rect 3516 28620 3568 28626
rect 3516 28562 3568 28568
rect 3148 28144 3200 28150
rect 3148 28086 3200 28092
rect 3056 28008 3108 28014
rect 3056 27950 3108 27956
rect 3516 28008 3568 28014
rect 3516 27950 3568 27956
rect 3068 26586 3096 27950
rect 3332 27872 3384 27878
rect 3332 27814 3384 27820
rect 3056 26580 3108 26586
rect 3056 26522 3108 26528
rect 2964 26240 3016 26246
rect 2964 26182 3016 26188
rect 2976 25362 3004 26182
rect 3068 26042 3096 26522
rect 3148 26376 3200 26382
rect 3148 26318 3200 26324
rect 3056 26036 3108 26042
rect 3056 25978 3108 25984
rect 3160 25945 3188 26318
rect 3146 25936 3202 25945
rect 3146 25871 3202 25880
rect 3344 25362 3372 27814
rect 3424 25696 3476 25702
rect 3424 25638 3476 25644
rect 2964 25356 3016 25362
rect 2964 25298 3016 25304
rect 3332 25356 3384 25362
rect 3332 25298 3384 25304
rect 3332 25220 3384 25226
rect 3332 25162 3384 25168
rect 2688 25152 2740 25158
rect 2688 25094 2740 25100
rect 2596 24744 2648 24750
rect 2596 24686 2648 24692
rect 2700 22710 2728 25094
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2792 23662 2820 24550
rect 2872 24200 2924 24206
rect 2872 24142 2924 24148
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2688 22704 2740 22710
rect 2688 22646 2740 22652
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2792 21010 2820 21286
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2884 20058 2912 24142
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 3344 18426 3372 25162
rect 3436 25158 3464 25638
rect 3528 25430 3556 27950
rect 3516 25424 3568 25430
rect 3516 25366 3568 25372
rect 3712 25226 3740 31622
rect 3896 30734 3924 37062
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 32434 4660 37062
rect 6184 32904 6236 32910
rect 6184 32846 6236 32852
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 5460 32026 5488 32302
rect 5448 32020 5500 32026
rect 5448 31962 5500 31968
rect 5264 31816 5316 31822
rect 5264 31758 5316 31764
rect 5276 31482 5304 31758
rect 5264 31476 5316 31482
rect 5264 31418 5316 31424
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3884 30728 3936 30734
rect 3884 30670 3936 30676
rect 4620 30660 4672 30666
rect 4620 30602 4672 30608
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 4172 30190 4200 30534
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3976 29640 4028 29646
rect 3976 29582 4028 29588
rect 3792 28144 3844 28150
rect 3792 28086 3844 28092
rect 3804 25498 3832 28086
rect 3988 27606 4016 29582
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3976 27600 4028 27606
rect 3976 27542 4028 27548
rect 4068 27396 4120 27402
rect 4068 27338 4120 27344
rect 4344 27396 4396 27402
rect 4344 27338 4396 27344
rect 3976 25832 4028 25838
rect 3976 25774 4028 25780
rect 3792 25492 3844 25498
rect 3792 25434 3844 25440
rect 3700 25220 3752 25226
rect 3700 25162 3752 25168
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3516 24608 3568 24614
rect 3516 24550 3568 24556
rect 3528 23594 3556 24550
rect 3988 24154 4016 25774
rect 4080 24410 4108 27338
rect 4252 27328 4304 27334
rect 4252 27270 4304 27276
rect 4264 26994 4292 27270
rect 4356 27130 4384 27338
rect 4344 27124 4396 27130
rect 4344 27066 4396 27072
rect 4252 26988 4304 26994
rect 4252 26930 4304 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 4068 24200 4120 24206
rect 3988 24148 4068 24154
rect 3988 24142 4120 24148
rect 3988 24126 4108 24142
rect 3988 23662 4016 24126
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3516 23588 3568 23594
rect 3516 23530 3568 23536
rect 3700 23520 3752 23526
rect 3700 23462 3752 23468
rect 3712 22234 3740 23462
rect 3988 23118 4016 23598
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23186 4660 30602
rect 5080 28552 5132 28558
rect 5080 28494 5132 28500
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3700 22228 3752 22234
rect 3700 22170 3752 22176
rect 3988 21010 4016 23054
rect 4620 22500 4672 22506
rect 4620 22442 4672 22448
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 21962 4660 22442
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 4804 21616 4856 21622
rect 4804 21558 4856 21564
rect 4620 21480 4672 21486
rect 4620 21422 4672 21428
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21010 4660 21422
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 3424 20868 3476 20874
rect 3424 20810 3476 20816
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 1766 17776 1822 17785
rect 1766 17711 1822 17720
rect 1768 16584 1820 16590
rect 2332 16574 2360 18022
rect 2332 16546 2452 16574
rect 1768 16526 1820 16532
rect 1780 16425 1808 16526
rect 1766 16416 1822 16425
rect 1766 16351 1822 16360
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 2148 14278 2176 14894
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 13025 1808 13126
rect 1766 13016 1822 13025
rect 1766 12951 1822 12960
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10985 1624 11086
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1596 9586 1624 10066
rect 1780 9625 1808 10406
rect 1766 9616 1822 9625
rect 1584 9580 1636 9586
rect 1766 9551 1822 9560
rect 1584 9522 1636 9528
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1872 9110 1900 9454
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1780 8265 1808 8298
rect 1766 8256 1822 8265
rect 1766 8191 1822 8200
rect 2424 6914 2452 16546
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2516 13938 2544 14418
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2516 12850 2544 13874
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2516 11762 2544 12786
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2516 10130 2544 11698
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2332 6886 2452 6914
rect 2332 6322 2360 6886
rect 2700 6662 2728 13262
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 3252 12442 3280 12854
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3344 12238 3372 14350
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3344 10062 3372 12174
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3160 8362 3188 9930
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 8430 3372 9318
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3436 7410 3464 20810
rect 4632 20466 4660 20946
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3988 19514 4016 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4632 19786 4660 20402
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3620 15706 3648 15982
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3804 12434 3832 18158
rect 3896 15026 3924 18362
rect 3988 16250 4016 19450
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4080 15638 4108 18294
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17746 4660 18770
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4356 17134 4384 17682
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4080 15026 4108 15438
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14414 4108 14962
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4724 14618 4752 20810
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4816 14550 4844 21558
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4908 18358 4936 18634
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 4896 15088 4948 15094
rect 4896 15030 4948 15036
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4908 14006 4936 15030
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3804 12406 3924 12434
rect 3896 10266 3924 12406
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3988 11218 4016 11698
rect 4080 11354 4108 13806
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3804 8022 3832 9590
rect 3988 8906 4016 9998
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9178 4660 10610
rect 5000 10198 5028 23122
rect 5092 17882 5120 28494
rect 5184 23526 5212 31282
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 5460 30326 5488 31078
rect 5724 30796 5776 30802
rect 5724 30738 5776 30744
rect 5448 30320 5500 30326
rect 5448 30262 5500 30268
rect 5540 29164 5592 29170
rect 5540 29106 5592 29112
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5368 28082 5396 28358
rect 5460 28218 5488 28358
rect 5448 28212 5500 28218
rect 5448 28154 5500 28160
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 5264 26036 5316 26042
rect 5264 25978 5316 25984
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5092 15094 5120 17682
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5184 16658 5212 17070
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 5184 14958 5212 16594
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5184 14482 5212 14894
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5276 14346 5304 25978
rect 5356 25900 5408 25906
rect 5356 25842 5408 25848
rect 5368 25498 5396 25842
rect 5356 25492 5408 25498
rect 5356 25434 5408 25440
rect 5448 25152 5500 25158
rect 5448 25094 5500 25100
rect 5460 23798 5488 25094
rect 5552 24070 5580 29106
rect 5632 28416 5684 28422
rect 5632 28358 5684 28364
rect 5644 27538 5672 28358
rect 5632 27532 5684 27538
rect 5632 27474 5684 27480
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5448 23792 5500 23798
rect 5448 23734 5500 23740
rect 5736 23322 5764 30738
rect 6000 30252 6052 30258
rect 6000 30194 6052 30200
rect 6012 29714 6040 30194
rect 6000 29708 6052 29714
rect 6000 29650 6052 29656
rect 5816 28008 5868 28014
rect 5816 27950 5868 27956
rect 5828 27538 5856 27950
rect 5908 27872 5960 27878
rect 5908 27814 5960 27820
rect 5816 27532 5868 27538
rect 5816 27474 5868 27480
rect 5920 27402 5948 27814
rect 5908 27396 5960 27402
rect 5908 27338 5960 27344
rect 5908 24404 5960 24410
rect 5908 24346 5960 24352
rect 5920 23866 5948 24346
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 5724 23316 5776 23322
rect 5724 23258 5776 23264
rect 5736 22094 5764 23258
rect 5552 22066 5764 22094
rect 5552 19718 5580 22066
rect 6012 21706 6040 29650
rect 6196 27402 6224 32846
rect 6552 32768 6604 32774
rect 6552 32710 6604 32716
rect 6564 32434 6592 32710
rect 6840 32434 6868 37130
rect 7196 37120 7248 37126
rect 7196 37062 7248 37068
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 10416 37120 10468 37126
rect 10416 37062 10468 37068
rect 11704 37120 11756 37126
rect 11704 37062 11756 37068
rect 6552 32428 6604 32434
rect 6552 32370 6604 32376
rect 6828 32428 6880 32434
rect 6828 32370 6880 32376
rect 6736 32360 6788 32366
rect 6736 32302 6788 32308
rect 6748 31482 6776 32302
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 7208 31346 7236 37062
rect 9140 32910 9168 37062
rect 9128 32904 9180 32910
rect 9128 32846 9180 32852
rect 7748 32224 7800 32230
rect 7748 32166 7800 32172
rect 10140 32224 10192 32230
rect 10140 32166 10192 32172
rect 7760 31958 7788 32166
rect 7380 31952 7432 31958
rect 7380 31894 7432 31900
rect 7748 31952 7800 31958
rect 7748 31894 7800 31900
rect 7196 31340 7248 31346
rect 7196 31282 7248 31288
rect 7392 31278 7420 31894
rect 9220 31884 9272 31890
rect 9220 31826 9272 31832
rect 7380 31272 7432 31278
rect 7380 31214 7432 31220
rect 7748 31272 7800 31278
rect 7748 31214 7800 31220
rect 7392 30802 7420 31214
rect 7760 30938 7788 31214
rect 7748 30932 7800 30938
rect 7748 30874 7800 30880
rect 7380 30796 7432 30802
rect 7380 30738 7432 30744
rect 8576 30728 8628 30734
rect 8576 30670 8628 30676
rect 6644 30660 6696 30666
rect 6644 30602 6696 30608
rect 7472 30660 7524 30666
rect 7472 30602 7524 30608
rect 6368 30048 6420 30054
rect 6368 29990 6420 29996
rect 6380 29646 6408 29990
rect 6656 29850 6684 30602
rect 6920 30320 6972 30326
rect 6920 30262 6972 30268
rect 6932 29850 6960 30262
rect 7484 30122 7512 30602
rect 8588 30326 8616 30670
rect 8576 30320 8628 30326
rect 8576 30262 8628 30268
rect 7472 30116 7524 30122
rect 7472 30058 7524 30064
rect 6644 29844 6696 29850
rect 6644 29786 6696 29792
rect 6920 29844 6972 29850
rect 6920 29786 6972 29792
rect 6368 29640 6420 29646
rect 6368 29582 6420 29588
rect 6828 29028 6880 29034
rect 6828 28970 6880 28976
rect 6184 27396 6236 27402
rect 6184 27338 6236 27344
rect 6460 27396 6512 27402
rect 6460 27338 6512 27344
rect 6184 24064 6236 24070
rect 6184 24006 6236 24012
rect 6012 21678 6132 21706
rect 6196 21690 6224 24006
rect 6472 22778 6500 27338
rect 6644 27056 6696 27062
rect 6644 26998 6696 27004
rect 6656 24342 6684 26998
rect 6644 24336 6696 24342
rect 6644 24278 6696 24284
rect 6840 23798 6868 28970
rect 6828 23792 6880 23798
rect 6828 23734 6880 23740
rect 6736 23588 6788 23594
rect 6736 23530 6788 23536
rect 6460 22772 6512 22778
rect 6460 22714 6512 22720
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6104 21146 6132 21678
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6564 21486 6592 21966
rect 6552 21480 6604 21486
rect 6552 21422 6604 21428
rect 6276 21412 6328 21418
rect 6276 21354 6328 21360
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5644 19718 5672 20742
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 6104 18902 6132 21082
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 5460 9178 5488 16390
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 11898 5580 14214
rect 6288 12782 6316 21354
rect 6458 19816 6514 19825
rect 6458 19751 6460 19760
rect 6512 19751 6514 19760
rect 6460 19722 6512 19728
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6380 12306 6408 17546
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5644 11218 5672 12174
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 9874 5580 11018
rect 5644 10674 5672 11154
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5644 9994 5672 10610
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5552 9846 5672 9874
rect 5644 9382 5672 9846
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 5368 7886 5396 8910
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 1766 6216 1822 6225
rect 1766 6151 1768 6160
rect 1820 6151 1822 6160
rect 1768 6122 1820 6128
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5846 2452 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 4632 5710 4660 7142
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4865 1808 4966
rect 1766 4856 1822 4865
rect 1766 4791 1822 4800
rect 2792 3738 2820 5578
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 20 2848 72 2854
rect 1780 2825 1808 3470
rect 2884 3126 2912 5510
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 20 2790 72 2796
rect 1766 2816 1822 2825
rect 32 800 60 2790
rect 1766 2751 1822 2760
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 2608 800 2636 2382
rect 2792 1465 2820 2994
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4724 2650 4752 6734
rect 5552 6390 5580 7142
rect 5644 6730 5672 9318
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4816 2582 4844 6054
rect 5736 5681 5764 11018
rect 5828 7954 5856 11834
rect 6380 11558 6408 12242
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6012 8838 6040 9522
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6012 7002 6040 7346
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5998 6896 6054 6905
rect 5998 6831 6054 6840
rect 6012 6798 6040 6831
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5828 6254 5856 6598
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 6288 5914 6316 9930
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9722 6408 9862
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6472 9518 6500 19722
rect 6748 19242 6776 23530
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7392 22642 7420 23258
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7484 21350 7512 30058
rect 7748 29640 7800 29646
rect 7748 29582 7800 29588
rect 7564 29504 7616 29510
rect 7564 29446 7616 29452
rect 7576 24818 7604 29446
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7760 24206 7788 29582
rect 8588 29238 8616 30262
rect 9128 29844 9180 29850
rect 9128 29786 9180 29792
rect 9140 29646 9168 29786
rect 9128 29640 9180 29646
rect 9128 29582 9180 29588
rect 9140 29306 9168 29582
rect 9128 29300 9180 29306
rect 9128 29242 9180 29248
rect 8576 29232 8628 29238
rect 8576 29174 8628 29180
rect 8208 29096 8260 29102
rect 8208 29038 8260 29044
rect 8220 28490 8248 29038
rect 8208 28484 8260 28490
rect 8208 28426 8260 28432
rect 8300 26784 8352 26790
rect 8300 26726 8352 26732
rect 8312 26450 8340 26726
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8208 25968 8260 25974
rect 8208 25910 8260 25916
rect 8220 25294 8248 25910
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 7748 24200 7800 24206
rect 7748 24142 7800 24148
rect 7760 23730 7788 24142
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 7760 22642 7788 23666
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7760 22438 7788 22578
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7472 21344 7524 21350
rect 7472 21286 7524 21292
rect 6736 19236 6788 19242
rect 6736 19178 6788 19184
rect 7576 18698 7604 22374
rect 7852 21962 7880 23462
rect 8220 22642 8248 25230
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 7840 21956 7892 21962
rect 7840 21898 7892 21904
rect 7932 20800 7984 20806
rect 7932 20742 7984 20748
rect 7838 20632 7894 20641
rect 7838 20567 7894 20576
rect 7852 20534 7880 20567
rect 7840 20528 7892 20534
rect 7840 20470 7892 20476
rect 7944 19854 7972 20742
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 6840 18426 6868 18634
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6748 9178 6776 11766
rect 6840 11762 6868 12718
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 9178 6868 11494
rect 6932 9382 6960 11698
rect 7300 10606 7328 18022
rect 7944 17270 7972 19790
rect 8312 18970 8340 22170
rect 8588 22098 8616 29174
rect 9232 28626 9260 31826
rect 10152 31414 10180 32166
rect 10428 31822 10456 37062
rect 11244 32768 11296 32774
rect 11244 32710 11296 32716
rect 11152 32428 11204 32434
rect 11152 32370 11204 32376
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 10876 31816 10928 31822
rect 10876 31758 10928 31764
rect 10600 31748 10652 31754
rect 10600 31690 10652 31696
rect 10140 31408 10192 31414
rect 10140 31350 10192 31356
rect 9588 31204 9640 31210
rect 9588 31146 9640 31152
rect 9404 30728 9456 30734
rect 9404 30670 9456 30676
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 9324 29714 9352 29990
rect 9312 29708 9364 29714
rect 9312 29650 9364 29656
rect 9220 28620 9272 28626
rect 9220 28562 9272 28568
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9140 26450 9168 27406
rect 9312 26852 9364 26858
rect 9312 26794 9364 26800
rect 9128 26444 9180 26450
rect 9128 26386 9180 26392
rect 9036 26036 9088 26042
rect 9036 25978 9088 25984
rect 9048 25226 9076 25978
rect 9140 25362 9168 26386
rect 9324 26382 9352 26794
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9128 25356 9180 25362
rect 9128 25298 9180 25304
rect 9036 25220 9088 25226
rect 9036 25162 9088 25168
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7576 12986 7604 16390
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7760 14618 7788 14894
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7944 12238 7972 17206
rect 8404 16794 8432 19110
rect 9048 18970 9076 25162
rect 9140 22710 9168 25298
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 9416 22094 9444 30670
rect 9600 30394 9628 31146
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10428 30802 10456 31078
rect 10416 30796 10468 30802
rect 10416 30738 10468 30744
rect 10612 30734 10640 31690
rect 10692 31340 10744 31346
rect 10692 31282 10744 31288
rect 10704 30938 10732 31282
rect 10692 30932 10744 30938
rect 10692 30874 10744 30880
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9496 30320 9548 30326
rect 9496 30262 9548 30268
rect 9508 30054 9536 30262
rect 9496 30048 9548 30054
rect 9496 29990 9548 29996
rect 9600 28150 9628 30330
rect 9864 29164 9916 29170
rect 9864 29106 9916 29112
rect 9876 28558 9904 29106
rect 9864 28552 9916 28558
rect 9864 28494 9916 28500
rect 9588 28144 9640 28150
rect 9588 28086 9640 28092
rect 10048 26920 10100 26926
rect 10046 26888 10048 26897
rect 10100 26888 10102 26897
rect 10046 26823 10102 26832
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9784 24750 9812 26182
rect 10060 25906 10088 26823
rect 10048 25900 10100 25906
rect 10048 25842 10100 25848
rect 9772 24744 9824 24750
rect 9772 24686 9824 24692
rect 10152 23594 10180 30670
rect 10888 30326 10916 31758
rect 11164 31686 11192 32370
rect 11152 31680 11204 31686
rect 11152 31622 11204 31628
rect 11060 31272 11112 31278
rect 11060 31214 11112 31220
rect 10876 30320 10928 30326
rect 10876 30262 10928 30268
rect 10692 30252 10744 30258
rect 10692 30194 10744 30200
rect 10508 29504 10560 29510
rect 10508 29446 10560 29452
rect 10520 29102 10548 29446
rect 10600 29232 10652 29238
rect 10600 29174 10652 29180
rect 10508 29096 10560 29102
rect 10508 29038 10560 29044
rect 10612 28762 10640 29174
rect 10704 29102 10732 30194
rect 11072 30122 11100 31214
rect 11164 30870 11192 31622
rect 11152 30864 11204 30870
rect 11152 30806 11204 30812
rect 11152 30660 11204 30666
rect 11152 30602 11204 30608
rect 11060 30116 11112 30122
rect 11060 30058 11112 30064
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 10600 28756 10652 28762
rect 10600 28698 10652 28704
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 10140 23588 10192 23594
rect 10140 23530 10192 23536
rect 10612 23526 10640 25774
rect 10704 23798 10732 29038
rect 10876 28552 10928 28558
rect 10876 28494 10928 28500
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10796 26382 10824 26726
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10888 25158 10916 28494
rect 11164 27062 11192 30602
rect 11256 29646 11284 32710
rect 11336 30184 11388 30190
rect 11336 30126 11388 30132
rect 11244 29640 11296 29646
rect 11244 29582 11296 29588
rect 11348 29170 11376 30126
rect 11716 30122 11744 37062
rect 11796 33312 11848 33318
rect 11796 33254 11848 33260
rect 11808 32434 11836 33254
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11888 32224 11940 32230
rect 11888 32166 11940 32172
rect 11704 30116 11756 30122
rect 11704 30058 11756 30064
rect 11520 30048 11572 30054
rect 11520 29990 11572 29996
rect 11532 29714 11560 29990
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 11520 29572 11572 29578
rect 11520 29514 11572 29520
rect 11336 29164 11388 29170
rect 11336 29106 11388 29112
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 11152 27056 11204 27062
rect 11152 26998 11204 27004
rect 10980 25430 11008 26998
rect 11428 26308 11480 26314
rect 11428 26250 11480 26256
rect 11440 26042 11468 26250
rect 11428 26036 11480 26042
rect 11428 25978 11480 25984
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 10968 25424 11020 25430
rect 10968 25366 11020 25372
rect 10876 25152 10928 25158
rect 10876 25094 10928 25100
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10692 23792 10744 23798
rect 10692 23734 10744 23740
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 9586 23352 9642 23361
rect 9586 23287 9642 23296
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9232 22066 9444 22094
rect 9508 22094 9536 22374
rect 9600 22234 9628 23287
rect 10612 22642 10640 23462
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9508 22066 9628 22094
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 9048 17796 9076 18906
rect 9232 18154 9260 22066
rect 9600 22030 9628 22066
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9496 21956 9548 21962
rect 9496 21898 9548 21904
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9416 21622 9444 21830
rect 9404 21616 9456 21622
rect 9404 21558 9456 21564
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9324 19310 9352 20334
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 8496 17768 9076 17796
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6656 8362 6684 8570
rect 6840 8498 6868 8910
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 6736 6792 6788 6798
rect 7208 6746 7236 6938
rect 7392 6798 7420 11630
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 7576 8906 7604 10678
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7852 7002 7880 12038
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8404 9042 8432 9454
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8566 8248 8842
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 6736 6734 6788 6740
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 5722 5672 5778 5681
rect 5722 5607 5778 5616
rect 6472 5234 6500 6598
rect 6748 6458 6776 6734
rect 7116 6718 7236 6746
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 3534 6684 4966
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 6564 2446 6592 3334
rect 7116 2514 7144 6718
rect 7392 6662 7420 6734
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7208 6322 7236 6598
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7208 5846 7236 6122
rect 7760 6118 7788 6326
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7392 5302 7420 6054
rect 7852 5914 7880 6326
rect 7944 5914 7972 6598
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8312 5778 8340 8434
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8496 5710 8524 17768
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8668 17264 8720 17270
rect 8668 17206 8720 17212
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8588 10266 8616 12582
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8680 8090 8708 17206
rect 8956 17134 8984 17614
rect 9232 17338 9260 18090
rect 9324 17338 9352 19246
rect 9416 17610 9444 21422
rect 9508 20942 9536 21898
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9508 19922 9536 20878
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8772 10810 8800 16730
rect 8956 16590 8984 17070
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8956 16114 8984 16526
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8956 14482 8984 16050
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 9232 14278 9260 15982
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9232 11286 9260 14214
rect 9416 13394 9444 14418
rect 9508 14074 9536 14894
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9508 13938 9536 14010
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 12170 9352 12582
rect 9600 12434 9628 21966
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9692 20874 9720 21830
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 10796 19514 10824 24006
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 16590 10364 18702
rect 10888 18698 10916 25094
rect 11164 23254 11192 25638
rect 11152 23248 11204 23254
rect 11152 23190 11204 23196
rect 11058 22128 11114 22137
rect 11058 22063 11114 22072
rect 11072 21962 11100 22063
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 11072 20058 11100 21898
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11164 19786 11192 21830
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11440 19446 11468 19926
rect 11532 19854 11560 29514
rect 11900 27402 11928 32166
rect 11992 32026 12020 37198
rect 12912 37126 12940 39200
rect 14844 37262 14872 39200
rect 16132 37262 16160 39200
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 16120 37256 16172 37262
rect 16120 37198 16172 37204
rect 17224 37256 17276 37262
rect 17224 37198 17276 37204
rect 12900 37120 12952 37126
rect 12900 37062 12952 37068
rect 14740 37120 14792 37126
rect 14740 37062 14792 37068
rect 16580 37120 16632 37126
rect 16580 37062 16632 37068
rect 12164 34060 12216 34066
rect 12164 34002 12216 34008
rect 12176 33522 12204 34002
rect 12624 33856 12676 33862
rect 12624 33798 12676 33804
rect 13544 33856 13596 33862
rect 13544 33798 13596 33804
rect 12636 33590 12664 33798
rect 12624 33584 12676 33590
rect 12624 33526 12676 33532
rect 13556 33522 13584 33798
rect 12164 33516 12216 33522
rect 12164 33458 12216 33464
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 11980 32020 12032 32026
rect 11980 31962 12032 31968
rect 12176 31754 12204 33458
rect 13912 33312 13964 33318
rect 13912 33254 13964 33260
rect 13360 32904 13412 32910
rect 13360 32846 13412 32852
rect 12992 31816 13044 31822
rect 12992 31758 13044 31764
rect 12176 31726 12296 31754
rect 12072 31136 12124 31142
rect 12072 31078 12124 31084
rect 12084 29510 12112 31078
rect 12072 29504 12124 29510
rect 12072 29446 12124 29452
rect 11888 27396 11940 27402
rect 11888 27338 11940 27344
rect 12164 27328 12216 27334
rect 12164 27270 12216 27276
rect 12176 26314 12204 27270
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 11704 25832 11756 25838
rect 11704 25774 11756 25780
rect 11716 24818 11744 25774
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 11808 22438 11836 22986
rect 12164 22500 12216 22506
rect 12164 22442 12216 22448
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 12176 21146 12204 22442
rect 12268 21622 12296 31726
rect 13004 30938 13032 31758
rect 13084 31136 13136 31142
rect 13084 31078 13136 31084
rect 12992 30932 13044 30938
rect 12992 30874 13044 30880
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 12360 29306 12388 30194
rect 12992 29708 13044 29714
rect 12992 29650 13044 29656
rect 12808 29572 12860 29578
rect 12808 29514 12860 29520
rect 12820 29306 12848 29514
rect 12348 29300 12400 29306
rect 12348 29242 12400 29248
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 12808 29300 12860 29306
rect 12808 29242 12860 29248
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 12452 27554 12480 29106
rect 12360 27526 12480 27554
rect 12360 26042 12388 27526
rect 12544 27062 12572 29242
rect 13004 29102 13032 29650
rect 12992 29096 13044 29102
rect 12992 29038 13044 29044
rect 13004 28626 13032 29038
rect 12992 28620 13044 28626
rect 12992 28562 13044 28568
rect 12808 27328 12860 27334
rect 13096 27282 13124 31078
rect 13372 30870 13400 32846
rect 13924 32570 13952 33254
rect 13912 32564 13964 32570
rect 13912 32506 13964 32512
rect 14752 32434 14780 37062
rect 15292 34604 15344 34610
rect 15292 34546 15344 34552
rect 15304 33318 15332 34546
rect 15292 33312 15344 33318
rect 15292 33254 15344 33260
rect 15384 32768 15436 32774
rect 15384 32710 15436 32716
rect 15660 32768 15712 32774
rect 15660 32710 15712 32716
rect 15396 32502 15424 32710
rect 15384 32496 15436 32502
rect 15384 32438 15436 32444
rect 15672 32434 15700 32710
rect 13452 32428 13504 32434
rect 13452 32370 13504 32376
rect 14188 32428 14240 32434
rect 14188 32370 14240 32376
rect 14740 32428 14792 32434
rect 14740 32370 14792 32376
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 16396 32428 16448 32434
rect 16396 32370 16448 32376
rect 13464 31482 13492 32370
rect 14004 32224 14056 32230
rect 14004 32166 14056 32172
rect 14096 32224 14148 32230
rect 14096 32166 14148 32172
rect 13636 31952 13688 31958
rect 13636 31894 13688 31900
rect 13452 31476 13504 31482
rect 13452 31418 13504 31424
rect 13648 31346 13676 31894
rect 14016 31822 14044 32166
rect 14004 31816 14056 31822
rect 14004 31758 14056 31764
rect 13636 31340 13688 31346
rect 13636 31282 13688 31288
rect 13728 31136 13780 31142
rect 13728 31078 13780 31084
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13740 30938 13768 31078
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 13360 30864 13412 30870
rect 13360 30806 13412 30812
rect 13372 30734 13400 30806
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 13176 30048 13228 30054
rect 13176 29990 13228 29996
rect 13188 29170 13216 29990
rect 13176 29164 13228 29170
rect 13176 29106 13228 29112
rect 13728 27668 13780 27674
rect 13728 27610 13780 27616
rect 12808 27270 12860 27276
rect 12714 27160 12770 27169
rect 12714 27095 12716 27104
rect 12768 27095 12770 27104
rect 12716 27066 12768 27072
rect 12532 27056 12584 27062
rect 12452 27004 12532 27010
rect 12452 26998 12584 27004
rect 12452 26982 12572 26998
rect 12820 26994 12848 27270
rect 12912 27254 13124 27282
rect 12808 26988 12860 26994
rect 12348 26036 12400 26042
rect 12348 25978 12400 25984
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11808 19446 11836 19654
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11796 19440 11848 19446
rect 11796 19382 11848 19388
rect 12256 19304 12308 19310
rect 12360 19292 12388 23598
rect 12308 19264 12388 19292
rect 12256 19246 12308 19252
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10336 15570 10364 16526
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14346 9720 14758
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10336 14006 10364 14214
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9416 12406 9628 12434
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9416 10810 9444 12406
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 9048 8090 9076 9590
rect 9416 8498 9444 10746
rect 9600 8566 9628 11630
rect 9784 11150 9812 13330
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 9722 9720 10406
rect 9784 10062 9812 11086
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9784 9722 9812 9998
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 10060 9382 10088 13330
rect 10520 13258 10548 15098
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10612 12434 10640 15846
rect 10612 12406 10732 12434
rect 10704 11898 10732 12406
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 10152 8430 10180 9930
rect 10796 9654 10824 17818
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10980 15570 11008 15982
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 11164 14618 11192 16594
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11348 14618 11376 16118
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10980 12918 11008 14486
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11440 13258 11468 14282
rect 11532 13530 11560 18566
rect 12164 15088 12216 15094
rect 12164 15030 12216 15036
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 11624 12850 11652 14350
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 12176 12442 12204 15030
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11624 11286 11652 11494
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11808 11150 11836 11494
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11440 10062 11468 10542
rect 11532 10198 11560 10950
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 10784 9648 10836 9654
rect 10782 9616 10784 9625
rect 10836 9616 10838 9625
rect 10782 9551 10838 9560
rect 11532 9382 11560 10134
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11808 9110 11836 11086
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 9518 12020 9862
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11992 8838 12020 9454
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9232 6866 9260 7278
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9784 6390 9812 7822
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10336 7478 10364 7686
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 9876 6866 9904 7414
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 10796 6458 10824 7210
rect 10980 6934 11008 7686
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 10152 5234 10180 6258
rect 11532 5574 11560 8774
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11624 6186 11652 6802
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11716 5846 11744 6734
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7300 3194 7328 5102
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 8312 2446 8340 2858
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9140 2446 9168 2790
rect 10152 2582 10180 5170
rect 11992 5166 12020 7278
rect 12268 6914 12296 19246
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12360 18426 12388 18634
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12452 17814 12480 26982
rect 12808 26930 12860 26936
rect 12912 26314 12940 27254
rect 13740 26926 13768 27610
rect 12992 26920 13044 26926
rect 13268 26920 13320 26926
rect 13044 26868 13216 26874
rect 12992 26862 13216 26868
rect 13268 26862 13320 26868
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13004 26846 13216 26862
rect 13188 26450 13216 26846
rect 13176 26444 13228 26450
rect 13176 26386 13228 26392
rect 12900 26308 12952 26314
rect 12900 26250 12952 26256
rect 13188 24750 13216 26386
rect 13176 24744 13228 24750
rect 13176 24686 13228 24692
rect 12992 24676 13044 24682
rect 12992 24618 13044 24624
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12544 21622 12572 21898
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12912 20398 12940 22034
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12912 19310 12940 20334
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12912 18222 12940 19246
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12912 17134 12940 18158
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12912 16046 12940 17070
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12346 13288 12402 13297
rect 12346 13223 12402 13232
rect 12360 12986 12388 13223
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12636 12374 12664 14826
rect 12820 13530 12848 15370
rect 12912 14958 12940 15982
rect 13004 15434 13032 24618
rect 13188 23662 13216 24686
rect 13176 23656 13228 23662
rect 13176 23598 13228 23604
rect 13188 23186 13216 23598
rect 13280 23186 13308 26862
rect 13832 26790 13860 31078
rect 14108 30410 14136 32166
rect 14016 30382 14136 30410
rect 13912 30048 13964 30054
rect 13912 29990 13964 29996
rect 13924 28150 13952 29990
rect 13912 28144 13964 28150
rect 13912 28086 13964 28092
rect 14016 27334 14044 30382
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 14108 29170 14136 30194
rect 14200 30190 14228 32370
rect 16028 32224 16080 32230
rect 16028 32166 16080 32172
rect 16040 32026 16068 32166
rect 16028 32020 16080 32026
rect 16028 31962 16080 31968
rect 15752 31952 15804 31958
rect 15752 31894 15804 31900
rect 15568 31272 15620 31278
rect 15568 31214 15620 31220
rect 14556 31204 14608 31210
rect 14556 31146 14608 31152
rect 14568 30666 14596 31146
rect 15580 30802 15608 31214
rect 15660 30932 15712 30938
rect 15660 30874 15712 30880
rect 15568 30796 15620 30802
rect 15568 30738 15620 30744
rect 14464 30660 14516 30666
rect 14464 30602 14516 30608
rect 14556 30660 14608 30666
rect 14556 30602 14608 30608
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 14280 30116 14332 30122
rect 14280 30058 14332 30064
rect 14292 29646 14320 30058
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14372 29504 14424 29510
rect 14372 29446 14424 29452
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14004 27328 14056 27334
rect 14004 27270 14056 27276
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13740 24410 13768 25434
rect 13636 24404 13688 24410
rect 13636 24346 13688 24352
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 13648 23866 13676 24346
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13176 23180 13228 23186
rect 13176 23122 13228 23128
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13188 22098 13216 23122
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13832 21554 13860 22986
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13464 20534 13492 20742
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 13372 18902 13400 19382
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13188 15706 13216 18158
rect 13556 17270 13584 21490
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13648 17134 13676 17478
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13280 16182 13308 16458
rect 13268 16176 13320 16182
rect 13268 16118 13320 16124
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12912 12782 12940 14894
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 12918 13400 13126
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13464 12782 13492 13262
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 12624 12368 12676 12374
rect 12624 12310 12676 12316
rect 12636 12238 12664 12310
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12532 11688 12584 11694
rect 12360 11636 12532 11642
rect 12360 11630 12584 11636
rect 12360 11614 12572 11630
rect 12360 10130 12388 11614
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12084 6886 12296 6914
rect 12084 6254 12112 6886
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6322 12204 6598
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4146 11192 4422
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 3058 11100 3334
rect 11808 3126 11836 4966
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4146 11928 4422
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11164 2650 11192 2994
rect 11992 2922 12020 5102
rect 12084 4622 12112 6054
rect 12268 5914 12296 6734
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12360 5234 12388 5850
rect 12452 5846 12480 6190
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12544 5642 12572 9590
rect 12636 7886 12664 12174
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12636 7410 12664 7822
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12820 5642 12848 12038
rect 12912 11898 12940 12718
rect 13464 12238 13492 12718
rect 13648 12434 13676 17070
rect 13832 14346 13860 21490
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13924 20058 13952 21286
rect 14108 21010 14136 29106
rect 14384 28014 14412 29446
rect 14476 29306 14504 30602
rect 14464 29300 14516 29306
rect 14464 29242 14516 29248
rect 15016 28960 15068 28966
rect 15016 28902 15068 28908
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 14476 28150 14504 28494
rect 14832 28484 14884 28490
rect 14832 28426 14884 28432
rect 14844 28218 14872 28426
rect 14832 28212 14884 28218
rect 14832 28154 14884 28160
rect 14464 28144 14516 28150
rect 14464 28086 14516 28092
rect 15028 28082 15056 28902
rect 15672 28626 15700 30874
rect 15764 30802 15792 31894
rect 16408 31822 16436 32370
rect 16396 31816 16448 31822
rect 16396 31758 16448 31764
rect 16408 31634 16436 31758
rect 16316 31606 16436 31634
rect 15752 30796 15804 30802
rect 15752 30738 15804 30744
rect 16028 28960 16080 28966
rect 16028 28902 16080 28908
rect 16040 28626 16068 28902
rect 15660 28620 15712 28626
rect 15660 28562 15712 28568
rect 16028 28620 16080 28626
rect 16028 28562 16080 28568
rect 15016 28076 15068 28082
rect 15016 28018 15068 28024
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14648 27532 14700 27538
rect 14648 27474 14700 27480
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14568 26926 14596 27066
rect 14556 26920 14608 26926
rect 14556 26862 14608 26868
rect 14568 26450 14596 26862
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14660 25974 14688 27474
rect 14924 27396 14976 27402
rect 14924 27338 14976 27344
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 14372 25968 14424 25974
rect 14372 25910 14424 25916
rect 14648 25968 14700 25974
rect 14648 25910 14700 25916
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 14108 19514 14136 20946
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13924 18834 13952 19246
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 14200 16046 14228 20402
rect 14384 19786 14412 25910
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14568 23118 14596 24006
rect 14752 23610 14780 26726
rect 14844 25226 14872 26726
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14936 23798 14964 27338
rect 15580 27169 15608 28018
rect 15566 27160 15622 27169
rect 15566 27095 15622 27104
rect 15016 26308 15068 26314
rect 15016 26250 15068 26256
rect 15028 26042 15056 26250
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 14924 23792 14976 23798
rect 14924 23734 14976 23740
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 14660 23582 14780 23610
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14476 21554 14504 21898
rect 14568 21690 14596 21898
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14292 15706 14320 16050
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 14016 13870 14044 14894
rect 14476 14414 14504 21490
rect 14660 21350 14688 23582
rect 14844 23474 14872 23598
rect 15016 23520 15068 23526
rect 14752 23468 15016 23474
rect 14752 23462 15068 23468
rect 14752 23446 15056 23462
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14660 20641 14688 21286
rect 14646 20632 14702 20641
rect 14752 20602 14780 23446
rect 15120 22094 15148 23666
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 14844 22066 15148 22094
rect 14844 21554 14872 22066
rect 15212 21894 15240 23462
rect 15304 23118 15332 24142
rect 15580 24070 15608 27095
rect 15672 24682 15700 28562
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15764 27878 15792 28358
rect 15856 28082 15884 28494
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15660 24676 15712 24682
rect 15660 24618 15712 24624
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15304 22642 15332 23054
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 14646 20567 14702 20576
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14936 19922 14964 21082
rect 15304 20942 15332 22578
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15212 20058 15240 20402
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 14924 19916 14976 19922
rect 14924 19858 14976 19864
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 14924 18352 14976 18358
rect 14924 18294 14976 18300
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14016 13462 14044 13806
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 13556 12406 13676 12434
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 13004 7546 13032 11018
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13188 8090 13216 9318
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 13096 7410 13124 7686
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12912 5302 12940 7346
rect 13280 6390 13308 9930
rect 13556 8430 13584 12406
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13648 8430 13676 12242
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13832 11762 13860 12174
rect 14476 11830 14504 13194
rect 14568 13190 14596 18022
rect 14936 17882 14964 18294
rect 14924 17876 14976 17882
rect 14924 17818 14976 17824
rect 14924 17740 14976 17746
rect 14844 17700 14924 17728
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12170 14596 12718
rect 14660 12646 14688 16934
rect 14844 16590 14872 17700
rect 15028 17728 15056 19722
rect 14976 17700 15056 17728
rect 14924 17682 14976 17688
rect 15488 17678 15516 20878
rect 15580 20398 15608 22578
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15580 18698 15608 20198
rect 15672 19990 15700 22918
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15764 18630 15792 27814
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15476 17672 15528 17678
rect 15856 17626 15884 28018
rect 16212 27328 16264 27334
rect 16212 27270 16264 27276
rect 15936 27056 15988 27062
rect 15936 26998 15988 27004
rect 15948 24750 15976 26998
rect 16120 26852 16172 26858
rect 16120 26794 16172 26800
rect 16132 26314 16160 26794
rect 16224 26314 16252 27270
rect 16120 26308 16172 26314
rect 16120 26250 16172 26256
rect 16212 26308 16264 26314
rect 16212 26250 16264 26256
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16028 25696 16080 25702
rect 16028 25638 16080 25644
rect 16040 24818 16068 25638
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15948 24410 15976 24550
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 15948 22098 15976 24346
rect 16132 24206 16160 24754
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 16120 24064 16172 24070
rect 16120 24006 16172 24012
rect 16028 22160 16080 22166
rect 16026 22128 16028 22137
rect 16080 22128 16082 22137
rect 15936 22092 15988 22098
rect 16026 22063 16082 22072
rect 15936 22034 15988 22040
rect 16132 20942 16160 24006
rect 16224 22094 16252 25842
rect 16316 23361 16344 31606
rect 16396 31476 16448 31482
rect 16396 31418 16448 31424
rect 16408 31346 16436 31418
rect 16592 31414 16620 37062
rect 17236 33658 17264 37198
rect 18064 37126 18092 39200
rect 18972 37256 19024 37262
rect 18972 37198 19024 37204
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 17408 34536 17460 34542
rect 17408 34478 17460 34484
rect 17224 33652 17276 33658
rect 17224 33594 17276 33600
rect 17420 33522 17448 34478
rect 17408 33516 17460 33522
rect 17408 33458 17460 33464
rect 18984 32570 19012 37198
rect 19352 37126 19380 39200
rect 20640 37210 20668 39200
rect 22572 37262 22600 39200
rect 20812 37256 20864 37262
rect 20640 37182 20760 37210
rect 20812 37198 20864 37204
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 20732 37126 20760 37182
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 18972 32564 19024 32570
rect 18972 32506 19024 32512
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19340 32360 19392 32366
rect 19340 32302 19392 32308
rect 17408 32224 17460 32230
rect 17408 32166 17460 32172
rect 16948 32020 17000 32026
rect 16948 31962 17000 31968
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16580 31408 16632 31414
rect 16580 31350 16632 31356
rect 16396 31340 16448 31346
rect 16396 31282 16448 31288
rect 16408 26994 16436 31282
rect 16580 30728 16632 30734
rect 16580 30670 16632 30676
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16408 25906 16436 26930
rect 16500 26518 16528 27406
rect 16488 26512 16540 26518
rect 16488 26454 16540 26460
rect 16592 26382 16620 30670
rect 16776 30326 16804 31758
rect 16960 31414 16988 31962
rect 17420 31822 17448 32166
rect 17592 31952 17644 31958
rect 17592 31894 17644 31900
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17224 31680 17276 31686
rect 17224 31622 17276 31628
rect 17236 31414 17264 31622
rect 16948 31408 17000 31414
rect 16948 31350 17000 31356
rect 17224 31408 17276 31414
rect 17224 31350 17276 31356
rect 17604 31278 17632 31894
rect 17592 31272 17644 31278
rect 17592 31214 17644 31220
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 16764 30320 16816 30326
rect 16764 30262 16816 30268
rect 17328 29646 17356 30534
rect 17604 30326 17632 31214
rect 19352 30870 19380 32302
rect 19444 31482 19472 32370
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 20732 31482 20760 31758
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 20720 31476 20772 31482
rect 20720 31418 20772 31424
rect 20824 30938 20852 37198
rect 20996 37120 21048 37126
rect 20996 37062 21048 37068
rect 20812 30932 20864 30938
rect 20812 30874 20864 30880
rect 19340 30864 19392 30870
rect 19340 30806 19392 30812
rect 17868 30728 17920 30734
rect 17868 30670 17920 30676
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 17592 30320 17644 30326
rect 17592 30262 17644 30268
rect 17880 30258 17908 30670
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 18972 30048 19024 30054
rect 18972 29990 19024 29996
rect 17316 29640 17368 29646
rect 17316 29582 17368 29588
rect 17132 29504 17184 29510
rect 17132 29446 17184 29452
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16868 28762 16896 29106
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 17144 28082 17172 29446
rect 18984 29170 19012 29990
rect 19156 29640 19208 29646
rect 19156 29582 19208 29588
rect 18972 29164 19024 29170
rect 18972 29106 19024 29112
rect 19168 29034 19196 29582
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 17592 28688 17644 28694
rect 17592 28630 17644 28636
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 16764 28008 16816 28014
rect 16764 27950 16816 27956
rect 16580 26376 16632 26382
rect 16580 26318 16632 26324
rect 16396 25900 16448 25906
rect 16396 25842 16448 25848
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16408 24206 16436 25230
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16408 23730 16436 24142
rect 16396 23724 16448 23730
rect 16396 23666 16448 23672
rect 16776 23662 16804 27950
rect 17040 27940 17092 27946
rect 17040 27882 17092 27888
rect 17052 27470 17080 27882
rect 17408 27872 17460 27878
rect 17408 27814 17460 27820
rect 17420 27538 17448 27814
rect 17408 27532 17460 27538
rect 17408 27474 17460 27480
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 16856 27328 16908 27334
rect 16856 27270 16908 27276
rect 16868 25974 16896 27270
rect 17316 26920 17368 26926
rect 17408 26920 17460 26926
rect 17316 26862 17368 26868
rect 17406 26888 17408 26897
rect 17460 26888 17462 26897
rect 17328 26450 17356 26862
rect 17406 26823 17462 26832
rect 17604 26450 17632 28630
rect 19168 28218 19196 28970
rect 19432 28484 19484 28490
rect 19432 28426 19484 28432
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19156 28212 19208 28218
rect 19156 28154 19208 28160
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18156 27538 18184 27950
rect 19352 27606 19380 28358
rect 19444 28218 19472 28426
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19432 28212 19484 28218
rect 19432 28154 19484 28160
rect 19996 28082 20024 30670
rect 20168 30592 20220 30598
rect 20168 30534 20220 30540
rect 20180 29714 20208 30534
rect 20456 29850 20484 30670
rect 20444 29844 20496 29850
rect 20444 29786 20496 29792
rect 20168 29708 20220 29714
rect 20168 29650 20220 29656
rect 21008 29646 21036 37062
rect 23308 33658 23336 37198
rect 23756 37188 23808 37194
rect 23756 37130 23808 37136
rect 23296 33652 23348 33658
rect 23296 33594 23348 33600
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 21364 31884 21416 31890
rect 21364 31826 21416 31832
rect 21376 31346 21404 31826
rect 21364 31340 21416 31346
rect 21364 31282 21416 31288
rect 22468 31340 22520 31346
rect 22468 31282 22520 31288
rect 21376 29850 21404 31282
rect 22480 30258 22508 31282
rect 22848 30938 22876 33458
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 23308 32570 23336 32846
rect 23296 32564 23348 32570
rect 23296 32506 23348 32512
rect 22928 31816 22980 31822
rect 22928 31758 22980 31764
rect 22940 31482 22968 31758
rect 22928 31476 22980 31482
rect 22928 31418 22980 31424
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 22744 30728 22796 30734
rect 22744 30670 22796 30676
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 21640 30048 21692 30054
rect 21640 29990 21692 29996
rect 21364 29844 21416 29850
rect 21364 29786 21416 29792
rect 21652 29714 21680 29990
rect 21640 29708 21692 29714
rect 21640 29650 21692 29656
rect 20628 29640 20680 29646
rect 20628 29582 20680 29588
rect 20996 29640 21048 29646
rect 20996 29582 21048 29588
rect 20076 29504 20128 29510
rect 20076 29446 20128 29452
rect 20088 29102 20116 29446
rect 20076 29096 20128 29102
rect 20076 29038 20128 29044
rect 20088 28762 20116 29038
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 20536 28144 20588 28150
rect 20536 28086 20588 28092
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 19444 27674 19472 28018
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 18144 27532 18196 27538
rect 18144 27474 18196 27480
rect 19444 26994 19472 27610
rect 20548 27606 20576 28086
rect 19984 27600 20036 27606
rect 19984 27542 20036 27548
rect 20536 27600 20588 27606
rect 20536 27542 20588 27548
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19616 26784 19668 26790
rect 19616 26726 19668 26732
rect 18696 26512 18748 26518
rect 18696 26454 18748 26460
rect 19432 26512 19484 26518
rect 19432 26454 19484 26460
rect 17316 26444 17368 26450
rect 17316 26386 17368 26392
rect 17592 26444 17644 26450
rect 17592 26386 17644 26392
rect 16856 25968 16908 25974
rect 16856 25910 16908 25916
rect 17604 25770 17632 26386
rect 18512 25832 18564 25838
rect 18512 25774 18564 25780
rect 17592 25764 17644 25770
rect 17592 25706 17644 25712
rect 17224 24880 17276 24886
rect 17224 24822 17276 24828
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 16302 23352 16358 23361
rect 16302 23287 16358 23296
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16488 23044 16540 23050
rect 16488 22986 16540 22992
rect 16500 22778 16528 22986
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 16224 22066 16344 22094
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 16316 20602 16344 22066
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16408 21146 16436 21898
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15476 17614 15528 17620
rect 15488 16658 15516 17614
rect 15580 17598 15884 17626
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14844 15502 14872 16526
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15396 16250 15424 16390
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14752 13870 14780 14350
rect 14844 14278 14872 15438
rect 15120 14890 15148 15982
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13740 9926 13768 11154
rect 13832 10674 13860 11698
rect 14568 11626 14596 12106
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13832 9586 13860 10610
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13556 5846 13584 6666
rect 13740 6254 13768 9454
rect 13832 8566 13860 9522
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 14016 6458 14044 10678
rect 14108 10606 14136 11222
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14108 9042 14136 10542
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14108 6914 14136 8978
rect 14660 8090 14688 12582
rect 14752 11898 14780 12854
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14844 10606 14872 14214
rect 15028 13326 15056 14418
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14936 9654 14964 12038
rect 15028 11762 15056 13262
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15120 11286 15148 13874
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15212 12170 15240 13126
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15304 12306 15332 12786
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15292 12096 15344 12102
rect 15212 12044 15292 12050
rect 15212 12038 15344 12044
rect 15212 12022 15332 12038
rect 15108 11280 15160 11286
rect 15108 11222 15160 11228
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15028 10810 15056 11086
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15028 10130 15056 10746
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 15108 9104 15160 9110
rect 15212 9092 15240 12022
rect 15396 11558 15424 15302
rect 15488 14482 15516 16594
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15580 13394 15608 17598
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15856 17270 15884 17478
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 15948 15502 15976 20334
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15660 13320 15712 13326
rect 15658 13288 15660 13297
rect 15712 13288 15714 13297
rect 15658 13223 15714 13232
rect 15672 11880 15700 13223
rect 15764 12850 15792 13874
rect 16040 12918 16068 20538
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16132 19825 16160 20402
rect 16118 19816 16174 19825
rect 16118 19751 16174 19760
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15764 12730 15792 12786
rect 15764 12702 15884 12730
rect 16040 12714 16068 12854
rect 15672 11852 15792 11880
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15304 9110 15332 11494
rect 15672 11150 15700 11698
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15764 10674 15792 11852
rect 15856 11150 15884 12702
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15160 9064 15240 9092
rect 15292 9104 15344 9110
rect 15108 9046 15160 9052
rect 15292 9046 15344 9052
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15108 8968 15160 8974
rect 15396 8956 15424 9046
rect 15160 8928 15424 8956
rect 15108 8910 15160 8916
rect 15488 8498 15516 10202
rect 15580 9450 15608 10406
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15764 8974 15792 9590
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15844 9376 15896 9382
rect 15842 9344 15844 9353
rect 15896 9344 15898 9353
rect 15842 9279 15898 9288
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15948 8906 15976 9522
rect 16040 9382 16068 11494
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16026 9208 16082 9217
rect 16026 9143 16082 9152
rect 16040 9042 16068 9143
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 14476 7546 14504 7754
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14108 6886 14228 6914
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12360 4282 12388 5170
rect 13740 4622 13768 6190
rect 14200 5778 14228 6886
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5778 14504 6054
rect 14568 5778 14596 6598
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14936 5710 14964 6258
rect 15120 6186 15148 7754
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15488 7002 15516 7686
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15672 6458 15700 6734
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15764 6390 15792 8298
rect 16040 8294 16068 8434
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16132 6798 16160 19751
rect 16500 18698 16528 20742
rect 16684 19174 16712 21830
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16488 18692 16540 18698
rect 16488 18634 16540 18640
rect 16684 18290 16712 19110
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16776 16726 16804 23122
rect 16960 20398 16988 23598
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16868 18834 16896 19246
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16396 16516 16448 16522
rect 16396 16458 16448 16464
rect 16408 15706 16436 16458
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16500 15586 16528 16662
rect 16960 16402 16988 20198
rect 17052 18698 17080 24618
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17144 21894 17172 23054
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 17144 21078 17172 21354
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17236 20058 17264 24822
rect 17868 24132 17920 24138
rect 17868 24074 17920 24080
rect 17880 23662 17908 24074
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 18064 23730 18092 24006
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17040 18692 17092 18698
rect 17040 18634 17092 18640
rect 16408 15558 16528 15586
rect 16868 16374 16988 16402
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16316 13938 16344 14350
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16224 11898 16252 12378
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16212 10736 16264 10742
rect 16212 10678 16264 10684
rect 16224 9994 16252 10678
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 16408 9110 16436 15558
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16500 12238 16528 13806
rect 16592 12442 16620 15030
rect 16764 14544 16816 14550
rect 16764 14486 16816 14492
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16500 11830 16528 12174
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16684 11218 16712 14282
rect 16776 14006 16804 14486
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16500 10742 16528 11086
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8294 16528 8774
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16488 8288 16540 8294
rect 16488 8230 16540 8236
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 6798 16344 7142
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 16408 6322 16436 8230
rect 16592 6914 16620 10474
rect 16684 9654 16712 11154
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16684 9058 16712 9590
rect 16764 9376 16816 9382
rect 16762 9344 16764 9353
rect 16816 9344 16818 9353
rect 16762 9279 16818 9288
rect 16684 9030 16804 9058
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8294 16712 8910
rect 16776 8498 16804 9030
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16684 7818 16712 8026
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16776 7410 16804 8434
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16776 6914 16804 7346
rect 16868 7018 16896 16374
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14482 16988 14894
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16960 9586 16988 12650
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 17052 9466 17080 18634
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17236 17746 17264 18022
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17236 15706 17264 16118
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17236 13530 17264 13942
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17328 13410 17356 21490
rect 17420 20505 17448 21830
rect 17512 21690 17540 22646
rect 17776 22500 17828 22506
rect 17776 22442 17828 22448
rect 17788 22234 17816 22442
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17880 22098 17908 23462
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17972 21622 18000 23054
rect 18236 23044 18288 23050
rect 18236 22986 18288 22992
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17684 20936 17736 20942
rect 17736 20884 17816 20890
rect 17684 20878 17816 20884
rect 17696 20862 17816 20878
rect 17406 20496 17462 20505
rect 17406 20431 17462 20440
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 17420 19446 17448 20266
rect 17788 19854 17816 20862
rect 17880 20754 17908 21422
rect 18052 20800 18104 20806
rect 17880 20748 18052 20754
rect 17880 20742 18104 20748
rect 17880 20726 18092 20742
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17408 19440 17460 19446
rect 17408 19382 17460 19388
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16658 17540 16934
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17406 16552 17462 16561
rect 17406 16487 17462 16496
rect 17420 16046 17448 16487
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17512 15162 17540 16594
rect 17604 15706 17632 17070
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17604 15042 17632 15642
rect 17236 13382 17356 13410
rect 17420 15014 17632 15042
rect 17236 9625 17264 13382
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17328 12306 17356 12718
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17420 10538 17448 15014
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17604 12782 17632 13806
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17604 11762 17632 12310
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17512 11218 17540 11630
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17408 10532 17460 10538
rect 17408 10474 17460 10480
rect 17512 9926 17540 10610
rect 17604 10266 17632 11018
rect 17696 10810 17724 11154
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17408 9648 17460 9654
rect 17222 9616 17278 9625
rect 17408 9590 17460 9596
rect 17222 9551 17278 9560
rect 17224 9512 17276 9518
rect 17052 9460 17224 9466
rect 17052 9454 17276 9460
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17052 9438 17264 9454
rect 16948 9104 17000 9110
rect 16948 9046 17000 9052
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 16960 8838 16988 9046
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 16960 7546 16988 7958
rect 17052 7886 17080 9046
rect 17040 7880 17092 7886
rect 17092 7828 17264 7834
rect 17040 7822 17264 7828
rect 17052 7806 17264 7822
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16868 7002 16988 7018
rect 16868 6996 17000 7002
rect 16868 6990 16948 6996
rect 16948 6938 17000 6944
rect 17052 6934 17080 7346
rect 17040 6928 17092 6934
rect 16592 6886 16712 6914
rect 16776 6886 16896 6914
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 16578 5672 16634 5681
rect 16578 5607 16580 5616
rect 16632 5607 16634 5616
rect 16580 5578 16632 5584
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 14292 2446 14320 4966
rect 16684 3194 16712 6886
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16776 2446 16804 6598
rect 16868 5710 16896 6886
rect 17040 6870 17092 6876
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16868 3194 16896 4082
rect 16960 4010 16988 6394
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17052 3058 17080 6870
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17144 2650 17172 6258
rect 17236 3058 17264 7806
rect 17328 7342 17356 9454
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17420 7274 17448 9590
rect 17512 8974 17540 9862
rect 17788 9382 17816 19790
rect 17880 17678 17908 20726
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17972 18698 18000 20198
rect 18156 19242 18184 22510
rect 18248 22234 18276 22986
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18248 20466 18276 22170
rect 18420 21888 18472 21894
rect 18420 21830 18472 21836
rect 18432 21010 18460 21830
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 18524 20874 18552 25774
rect 18708 24206 18736 26454
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19248 25832 19300 25838
rect 19248 25774 19300 25780
rect 19260 25362 19288 25774
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19352 24954 19380 25910
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18616 21894 18644 23462
rect 18708 23118 18736 24142
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18800 23322 18828 23598
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 19444 23254 19472 26454
rect 19628 26314 19656 26726
rect 19616 26308 19668 26314
rect 19616 26250 19668 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 19536 25430 19564 25774
rect 19524 25424 19576 25430
rect 19524 25366 19576 25372
rect 19536 25265 19564 25366
rect 19522 25256 19578 25265
rect 19522 25191 19578 25200
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23848 20024 27542
rect 20260 26988 20312 26994
rect 20260 26930 20312 26936
rect 20272 25498 20300 26930
rect 20640 26450 20668 29582
rect 20812 28416 20864 28422
rect 20812 28358 20864 28364
rect 21824 28416 21876 28422
rect 21824 28358 21876 28364
rect 20824 28082 20852 28358
rect 21836 28082 21864 28358
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20824 27538 20852 27814
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 21180 27464 21232 27470
rect 21180 27406 21232 27412
rect 20732 27130 20760 27406
rect 20720 27124 20772 27130
rect 20720 27066 20772 27072
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20732 25906 20760 26862
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20824 26450 20852 26726
rect 20812 26444 20864 26450
rect 20812 26386 20864 26392
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20628 25696 20680 25702
rect 20628 25638 20680 25644
rect 20260 25492 20312 25498
rect 20260 25434 20312 25440
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20352 24268 20404 24274
rect 20352 24210 20404 24216
rect 19536 23820 20024 23848
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 18696 23112 18748 23118
rect 19536 23066 19564 23820
rect 20364 23730 20392 24210
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 19708 23520 19760 23526
rect 19708 23462 19760 23468
rect 19720 23186 19748 23462
rect 19800 23248 19852 23254
rect 19798 23216 19800 23225
rect 19852 23216 19854 23225
rect 19708 23180 19760 23186
rect 19798 23151 19854 23160
rect 19708 23122 19760 23128
rect 19812 23118 19840 23151
rect 18696 23054 18748 23060
rect 19444 23038 19564 23066
rect 19800 23112 19852 23118
rect 19800 23054 19852 23060
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 18708 22642 18736 22918
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18512 20868 18564 20874
rect 18512 20810 18564 20816
rect 18788 20868 18840 20874
rect 18788 20810 18840 20816
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17972 17270 18000 17478
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17972 16674 18000 17206
rect 17972 16646 18184 16674
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 18064 15502 18092 16526
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18064 15094 18092 15438
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17972 13530 18000 14894
rect 18156 14414 18184 16646
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18156 13326 18184 14214
rect 18248 13870 18276 17818
rect 18328 17604 18380 17610
rect 18328 17546 18380 17552
rect 18340 17338 18368 17546
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18432 12238 18460 17138
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18524 15978 18552 17002
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18512 15972 18564 15978
rect 18512 15914 18564 15920
rect 18420 12232 18472 12238
rect 18340 12192 18420 12220
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 11898 18184 12038
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17880 11082 17908 11630
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17880 9160 17908 11018
rect 18248 10810 18276 11766
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9178 18000 9998
rect 18340 9994 18368 12192
rect 18420 12174 18472 12180
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18432 11354 18460 11834
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18064 9217 18092 9318
rect 18050 9208 18106 9217
rect 17788 9132 17908 9160
rect 17960 9172 18012 9178
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17512 8566 17540 8910
rect 17696 8566 17724 8910
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 17512 6866 17540 8366
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 7886 17724 8230
rect 17788 7954 17816 9132
rect 18248 9178 18276 9590
rect 18050 9143 18106 9152
rect 18236 9172 18288 9178
rect 17960 9114 18012 9120
rect 18236 9114 18288 9120
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17880 6730 17908 7142
rect 18524 6914 18552 15914
rect 18708 15570 18736 15982
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18616 11354 18644 12854
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18432 6886 18552 6914
rect 18800 6914 18828 20810
rect 18892 17882 18920 22374
rect 19156 22024 19208 22030
rect 19156 21966 19208 21972
rect 19168 18834 19196 21966
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19260 20398 19288 21286
rect 19352 20942 19380 22918
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20534 19380 20742
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19260 19514 19288 20334
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 19168 18290 19196 18770
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 18984 16794 19012 17206
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 19260 16114 19288 19110
rect 19352 18970 19380 19382
rect 19444 19310 19472 23038
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22778 20024 23666
rect 20260 23248 20312 23254
rect 20260 23190 20312 23196
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 20088 21554 20116 22578
rect 20272 22234 20300 23190
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20180 21690 20208 21966
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19352 18154 19380 18702
rect 19996 18698 20024 20334
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18892 14006 18920 14214
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 18984 12986 19012 13942
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18892 12442 18920 12786
rect 18880 12436 18932 12442
rect 19260 12434 19288 16050
rect 19352 13870 19380 17546
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 18880 12378 18932 12384
rect 19076 12406 19288 12434
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 18984 11626 19012 11766
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18984 9042 19012 9454
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 19076 6914 19104 12406
rect 19352 11098 19380 13806
rect 19444 11257 19472 18634
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20088 18306 20116 21490
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 20180 18426 20208 18838
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 19996 18278 20116 18306
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19996 16454 20024 18278
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15026 20116 18090
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20180 15162 20208 16050
rect 20272 15570 20300 22170
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19996 13394 20024 13806
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20364 12434 20392 22646
rect 20548 22094 20576 25230
rect 20640 24818 20668 25638
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20732 24154 20760 25842
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 20824 24274 20852 24550
rect 20916 24274 20944 25230
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 21008 24818 21036 25094
rect 20996 24812 21048 24818
rect 20996 24754 21048 24760
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20732 24126 20944 24154
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20640 22642 20668 22986
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20548 22066 20668 22094
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20456 20602 20484 21422
rect 20548 20777 20576 21966
rect 20534 20768 20590 20777
rect 20534 20703 20590 20712
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20640 19394 20668 22066
rect 20732 21010 20760 23666
rect 20812 23044 20864 23050
rect 20812 22986 20864 22992
rect 20824 22166 20852 22986
rect 20812 22160 20864 22166
rect 20812 22102 20864 22108
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20548 19366 20668 19394
rect 20444 17604 20496 17610
rect 20444 17546 20496 17552
rect 20456 17338 20484 17546
rect 20548 17542 20576 19366
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20640 18834 20668 19246
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20640 17202 20668 18022
rect 20824 17814 20852 21830
rect 20916 18290 20944 24126
rect 21100 23594 21128 26930
rect 21192 25906 21220 27406
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21192 23866 21220 25842
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 21088 23588 21140 23594
rect 21088 23530 21140 23536
rect 21100 21418 21128 23530
rect 21284 22098 21312 26318
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21376 23866 21404 24006
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 21376 22778 21404 23054
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21560 21146 21588 24210
rect 21928 21622 21956 30194
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 22020 27674 22048 28494
rect 22008 27668 22060 27674
rect 22008 27610 22060 27616
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 22112 26042 22140 26318
rect 22204 26314 22232 29446
rect 22756 28218 22784 30670
rect 23584 29850 23612 30670
rect 23572 29844 23624 29850
rect 23572 29786 23624 29792
rect 23768 29646 23796 37130
rect 23860 37126 23888 39200
rect 25792 37262 25820 39200
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 27080 37126 27108 39200
rect 29012 37262 29040 39200
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 29000 37256 29052 37262
rect 30300 37244 30328 39200
rect 30380 37256 30432 37262
rect 30300 37216 30380 37244
rect 29000 37198 29052 37204
rect 31588 37244 31616 39200
rect 33520 37262 33548 39200
rect 34808 37262 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 31760 37256 31812 37262
rect 31588 37216 31760 37244
rect 30380 37198 30432 37204
rect 31760 37198 31812 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 36636 37256 36688 37262
rect 36636 37198 36688 37204
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 27172 33114 27200 37198
rect 27436 37188 27488 37194
rect 27436 37130 27488 37136
rect 27160 33108 27212 33114
rect 27160 33050 27212 33056
rect 25044 32224 25096 32230
rect 25044 32166 25096 32172
rect 23848 30796 23900 30802
rect 23848 30738 23900 30744
rect 23860 29850 23888 30738
rect 24032 30592 24084 30598
rect 24032 30534 24084 30540
rect 23848 29844 23900 29850
rect 23848 29786 23900 29792
rect 23020 29640 23072 29646
rect 23020 29582 23072 29588
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 22744 28212 22796 28218
rect 22744 28154 22796 28160
rect 22560 27124 22612 27130
rect 22560 27066 22612 27072
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 22192 26308 22244 26314
rect 22192 26250 22244 26256
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22112 23866 22140 24074
rect 22100 23860 22152 23866
rect 22100 23802 22152 23808
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22020 23050 22048 23666
rect 22204 23186 22232 26250
rect 22296 24410 22324 26318
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22388 25498 22416 25842
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22296 24188 22324 24346
rect 22296 24160 22416 24188
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22296 23662 22324 24006
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22204 21622 22232 23122
rect 22388 22030 22416 24160
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21468 20602 21496 20878
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20272 12406 20392 12434
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19430 11248 19486 11257
rect 19430 11183 19486 11192
rect 19260 11070 19380 11098
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19260 10554 19288 11070
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10742 19380 10950
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19260 10526 19380 10554
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9586 19288 9998
rect 19352 9654 19380 10526
rect 19444 10266 19472 11086
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19522 10704 19578 10713
rect 19522 10639 19578 10648
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19536 10146 19564 10639
rect 19444 10118 19564 10146
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19444 8922 19472 10118
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9654 20024 11766
rect 20272 11762 20300 12406
rect 20456 12238 20484 15914
rect 20824 14414 20852 17750
rect 20916 16114 20944 18226
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 21008 16794 21036 17070
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21100 16726 21128 17138
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 21008 16250 21036 16526
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 21100 15586 21128 16662
rect 21100 15558 21220 15586
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21008 15162 21036 15302
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 21192 15026 21220 15558
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20548 14074 20576 14282
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20916 13938 20944 14418
rect 21284 14006 21312 15370
rect 21376 14618 21404 15438
rect 21560 14890 21588 21082
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21928 20058 21956 20402
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 22020 15094 22048 17614
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 22296 16794 22324 16934
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22008 15088 22060 15094
rect 22008 15030 22060 15036
rect 21548 14884 21600 14890
rect 21548 14826 21600 14832
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21272 14000 21324 14006
rect 21272 13942 21324 13948
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 22204 13870 22232 15982
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20824 12782 20852 13126
rect 20916 12918 20944 13126
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 20824 12442 20852 12718
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20272 10742 20300 11698
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20456 10130 20484 12174
rect 21192 11082 21220 12718
rect 21744 12442 21772 13262
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21376 11694 21404 12174
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21652 11150 21680 12106
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19352 8894 19472 8922
rect 19352 7546 19380 8894
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19444 7426 19472 8774
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19444 7398 19564 7426
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19352 7018 19380 7210
rect 19260 7002 19380 7018
rect 19248 6996 19380 7002
rect 19300 6990 19380 6996
rect 19248 6938 19300 6944
rect 18800 6905 18920 6914
rect 18800 6896 18934 6905
rect 18800 6886 18878 6896
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 18052 6724 18104 6730
rect 18052 6666 18104 6672
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17420 5914 17448 6190
rect 17788 6186 17816 6666
rect 18064 6610 18092 6666
rect 17880 6582 18092 6610
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17880 5370 17908 6582
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 18432 5234 18460 6886
rect 18878 6831 18934 6840
rect 18984 6886 19104 6914
rect 18984 6322 19012 6886
rect 19260 6780 19288 6938
rect 19536 6866 19564 7398
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19260 6752 19380 6780
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19076 6322 19104 6598
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18892 5710 18920 6054
rect 19352 5846 19380 6752
rect 19444 6730 19564 6746
rect 19444 6724 19576 6730
rect 19444 6718 19524 6724
rect 19444 6458 19472 6718
rect 19524 6666 19576 6672
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 20088 6254 20116 10066
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20272 8838 20300 9862
rect 20626 9616 20682 9625
rect 20626 9551 20682 9560
rect 20640 9518 20668 9551
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20364 6458 20392 7414
rect 20548 6798 20576 9386
rect 20732 9382 20760 9454
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20824 8974 20852 9998
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 21008 8906 21036 9318
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20640 6934 20668 7278
rect 20628 6928 20680 6934
rect 20628 6870 20680 6876
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20076 6248 20128 6254
rect 20076 6190 20128 6196
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 21008 5778 21036 8842
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17604 3194 17632 3470
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 18340 3126 18368 4422
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 18616 2446 18644 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20088 2446 20116 5510
rect 21192 3466 21220 11018
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21928 8634 21956 9998
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 21916 8628 21968 8634
rect 21916 8570 21968 8576
rect 22020 7546 22048 8978
rect 22112 8906 22140 9318
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 22204 7546 22232 13806
rect 22388 12782 22416 21422
rect 22572 19854 22600 27066
rect 22756 26518 22784 28154
rect 23032 28082 23060 29582
rect 24044 29578 24072 30534
rect 24032 29572 24084 29578
rect 24032 29514 24084 29520
rect 24044 28218 24072 29514
rect 24216 29096 24268 29102
rect 24216 29038 24268 29044
rect 24228 28762 24256 29038
rect 24676 28960 24728 28966
rect 24676 28902 24728 28908
rect 24952 28960 25004 28966
rect 24952 28902 25004 28908
rect 24216 28756 24268 28762
rect 24216 28698 24268 28704
rect 24584 28620 24636 28626
rect 24584 28562 24636 28568
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 23020 28076 23072 28082
rect 23020 28018 23072 28024
rect 22928 27056 22980 27062
rect 22928 26998 22980 27004
rect 22744 26512 22796 26518
rect 22744 26454 22796 26460
rect 22940 25294 22968 26998
rect 22928 25288 22980 25294
rect 22928 25230 22980 25236
rect 22940 24818 22968 25230
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 22848 21146 22876 21558
rect 22836 21140 22888 21146
rect 22836 21082 22888 21088
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22756 19854 22784 20334
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22560 19848 22612 19854
rect 22744 19848 22796 19854
rect 22612 19796 22692 19802
rect 22560 19790 22692 19796
rect 22744 19790 22796 19796
rect 22572 19774 22692 19790
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22572 19378 22600 19654
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22664 18714 22692 19774
rect 22664 18686 22784 18714
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22480 17746 22508 18022
rect 22572 17882 22600 18158
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22664 17746 22692 18566
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22480 16998 22508 17682
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22756 16574 22784 18686
rect 22664 16546 22784 16574
rect 22664 15502 22692 16546
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22756 15706 22784 15982
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22848 14906 22876 20198
rect 22940 15434 22968 24754
rect 23032 21078 23060 28018
rect 23848 28008 23900 28014
rect 23848 27950 23900 27956
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23584 27470 23612 27814
rect 23860 27606 23888 27950
rect 24596 27674 24624 28562
rect 24688 28218 24716 28902
rect 24964 28558 24992 28902
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 24676 28212 24728 28218
rect 24676 28154 24728 28160
rect 23940 27668 23992 27674
rect 23940 27610 23992 27616
rect 24584 27668 24636 27674
rect 24584 27610 24636 27616
rect 23848 27600 23900 27606
rect 23848 27542 23900 27548
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23480 25696 23532 25702
rect 23480 25638 23532 25644
rect 23492 24818 23520 25638
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23388 24744 23440 24750
rect 23440 24692 23520 24698
rect 23388 24686 23520 24692
rect 23400 24670 23520 24686
rect 23584 24682 23612 25230
rect 23952 24750 23980 27610
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24124 26852 24176 26858
rect 24124 26794 24176 26800
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 24044 24954 24072 25094
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 24044 24750 24072 24890
rect 23940 24744 23992 24750
rect 23940 24686 23992 24692
rect 24032 24744 24084 24750
rect 24032 24686 24084 24692
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 23308 23186 23336 23598
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 23492 22114 23520 24670
rect 23572 24676 23624 24682
rect 23572 24618 23624 24624
rect 23124 22086 23520 22114
rect 24136 22098 24164 26794
rect 24504 26314 24532 26862
rect 24596 26518 24624 27270
rect 24688 26926 24716 28154
rect 25056 28082 25084 32166
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 25228 28008 25280 28014
rect 25228 27950 25280 27956
rect 25240 27674 25268 27950
rect 25228 27668 25280 27674
rect 25228 27610 25280 27616
rect 25228 27464 25280 27470
rect 25332 27452 25360 29106
rect 27160 27940 27212 27946
rect 27160 27882 27212 27888
rect 25280 27424 25360 27452
rect 25228 27406 25280 27412
rect 24768 27328 24820 27334
rect 24768 27270 24820 27276
rect 24780 27062 24808 27270
rect 25240 27130 25268 27406
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 25228 27124 25280 27130
rect 25228 27066 25280 27072
rect 24768 27056 24820 27062
rect 24768 26998 24820 27004
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 24584 26512 24636 26518
rect 24584 26454 24636 26460
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24504 25294 24532 26250
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 25320 25152 25372 25158
rect 25320 25094 25372 25100
rect 25332 24886 25360 25094
rect 25320 24880 25372 24886
rect 25320 24822 25372 24828
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25148 23730 25176 24006
rect 25136 23724 25188 23730
rect 25136 23666 25188 23672
rect 25228 23656 25280 23662
rect 25228 23598 25280 23604
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 24780 22710 24808 23190
rect 24964 23186 24992 23462
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24124 22092 24176 22098
rect 23124 21962 23152 22086
rect 24124 22034 24176 22040
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 23112 21956 23164 21962
rect 23112 21898 23164 21904
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23020 21072 23072 21078
rect 23020 21014 23072 21020
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 23032 20058 23060 20878
rect 23216 20806 23244 21898
rect 23584 21690 23612 21898
rect 24228 21690 24256 21966
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 23204 20800 23256 20806
rect 23204 20742 23256 20748
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23112 20392 23164 20398
rect 23112 20334 23164 20340
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 23124 19922 23152 20334
rect 23112 19916 23164 19922
rect 23112 19858 23164 19864
rect 23216 19802 23244 20742
rect 23584 20466 23612 20742
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23124 19774 23244 19802
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23124 16250 23152 19774
rect 23308 19666 23336 19790
rect 23216 19638 23336 19666
rect 23216 16794 23244 19638
rect 24780 18902 24808 20878
rect 24768 18896 24820 18902
rect 24768 18838 24820 18844
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24320 18358 24348 18566
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 24308 18352 24360 18358
rect 24308 18294 24360 18300
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 22756 14878 22876 14906
rect 22756 14074 22784 14878
rect 22836 14816 22888 14822
rect 22836 14758 22888 14764
rect 22848 14414 22876 14758
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22388 12102 22416 12718
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22664 11150 22692 11494
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22756 10606 22784 14010
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 23032 11626 23060 13874
rect 23112 13252 23164 13258
rect 23112 13194 23164 13200
rect 23020 11620 23072 11626
rect 23020 11562 23072 11568
rect 22836 11008 22888 11014
rect 22836 10950 22888 10956
rect 22848 10674 22876 10950
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 23124 10266 23152 13194
rect 23216 12850 23244 16730
rect 23860 16522 23888 18294
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 24228 17542 24256 18158
rect 24780 17898 24808 18838
rect 25044 18692 25096 18698
rect 25044 18634 25096 18640
rect 25056 18086 25084 18634
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 24780 17870 24900 17898
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23860 15502 23888 16458
rect 24228 16250 24256 17478
rect 24768 17060 24820 17066
rect 24768 17002 24820 17008
rect 24780 16454 24808 17002
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 23952 15706 23980 15982
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 24596 15570 24624 15982
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23860 14482 23888 15438
rect 24780 15094 24808 16050
rect 24400 15088 24452 15094
rect 24400 15030 24452 15036
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23400 13394 23428 13806
rect 23492 13530 23520 13942
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 23860 12714 23888 13738
rect 24412 12850 24440 15030
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 24584 14884 24636 14890
rect 24584 14826 24636 14832
rect 24596 14414 24624 14826
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24688 13938 24716 14894
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24872 12918 24900 17870
rect 25056 17678 25084 18022
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 25240 15706 25268 23598
rect 25424 22574 25452 24142
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 25872 19848 25924 19854
rect 25872 19790 25924 19796
rect 25332 19514 25360 19790
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25320 19508 25372 19514
rect 25320 19450 25372 19456
rect 25424 18222 25452 19654
rect 25884 19378 25912 19790
rect 25872 19372 25924 19378
rect 25872 19314 25924 19320
rect 25504 18352 25556 18358
rect 25504 18294 25556 18300
rect 25412 18216 25464 18222
rect 25412 18158 25464 18164
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 25240 15162 25268 15642
rect 25424 15638 25452 18158
rect 25516 17882 25544 18294
rect 25504 17876 25556 17882
rect 25504 17818 25556 17824
rect 25884 16590 25912 19314
rect 25976 17270 26004 26726
rect 26252 25362 26280 27338
rect 27172 25906 27200 27882
rect 27448 27470 27476 37130
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 32404 37120 32456 37126
rect 32404 37062 32456 37068
rect 34612 37120 34664 37126
rect 34612 37062 34664 37068
rect 29460 33312 29512 33318
rect 29460 33254 29512 33260
rect 27896 30592 27948 30598
rect 27896 30534 27948 30540
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 27068 25900 27120 25906
rect 27068 25842 27120 25848
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 27080 25498 27108 25842
rect 27068 25492 27120 25498
rect 27068 25434 27120 25440
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 26056 22636 26108 22642
rect 26056 22578 26108 22584
rect 26068 22234 26096 22578
rect 26056 22228 26108 22234
rect 26056 22170 26108 22176
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25872 16584 25924 16590
rect 25872 16526 25924 16532
rect 25516 16250 25544 16526
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25412 15632 25464 15638
rect 25412 15574 25464 15580
rect 25872 15496 25924 15502
rect 25872 15438 25924 15444
rect 25884 15162 25912 15438
rect 25228 15156 25280 15162
rect 25228 15098 25280 15104
rect 25872 15156 25924 15162
rect 25872 15098 25924 15104
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25608 14550 25636 14962
rect 25596 14544 25648 14550
rect 25596 14486 25648 14492
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 24964 13326 24992 14010
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24400 12844 24452 12850
rect 25780 12844 25832 12850
rect 24400 12786 24452 12792
rect 25700 12804 25780 12832
rect 23848 12708 23900 12714
rect 23848 12650 23900 12656
rect 24412 12238 24440 12786
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23216 11762 23244 12038
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23388 11688 23440 11694
rect 23388 11630 23440 11636
rect 23400 11354 23428 11630
rect 23388 11348 23440 11354
rect 23388 11290 23440 11296
rect 23584 11150 23612 12038
rect 24964 11218 24992 12582
rect 25228 11620 25280 11626
rect 25228 11562 25280 11568
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 24768 11076 24820 11082
rect 24768 11018 24820 11024
rect 24780 10674 24808 11018
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22388 8566 22416 9862
rect 23584 9722 23612 10406
rect 24044 10062 24072 10406
rect 24872 10130 24900 10406
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 23572 9716 23624 9722
rect 23572 9658 23624 9664
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22848 8566 22876 8774
rect 22376 8560 22428 8566
rect 22376 8502 22428 8508
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22848 7410 22876 8502
rect 23032 8498 23060 9522
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 23216 9042 23244 9454
rect 23204 9036 23256 9042
rect 23204 8978 23256 8984
rect 23572 8900 23624 8906
rect 23572 8842 23624 8848
rect 23584 8634 23612 8842
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 24688 8090 24716 9998
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 24780 9042 24808 9658
rect 24964 9178 24992 10542
rect 25056 9178 25084 11494
rect 25240 11354 25268 11562
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25700 10606 25728 12804
rect 25780 12786 25832 12792
rect 26068 12238 26096 18566
rect 26252 18426 26280 25298
rect 27160 25288 27212 25294
rect 27160 25230 27212 25236
rect 27172 24206 27200 25230
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 26332 24132 26384 24138
rect 26332 24074 26384 24080
rect 26344 23730 26372 24074
rect 26608 23792 26660 23798
rect 26608 23734 26660 23740
rect 26332 23724 26384 23730
rect 26332 23666 26384 23672
rect 26620 23322 26648 23734
rect 26608 23316 26660 23322
rect 26608 23258 26660 23264
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26344 17814 26372 19654
rect 27264 19310 27292 27270
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 27344 26376 27396 26382
rect 27344 26318 27396 26324
rect 27356 25294 27384 26318
rect 27620 26240 27672 26246
rect 27620 26182 27672 26188
rect 27632 25702 27660 26182
rect 27620 25696 27672 25702
rect 27620 25638 27672 25644
rect 27344 25288 27396 25294
rect 27344 25230 27396 25236
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 27540 23866 27568 24142
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27356 22234 27384 22646
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27540 21554 27568 23802
rect 27632 22574 27660 25638
rect 27816 25294 27844 26522
rect 27908 26450 27936 30534
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 27896 26444 27948 26450
rect 27896 26386 27948 26392
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27712 25152 27764 25158
rect 27712 25094 27764 25100
rect 27724 23798 27752 25094
rect 28000 24818 28028 29106
rect 28540 25968 28592 25974
rect 28540 25910 28592 25916
rect 28172 25696 28224 25702
rect 28172 25638 28224 25644
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 28000 23798 28028 24754
rect 27712 23792 27764 23798
rect 27712 23734 27764 23740
rect 27988 23792 28040 23798
rect 27988 23734 28040 23740
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27540 20942 27568 21490
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 27724 20482 27752 22510
rect 27988 21004 28040 21010
rect 27988 20946 28040 20952
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27632 20454 27752 20482
rect 27908 20466 27936 20742
rect 27896 20460 27948 20466
rect 27344 19440 27396 19446
rect 27344 19382 27396 19388
rect 27252 19304 27304 19310
rect 27252 19246 27304 19252
rect 27356 18970 27384 19382
rect 27344 18964 27396 18970
rect 27344 18906 27396 18912
rect 26608 18420 26660 18426
rect 26608 18362 26660 18368
rect 26332 17808 26384 17814
rect 26332 17750 26384 17756
rect 26424 17808 26476 17814
rect 26424 17750 26476 17756
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26252 17134 26280 17546
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26252 13326 26280 17070
rect 26344 16454 26372 17614
rect 26332 16448 26384 16454
rect 26332 16390 26384 16396
rect 26436 15570 26464 17750
rect 26620 17746 26648 18362
rect 26792 18284 26844 18290
rect 26792 18226 26844 18232
rect 26608 17740 26660 17746
rect 26608 17682 26660 17688
rect 26608 17264 26660 17270
rect 26608 17206 26660 17212
rect 26516 17060 26568 17066
rect 26516 17002 26568 17008
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26344 14618 26372 14894
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 26344 13938 26372 14282
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26056 12232 26108 12238
rect 26056 12174 26108 12180
rect 25964 11824 26016 11830
rect 25964 11766 26016 11772
rect 25780 11688 25832 11694
rect 25780 11630 25832 11636
rect 25792 11286 25820 11630
rect 25872 11620 25924 11626
rect 25872 11562 25924 11568
rect 25780 11280 25832 11286
rect 25780 11222 25832 11228
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 25884 10538 25912 11562
rect 25976 11354 26004 11766
rect 25964 11348 26016 11354
rect 25964 11290 26016 11296
rect 26068 10742 26096 12174
rect 26148 12096 26200 12102
rect 26148 12038 26200 12044
rect 26160 11150 26188 12038
rect 26148 11144 26200 11150
rect 26148 11086 26200 11092
rect 26056 10736 26108 10742
rect 26056 10678 26108 10684
rect 25872 10532 25924 10538
rect 25872 10474 25924 10480
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 25332 9586 25360 10406
rect 25884 9994 25912 10474
rect 25872 9988 25924 9994
rect 25872 9930 25924 9936
rect 26240 9988 26292 9994
rect 26240 9930 26292 9936
rect 25504 9920 25556 9926
rect 25504 9862 25556 9868
rect 25516 9654 25544 9862
rect 26252 9722 26280 9930
rect 26240 9716 26292 9722
rect 26240 9658 26292 9664
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 24964 8974 24992 9114
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25240 8498 25268 8774
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 24676 8084 24728 8090
rect 24676 8026 24728 8032
rect 25148 7954 25176 8366
rect 25516 8362 25544 9590
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 25504 8356 25556 8362
rect 25504 8298 25556 8304
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23480 7812 23532 7818
rect 23480 7754 23532 7760
rect 23492 7426 23520 7754
rect 23400 7410 23520 7426
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 23388 7404 23520 7410
rect 23440 7398 23520 7404
rect 23388 7346 23440 7352
rect 23492 6798 23520 7398
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 21284 2650 21312 5646
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 22296 2446 22324 6598
rect 23400 6458 23428 6734
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23388 6452 23440 6458
rect 23388 6394 23440 6400
rect 23492 6390 23520 6598
rect 23480 6384 23532 6390
rect 23480 6326 23532 6332
rect 23492 5846 23520 6326
rect 23768 6322 23796 6598
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23480 5840 23532 5846
rect 23480 5782 23532 5788
rect 23860 2650 23888 7822
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 24044 6458 24072 7278
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24412 6390 24440 7142
rect 24400 6384 24452 6390
rect 24400 6326 24452 6332
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 4540 800 4568 2246
rect 5828 800 5856 2246
rect 7760 800 7788 2246
rect 9048 800 9076 2246
rect 10336 800 10364 2382
rect 12268 800 12296 2382
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 800 13584 2246
rect 15488 800 15516 2382
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 16776 800 16804 2246
rect 18708 800 18736 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2246
rect 21284 800 21312 2382
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 23216 800 23244 2246
rect 24504 800 24532 2382
rect 26160 2378 26188 8910
rect 26344 5778 26372 12786
rect 26528 10130 26556 17002
rect 26620 16454 26648 17206
rect 26608 16448 26660 16454
rect 26608 16390 26660 16396
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26620 15162 26648 15438
rect 26608 15156 26660 15162
rect 26608 15098 26660 15104
rect 26804 14346 26832 18226
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27356 17202 27384 17546
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27356 16590 27384 17138
rect 27344 16584 27396 16590
rect 27344 16526 27396 16532
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 26792 14340 26844 14346
rect 26792 14282 26844 14288
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26528 6186 26556 10066
rect 26516 6180 26568 6186
rect 26516 6122 26568 6128
rect 26620 5914 26648 13262
rect 26804 12850 26832 14282
rect 26976 13864 27028 13870
rect 26976 13806 27028 13812
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 26988 11218 27016 13806
rect 27080 11898 27108 14962
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27172 13394 27200 13670
rect 27160 13388 27212 13394
rect 27160 13330 27212 13336
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 27068 11892 27120 11898
rect 27068 11834 27120 11840
rect 27264 11762 27292 12582
rect 27356 12374 27384 16526
rect 27528 14884 27580 14890
rect 27528 14826 27580 14832
rect 27344 12368 27396 12374
rect 27344 12310 27396 12316
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27160 11688 27212 11694
rect 27160 11630 27212 11636
rect 26976 11212 27028 11218
rect 26976 11154 27028 11160
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26712 8090 26740 11018
rect 27172 9625 27200 11630
rect 27540 11354 27568 14826
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27632 10674 27660 20454
rect 27896 20402 27948 20408
rect 27804 19236 27856 19242
rect 27804 19178 27856 19184
rect 27896 19236 27948 19242
rect 27896 19178 27948 19184
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27724 14414 27752 18702
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27816 13546 27844 19178
rect 27908 18970 27936 19178
rect 27896 18964 27948 18970
rect 27896 18906 27948 18912
rect 27896 17672 27948 17678
rect 27896 17614 27948 17620
rect 27908 17338 27936 17614
rect 27896 17332 27948 17338
rect 27896 17274 27948 17280
rect 27896 16652 27948 16658
rect 27896 16594 27948 16600
rect 27724 13518 27844 13546
rect 27724 11830 27752 13518
rect 27804 13456 27856 13462
rect 27804 13398 27856 13404
rect 27816 12850 27844 13398
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27712 11824 27764 11830
rect 27712 11766 27764 11772
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27158 9616 27214 9625
rect 27908 9586 27936 16594
rect 28000 16574 28028 20946
rect 28080 20936 28132 20942
rect 28080 20878 28132 20884
rect 28092 20602 28120 20878
rect 28080 20596 28132 20602
rect 28080 20538 28132 20544
rect 28184 20058 28212 25638
rect 28552 25362 28580 25910
rect 29472 25906 29500 33254
rect 29748 28150 29776 37062
rect 29828 36168 29880 36174
rect 29828 36110 29880 36116
rect 29840 31890 29868 36110
rect 29828 31884 29880 31890
rect 29828 31826 29880 31832
rect 29736 28144 29788 28150
rect 29736 28086 29788 28092
rect 30392 27606 30420 37062
rect 32416 30734 32444 37062
rect 34336 36780 34388 36786
rect 34336 36722 34388 36728
rect 34348 35834 34376 36722
rect 34336 35828 34388 35834
rect 34336 35770 34388 35776
rect 33324 35692 33376 35698
rect 33324 35634 33376 35640
rect 32404 30728 32456 30734
rect 32404 30670 32456 30676
rect 30472 30252 30524 30258
rect 30472 30194 30524 30200
rect 31760 30252 31812 30258
rect 31760 30194 31812 30200
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 29460 25900 29512 25906
rect 29460 25842 29512 25848
rect 28540 25356 28592 25362
rect 28540 25298 28592 25304
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 28908 25220 28960 25226
rect 28908 25162 28960 25168
rect 28356 24812 28408 24818
rect 28356 24754 28408 24760
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28264 24064 28316 24070
rect 28264 24006 28316 24012
rect 28276 23118 28304 24006
rect 28368 23866 28396 24754
rect 28644 24698 28672 24754
rect 28552 24670 28672 24698
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28552 23730 28580 24670
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28356 22568 28408 22574
rect 28356 22510 28408 22516
rect 28368 22098 28396 22510
rect 28552 22438 28580 23666
rect 28540 22432 28592 22438
rect 28540 22374 28592 22380
rect 28920 22166 28948 25162
rect 29012 24410 29040 25230
rect 29828 25152 29880 25158
rect 29828 25094 29880 25100
rect 29552 24744 29604 24750
rect 29552 24686 29604 24692
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 28908 22160 28960 22166
rect 28908 22102 28960 22108
rect 28356 22092 28408 22098
rect 28356 22034 28408 22040
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28460 21146 28488 21898
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 28920 19922 28948 22102
rect 29564 21690 29592 24686
rect 29840 23662 29868 25094
rect 30484 24750 30512 30194
rect 31772 26858 31800 30194
rect 31760 26852 31812 26858
rect 31760 26794 31812 26800
rect 30472 24744 30524 24750
rect 30472 24686 30524 24692
rect 29920 24608 29972 24614
rect 29920 24550 29972 24556
rect 29932 23798 29960 24550
rect 30484 23798 30512 24686
rect 33336 24342 33364 35634
rect 34520 33992 34572 33998
rect 34520 33934 34572 33940
rect 34532 30326 34560 33934
rect 34624 32434 34652 37062
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35452 34202 35480 37198
rect 36648 36378 36676 37198
rect 36740 37126 36768 39200
rect 37462 38176 37518 38185
rect 37462 38111 37518 38120
rect 37476 37330 37504 38111
rect 37464 37324 37516 37330
rect 37464 37266 37516 37272
rect 37740 37256 37792 37262
rect 37740 37198 37792 37204
rect 36728 37120 36780 37126
rect 36728 37062 36780 37068
rect 36636 36372 36688 36378
rect 36636 36314 36688 36320
rect 37280 34944 37332 34950
rect 37280 34886 37332 34892
rect 36452 34604 36504 34610
rect 36452 34546 36504 34552
rect 35440 34196 35492 34202
rect 35440 34138 35492 34144
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34612 32428 34664 32434
rect 34612 32370 34664 32376
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34520 30320 34572 30326
rect 34520 30262 34572 30268
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 36464 29306 36492 34546
rect 36452 29300 36504 29306
rect 36452 29242 36504 29248
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36648 25498 36676 29106
rect 37292 26994 37320 34886
rect 37372 31884 37424 31890
rect 37372 31826 37424 31832
rect 37280 26988 37332 26994
rect 37280 26930 37332 26936
rect 37280 26784 37332 26790
rect 37280 26726 37332 26732
rect 36636 25492 36688 25498
rect 36636 25434 36688 25440
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33324 24336 33376 24342
rect 33324 24278 33376 24284
rect 29920 23792 29972 23798
rect 29920 23734 29972 23740
rect 30472 23792 30524 23798
rect 30472 23734 30524 23740
rect 29828 23656 29880 23662
rect 29828 23598 29880 23604
rect 29840 23322 29868 23598
rect 30104 23588 30156 23594
rect 30104 23530 30156 23536
rect 29828 23316 29880 23322
rect 29828 23258 29880 23264
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29564 21078 29592 21626
rect 29552 21072 29604 21078
rect 29552 21014 29604 21020
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29932 20602 29960 20878
rect 29920 20596 29972 20602
rect 29920 20538 29972 20544
rect 29460 20460 29512 20466
rect 29460 20402 29512 20408
rect 28632 19916 28684 19922
rect 28632 19858 28684 19864
rect 28908 19916 28960 19922
rect 28908 19858 28960 19864
rect 28356 19780 28408 19786
rect 28356 19722 28408 19728
rect 28368 18970 28396 19722
rect 28644 19378 28672 19858
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28632 19372 28684 19378
rect 28632 19314 28684 19320
rect 28356 18964 28408 18970
rect 28356 18906 28408 18912
rect 28460 18834 28488 19314
rect 28448 18828 28500 18834
rect 28448 18770 28500 18776
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 28000 16546 28120 16574
rect 27988 15496 28040 15502
rect 27988 15438 28040 15444
rect 28000 15162 28028 15438
rect 28092 15366 28120 16546
rect 28368 15910 28396 18702
rect 28448 16040 28500 16046
rect 28448 15982 28500 15988
rect 28540 16040 28592 16046
rect 28540 15982 28592 15988
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28460 15570 28488 15982
rect 28552 15706 28580 15982
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 28448 15564 28500 15570
rect 28448 15506 28500 15512
rect 28540 15428 28592 15434
rect 28540 15370 28592 15376
rect 28080 15360 28132 15366
rect 28080 15302 28132 15308
rect 27988 15156 28040 15162
rect 27988 15098 28040 15104
rect 28552 15026 28580 15370
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28644 14618 28672 19314
rect 29472 18766 29500 20402
rect 29460 18760 29512 18766
rect 29460 18702 29512 18708
rect 29644 18760 29696 18766
rect 29644 18702 29696 18708
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29656 18426 29684 18702
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29840 17882 29868 18702
rect 29920 18080 29972 18086
rect 29920 18022 29972 18028
rect 29828 17876 29880 17882
rect 29828 17818 29880 17824
rect 29932 17678 29960 18022
rect 29920 17672 29972 17678
rect 29920 17614 29972 17620
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29012 17202 29040 17478
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 29828 16040 29880 16046
rect 29828 15982 29880 15988
rect 28632 14612 28684 14618
rect 28632 14554 28684 14560
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 28276 14074 28304 14350
rect 28448 14272 28500 14278
rect 28448 14214 28500 14220
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28460 13938 28488 14214
rect 28448 13932 28500 13938
rect 28448 13874 28500 13880
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 28092 12782 28120 13126
rect 28080 12776 28132 12782
rect 28080 12718 28132 12724
rect 28092 11898 28120 12718
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 29564 9654 29592 15982
rect 29840 15706 29868 15982
rect 30116 15978 30144 23530
rect 36452 23520 36504 23526
rect 36452 23462 36504 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30196 21888 30248 21894
rect 30196 21830 30248 21836
rect 30208 20466 30236 21830
rect 30944 21146 30972 21966
rect 33048 21548 33100 21554
rect 33048 21490 33100 21496
rect 30932 21140 30984 21146
rect 30932 21082 30984 21088
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 31128 20602 31156 20878
rect 31116 20596 31168 20602
rect 31116 20538 31168 20544
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 31024 20460 31076 20466
rect 31024 20402 31076 20408
rect 30380 20392 30432 20398
rect 30380 20334 30432 20340
rect 30392 20058 30420 20334
rect 30472 20256 30524 20262
rect 30472 20198 30524 20204
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 30300 18290 30328 19790
rect 30484 18970 30512 20198
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30288 18284 30340 18290
rect 30288 18226 30340 18232
rect 30380 17604 30432 17610
rect 30380 17546 30432 17552
rect 30392 17202 30420 17546
rect 30380 17196 30432 17202
rect 30380 17138 30432 17144
rect 30104 15972 30156 15978
rect 30104 15914 30156 15920
rect 29828 15700 29880 15706
rect 29828 15642 29880 15648
rect 29920 14476 29972 14482
rect 29920 14418 29972 14424
rect 29932 13530 29960 14418
rect 29920 13524 29972 13530
rect 29920 13466 29972 13472
rect 30484 13394 30512 18906
rect 30932 18216 30984 18222
rect 30932 18158 30984 18164
rect 30944 17746 30972 18158
rect 31036 18154 31064 20402
rect 31760 20256 31812 20262
rect 31760 20198 31812 20204
rect 31024 18148 31076 18154
rect 31024 18090 31076 18096
rect 30932 17740 30984 17746
rect 30932 17682 30984 17688
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30576 17338 30604 17614
rect 31024 17536 31076 17542
rect 31024 17478 31076 17484
rect 31036 17338 31064 17478
rect 30564 17332 30616 17338
rect 30564 17274 30616 17280
rect 31024 17332 31076 17338
rect 31024 17274 31076 17280
rect 31036 16658 31064 17274
rect 31772 17270 31800 20198
rect 33060 20058 33088 21490
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 36464 20466 36492 23462
rect 37292 22098 37320 26726
rect 37384 26450 37412 31826
rect 37752 27470 37780 37198
rect 38028 36922 38056 39200
rect 39316 37466 39344 39200
rect 39304 37460 39356 37466
rect 39304 37402 39356 37408
rect 38016 36916 38068 36922
rect 38016 36858 38068 36864
rect 38198 36816 38254 36825
rect 38198 36751 38254 36760
rect 38212 36378 38240 36751
rect 38200 36372 38252 36378
rect 38200 36314 38252 36320
rect 38016 36168 38068 36174
rect 38016 36110 38068 36116
rect 38028 34746 38056 36110
rect 38292 35080 38344 35086
rect 38292 35022 38344 35028
rect 38304 34785 38332 35022
rect 38290 34776 38346 34785
rect 38016 34740 38068 34746
rect 38290 34711 38346 34720
rect 38016 34682 38068 34688
rect 38292 33516 38344 33522
rect 38292 33458 38344 33464
rect 38304 33425 38332 33458
rect 38290 33416 38346 33425
rect 38290 33351 38346 33360
rect 38108 31816 38160 31822
rect 38108 31758 38160 31764
rect 38120 31385 38148 31758
rect 38106 31376 38162 31385
rect 38106 31311 38162 31320
rect 38200 30048 38252 30054
rect 38198 30016 38200 30025
rect 38252 30016 38254 30025
rect 38198 29951 38254 29960
rect 38200 29028 38252 29034
rect 38200 28970 38252 28976
rect 38212 28665 38240 28970
rect 38198 28656 38254 28665
rect 38198 28591 38254 28600
rect 37740 27464 37792 27470
rect 37740 27406 37792 27412
rect 38292 26988 38344 26994
rect 38292 26930 38344 26936
rect 38304 26625 38332 26930
rect 38290 26616 38346 26625
rect 38290 26551 38346 26560
rect 37372 26444 37424 26450
rect 37372 26386 37424 26392
rect 38108 25832 38160 25838
rect 38108 25774 38160 25780
rect 38120 25498 38148 25774
rect 38108 25492 38160 25498
rect 38108 25434 38160 25440
rect 38292 25288 38344 25294
rect 38290 25256 38292 25265
rect 38344 25256 38346 25265
rect 38290 25191 38346 25200
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 38304 23225 38332 23666
rect 38290 23216 38346 23225
rect 38290 23151 38346 23160
rect 37280 22092 37332 22098
rect 37280 22034 37332 22040
rect 38200 21888 38252 21894
rect 38198 21856 38200 21865
rect 38252 21856 38254 21865
rect 38198 21791 38254 21800
rect 36452 20460 36504 20466
rect 36452 20402 36504 20408
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 33048 20052 33100 20058
rect 33048 19994 33100 20000
rect 38292 19848 38344 19854
rect 38290 19816 38292 19825
rect 38344 19816 38346 19825
rect 38290 19751 38346 19760
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 38292 18760 38344 18766
rect 38292 18702 38344 18708
rect 38304 18465 38332 18702
rect 38290 18456 38346 18465
rect 38290 18391 38346 18400
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 31760 17264 31812 17270
rect 31760 17206 31812 17212
rect 31024 16652 31076 16658
rect 31024 16594 31076 16600
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 30668 15706 30696 16526
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 30656 15700 30708 15706
rect 30656 15642 30708 15648
rect 31128 15638 31156 16390
rect 31116 15632 31168 15638
rect 31116 15574 31168 15580
rect 30564 15496 30616 15502
rect 30564 15438 30616 15444
rect 30576 15162 30604 15438
rect 30564 15156 30616 15162
rect 30564 15098 30616 15104
rect 30840 13456 30892 13462
rect 30840 13398 30892 13404
rect 30472 13388 30524 13394
rect 30472 13330 30524 13336
rect 30852 12986 30880 13398
rect 30840 12980 30892 12986
rect 30840 12922 30892 12928
rect 30852 12238 30880 12922
rect 30840 12232 30892 12238
rect 30840 12174 30892 12180
rect 31772 11694 31800 17206
rect 38292 17196 38344 17202
rect 38292 17138 38344 17144
rect 32404 17128 32456 17134
rect 38304 17105 38332 17138
rect 32404 17070 32456 17076
rect 38290 17096 38346 17105
rect 32416 16794 32444 17070
rect 38290 17031 38346 17040
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 32404 16788 32456 16794
rect 32404 16730 32456 16736
rect 33598 16552 33654 16561
rect 33598 16487 33654 16496
rect 33612 16454 33640 16487
rect 35912 16454 35940 16934
rect 37096 16652 37148 16658
rect 37096 16594 37148 16600
rect 33600 16448 33652 16454
rect 33600 16390 33652 16396
rect 35900 16448 35952 16454
rect 35900 16390 35952 16396
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 32404 15496 32456 15502
rect 32404 15438 32456 15444
rect 32416 11898 32444 15438
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 37108 14074 37136 16594
rect 38200 15360 38252 15366
rect 38200 15302 38252 15308
rect 38212 15065 38240 15302
rect 38198 15056 38254 15065
rect 38198 14991 38254 15000
rect 37096 14068 37148 14074
rect 37096 14010 37148 14016
rect 38292 13932 38344 13938
rect 38292 13874 38344 13880
rect 38304 13705 38332 13874
rect 38290 13696 38346 13705
rect 34934 13628 35242 13637
rect 38290 13631 38346 13640
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 36912 13388 36964 13394
rect 36912 13330 36964 13336
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 32496 12096 32548 12102
rect 32496 12038 32548 12044
rect 32404 11892 32456 11898
rect 32404 11834 32456 11840
rect 32508 11762 32536 12038
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 31760 11688 31812 11694
rect 31760 11630 31812 11636
rect 34060 11552 34112 11558
rect 34060 11494 34112 11500
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29552 9648 29604 9654
rect 29552 9590 29604 9596
rect 27158 9551 27214 9560
rect 27896 9580 27948 9586
rect 27896 9522 27948 9528
rect 27908 8566 27936 9522
rect 28724 8900 28776 8906
rect 28724 8842 28776 8848
rect 27896 8560 27948 8566
rect 27896 8502 27948 8508
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 28736 7886 28764 8842
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 26608 5908 26660 5914
rect 26608 5850 26660 5856
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 27172 2650 27200 6258
rect 27540 2650 27568 6734
rect 27804 4480 27856 4486
rect 27804 4422 27856 4428
rect 27816 2990 27844 4422
rect 27804 2984 27856 2990
rect 27804 2926 27856 2932
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 27908 2582 27936 7822
rect 29748 2650 29776 11086
rect 31392 11008 31444 11014
rect 31392 10950 31444 10956
rect 31404 10062 31432 10950
rect 32312 10600 32364 10606
rect 32312 10542 32364 10548
rect 31392 10056 31444 10062
rect 31392 9998 31444 10004
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 29828 6724 29880 6730
rect 29828 6666 29880 6672
rect 29840 5914 29868 6666
rect 29828 5908 29880 5914
rect 29828 5850 29880 5856
rect 30300 5302 30328 8774
rect 31668 7744 31720 7750
rect 31668 7686 31720 7692
rect 30288 5296 30340 5302
rect 30288 5238 30340 5244
rect 31680 5234 31708 7686
rect 31668 5228 31720 5234
rect 31668 5170 31720 5176
rect 32324 2650 32352 10542
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 33152 10062 33180 10406
rect 33140 10056 33192 10062
rect 33140 9998 33192 10004
rect 32864 9920 32916 9926
rect 32864 9862 32916 9868
rect 32876 8974 32904 9862
rect 33048 9580 33100 9586
rect 33048 9522 33100 9528
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 33060 2650 33088 9522
rect 34072 7410 34100 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 36924 10810 36952 13330
rect 38292 11756 38344 11762
rect 38292 11698 38344 11704
rect 38304 11665 38332 11698
rect 38290 11656 38346 11665
rect 38290 11591 38346 11600
rect 36912 10804 36964 10810
rect 36912 10746 36964 10752
rect 38292 10668 38344 10674
rect 38292 10610 38344 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 38304 10305 38332 10610
rect 38290 10296 38346 10305
rect 38290 10231 38346 10240
rect 38016 9920 38068 9926
rect 38016 9862 38068 9868
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34060 7404 34112 7410
rect 34060 7346 34112 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 36728 5704 36780 5710
rect 36728 5646 36780 5652
rect 37188 5704 37240 5710
rect 37188 5646 37240 5652
rect 33692 5092 33744 5098
rect 33692 5034 33744 5040
rect 29736 2644 29788 2650
rect 29736 2586 29788 2592
rect 32312 2644 32364 2650
rect 32312 2586 32364 2592
rect 33048 2644 33100 2650
rect 33048 2586 33100 2592
rect 27896 2576 27948 2582
rect 27896 2518 27948 2524
rect 33704 2514 33732 5034
rect 34060 5024 34112 5030
rect 34060 4966 34112 4972
rect 34072 3126 34100 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35624 4616 35676 4622
rect 35624 4558 35676 4564
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34060 3120 34112 3126
rect 34060 3062 34112 3068
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35636 2650 35664 4558
rect 36740 3194 36768 5646
rect 37200 5545 37228 5646
rect 37186 5536 37242 5545
rect 37186 5471 37242 5480
rect 38028 3534 38056 9862
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38200 7200 38252 7206
rect 38200 7142 38252 7148
rect 38212 6905 38240 7142
rect 38198 6896 38254 6905
rect 38198 6831 38254 6840
rect 38016 3528 38068 3534
rect 38016 3470 38068 3476
rect 38198 3496 38254 3505
rect 38198 3431 38254 3440
rect 38212 3398 38240 3431
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 36728 3188 36780 3194
rect 36728 3130 36780 3136
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 35624 2644 35676 2650
rect 35624 2586 35676 2592
rect 33692 2508 33744 2514
rect 33692 2450 33744 2456
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 26148 2372 26200 2378
rect 26148 2314 26200 2320
rect 26436 800 26464 2382
rect 27724 800 27752 2382
rect 29012 800 29040 2382
rect 30944 800 30972 2382
rect 32232 800 32260 2382
rect 34164 800 34192 2382
rect 35452 800 35480 2382
rect 36924 2145 36952 2994
rect 38200 2848 38252 2854
rect 38200 2790 38252 2796
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 36910 2136 36966 2145
rect 36910 2071 36966 2080
rect 37384 800 37412 2246
rect 18 200 74 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 7746 200 7802 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 12254 200 12310 800
rect 13542 200 13598 800
rect 15474 200 15530 800
rect 16762 200 16818 800
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 26422 200 26478 800
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 37370 200 37426 800
rect 38212 105 38240 2790
rect 38660 2372 38712 2378
rect 38660 2314 38712 2320
rect 38672 800 38700 2314
rect 38658 200 38714 800
rect 38198 96 38254 105
rect 38198 31 38254 40
<< via2 >>
rect 2778 39480 2834 39536
rect 3146 37440 3202 37496
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1766 36116 1768 36136
rect 1768 36116 1820 36136
rect 1820 36116 1822 36136
rect 1766 36080 1822 36116
rect 1766 34040 1822 34096
rect 1766 32680 1822 32736
rect 1766 30640 1822 30696
rect 1950 31728 2006 31784
rect 1766 29280 1822 29336
rect 1766 27920 1822 27976
rect 1582 14320 1638 14376
rect 1766 24520 1822 24576
rect 1766 22480 1822 22536
rect 1766 21120 1822 21176
rect 1950 20460 2006 20496
rect 1950 20440 1952 20460
rect 1952 20440 2004 20460
rect 2004 20440 2006 20460
rect 1766 19796 1768 19816
rect 1768 19796 1820 19816
rect 1820 19796 1822 19816
rect 1766 19760 1822 19796
rect 3146 25880 3202 25936
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 1766 17720 1822 17776
rect 1766 16360 1822 16416
rect 1766 12960 1822 13016
rect 1582 10920 1638 10976
rect 1766 9560 1822 9616
rect 1766 8200 1822 8256
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 6458 19780 6514 19816
rect 6458 19760 6460 19780
rect 6460 19760 6512 19780
rect 6512 19760 6514 19780
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1766 6180 1822 6216
rect 1766 6160 1768 6180
rect 1768 6160 1820 6180
rect 1820 6160 1822 6180
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1766 4800 1822 4856
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1766 2760 1822 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5998 6840 6054 6896
rect 7838 20576 7894 20632
rect 10046 26868 10048 26888
rect 10048 26868 10100 26888
rect 10100 26868 10102 26888
rect 10046 26832 10102 26868
rect 9586 23296 9642 23352
rect 5722 5616 5778 5672
rect 11058 22072 11114 22128
rect 12714 27124 12770 27160
rect 12714 27104 12716 27124
rect 12716 27104 12768 27124
rect 12768 27104 12770 27124
rect 10782 9596 10784 9616
rect 10784 9596 10836 9616
rect 10836 9596 10838 9616
rect 10782 9560 10838 9596
rect 12346 13232 12402 13288
rect 15566 27104 15622 27160
rect 14646 20576 14702 20632
rect 16026 22108 16028 22128
rect 16028 22108 16080 22128
rect 16080 22108 16082 22128
rect 16026 22072 16082 22108
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 17406 26868 17408 26888
rect 17408 26868 17460 26888
rect 17460 26868 17462 26888
rect 17406 26832 17462 26868
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 16302 23296 16358 23352
rect 15658 13268 15660 13288
rect 15660 13268 15712 13288
rect 15712 13268 15714 13288
rect 15658 13232 15714 13268
rect 16118 19760 16174 19816
rect 15842 9324 15844 9344
rect 15844 9324 15896 9344
rect 15896 9324 15898 9344
rect 15842 9288 15898 9324
rect 16026 9152 16082 9208
rect 16762 9324 16764 9344
rect 16764 9324 16816 9344
rect 16816 9324 16818 9344
rect 16762 9288 16818 9324
rect 17406 20440 17462 20496
rect 17406 16496 17462 16552
rect 17222 9560 17278 9616
rect 16578 5636 16634 5672
rect 16578 5616 16580 5636
rect 16580 5616 16632 5636
rect 16632 5616 16634 5636
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19522 25200 19578 25256
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19798 23196 19800 23216
rect 19800 23196 19852 23216
rect 19852 23196 19854 23216
rect 19798 23160 19854 23196
rect 18050 9152 18106 9208
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 20534 20712 20590 20768
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19430 11192 19486 11248
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19522 10648 19578 10704
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 18878 6840 18934 6896
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20626 9560 20682 9616
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 2778 1400 2834 1456
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 27158 9560 27214 9616
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 37462 38120 37518 38176
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 38198 36760 38254 36816
rect 38290 34720 38346 34776
rect 38290 33360 38346 33416
rect 38106 31320 38162 31376
rect 38198 29996 38200 30016
rect 38200 29996 38252 30016
rect 38252 29996 38254 30016
rect 38198 29960 38254 29996
rect 38198 28600 38254 28656
rect 38290 26560 38346 26616
rect 38290 25236 38292 25256
rect 38292 25236 38344 25256
rect 38344 25236 38346 25256
rect 38290 25200 38346 25236
rect 38290 23160 38346 23216
rect 38198 21836 38200 21856
rect 38200 21836 38252 21856
rect 38252 21836 38254 21856
rect 38198 21800 38254 21836
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 38290 19796 38292 19816
rect 38292 19796 38344 19816
rect 38344 19796 38346 19816
rect 38290 19760 38346 19796
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 38290 18400 38346 18456
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 38290 17040 38346 17096
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 33598 16496 33654 16552
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 38198 15000 38254 15056
rect 38290 13640 38346 13696
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 38290 11600 38346 11656
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 38290 10240 38346 10296
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37186 5480 37242 5536
rect 38198 8880 38254 8936
rect 38198 6840 38254 6896
rect 38198 3440 38254 3496
rect 36910 2080 36966 2136
rect 38198 40 38254 96
<< metal3 >>
rect 200 39538 800 39568
rect 2773 39538 2839 39541
rect 200 39536 2839 39538
rect 200 39480 2778 39536
rect 2834 39480 2839 39536
rect 200 39478 2839 39480
rect 200 39448 800 39478
rect 2773 39475 2839 39478
rect 37457 38178 37523 38181
rect 39200 38178 39800 38208
rect 37457 38176 39800 38178
rect 37457 38120 37462 38176
rect 37518 38120 39800 38176
rect 37457 38118 39800 38120
rect 37457 38115 37523 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 3141 37498 3207 37501
rect 200 37496 3207 37498
rect 200 37440 3146 37496
rect 3202 37440 3207 37496
rect 200 37438 3207 37440
rect 200 37408 800 37438
rect 3141 37435 3207 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 38193 36818 38259 36821
rect 39200 36818 39800 36848
rect 38193 36816 39800 36818
rect 38193 36760 38198 36816
rect 38254 36760 39800 36816
rect 38193 36758 39800 36760
rect 38193 36755 38259 36758
rect 39200 36728 39800 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1761 36138 1827 36141
rect 200 36136 1827 36138
rect 200 36080 1766 36136
rect 1822 36080 1827 36136
rect 200 36078 1827 36080
rect 200 36048 800 36078
rect 1761 36075 1827 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 38285 34778 38351 34781
rect 39200 34778 39800 34808
rect 38285 34776 39800 34778
rect 38285 34720 38290 34776
rect 38346 34720 39800 34776
rect 38285 34718 39800 34720
rect 38285 34715 38351 34718
rect 39200 34688 39800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1761 34098 1827 34101
rect 200 34096 1827 34098
rect 200 34040 1766 34096
rect 1822 34040 1827 34096
rect 200 34038 1827 34040
rect 200 34008 800 34038
rect 1761 34035 1827 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 38285 33418 38351 33421
rect 39200 33418 39800 33448
rect 38285 33416 39800 33418
rect 38285 33360 38290 33416
rect 38346 33360 39800 33416
rect 38285 33358 39800 33360
rect 38285 33355 38351 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32768
rect 1761 32738 1827 32741
rect 200 32736 1827 32738
rect 200 32680 1766 32736
rect 1822 32680 1827 32736
rect 200 32678 1827 32680
rect 200 32648 800 32678
rect 1761 32675 1827 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1945 31786 2011 31789
rect 2078 31786 2084 31788
rect 1945 31784 2084 31786
rect 1945 31728 1950 31784
rect 2006 31728 2084 31784
rect 1945 31726 2084 31728
rect 1945 31723 2011 31726
rect 2078 31724 2084 31726
rect 2148 31724 2154 31788
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 38101 31378 38167 31381
rect 39200 31378 39800 31408
rect 38101 31376 39800 31378
rect 38101 31320 38106 31376
rect 38162 31320 39800 31376
rect 38101 31318 39800 31320
rect 38101 31315 38167 31318
rect 39200 31288 39800 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38193 30018 38259 30021
rect 39200 30018 39800 30048
rect 38193 30016 39800 30018
rect 38193 29960 38198 30016
rect 38254 29960 39800 30016
rect 38193 29958 39800 29960
rect 38193 29955 38259 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1761 29338 1827 29341
rect 200 29336 1827 29338
rect 200 29280 1766 29336
rect 1822 29280 1827 29336
rect 200 29278 1827 29280
rect 200 29248 800 29278
rect 1761 29275 1827 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 38193 28658 38259 28661
rect 39200 28658 39800 28688
rect 38193 28656 39800 28658
rect 38193 28600 38198 28656
rect 38254 28600 39800 28656
rect 38193 28598 39800 28600
rect 38193 28595 38259 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 200 27978 800 28008
rect 1761 27978 1827 27981
rect 200 27976 1827 27978
rect 200 27920 1766 27976
rect 1822 27920 1827 27976
rect 200 27918 1827 27920
rect 200 27888 800 27918
rect 1761 27915 1827 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 12709 27162 12775 27165
rect 15561 27162 15627 27165
rect 12709 27160 15627 27162
rect 12709 27104 12714 27160
rect 12770 27104 15566 27160
rect 15622 27104 15627 27160
rect 12709 27102 15627 27104
rect 12709 27099 12775 27102
rect 15561 27099 15627 27102
rect 10041 26890 10107 26893
rect 17401 26890 17467 26893
rect 10041 26888 17467 26890
rect 10041 26832 10046 26888
rect 10102 26832 17406 26888
rect 17462 26832 17467 26888
rect 10041 26830 17467 26832
rect 10041 26827 10107 26830
rect 17401 26827 17467 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 38285 26618 38351 26621
rect 39200 26618 39800 26648
rect 38285 26616 39800 26618
rect 38285 26560 38290 26616
rect 38346 26560 39800 26616
rect 38285 26558 39800 26560
rect 38285 26555 38351 26558
rect 39200 26528 39800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25938 800 25968
rect 3141 25938 3207 25941
rect 200 25936 3207 25938
rect 200 25880 3146 25936
rect 3202 25880 3207 25936
rect 200 25878 3207 25880
rect 200 25848 800 25878
rect 3141 25875 3207 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19517 25258 19583 25261
rect 20110 25258 20116 25260
rect 19517 25256 20116 25258
rect 19517 25200 19522 25256
rect 19578 25200 20116 25256
rect 19517 25198 20116 25200
rect 19517 25195 19583 25198
rect 20110 25196 20116 25198
rect 20180 25196 20186 25260
rect 38285 25258 38351 25261
rect 39200 25258 39800 25288
rect 38285 25256 39800 25258
rect 38285 25200 38290 25256
rect 38346 25200 39800 25256
rect 38285 25198 39800 25200
rect 38285 25195 38351 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 200 24578 800 24608
rect 1761 24578 1827 24581
rect 200 24576 1827 24578
rect 200 24520 1766 24576
rect 1822 24520 1827 24576
rect 200 24518 1827 24520
rect 200 24488 800 24518
rect 1761 24515 1827 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 9581 23354 9647 23357
rect 16297 23354 16363 23357
rect 9581 23352 16363 23354
rect 9581 23296 9586 23352
rect 9642 23296 16302 23352
rect 16358 23296 16363 23352
rect 9581 23294 16363 23296
rect 9581 23291 9647 23294
rect 16297 23291 16363 23294
rect 2078 23156 2084 23220
rect 2148 23218 2154 23220
rect 19793 23218 19859 23221
rect 2148 23216 19859 23218
rect 2148 23160 19798 23216
rect 19854 23160 19859 23216
rect 2148 23158 19859 23160
rect 2148 23156 2154 23158
rect 19793 23155 19859 23158
rect 38285 23218 38351 23221
rect 39200 23218 39800 23248
rect 38285 23216 39800 23218
rect 38285 23160 38290 23216
rect 38346 23160 39800 23216
rect 38285 23158 39800 23160
rect 38285 23155 38351 23158
rect 39200 23128 39800 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 11053 22130 11119 22133
rect 16021 22130 16087 22133
rect 11053 22128 16087 22130
rect 11053 22072 11058 22128
rect 11114 22072 16026 22128
rect 16082 22072 16087 22128
rect 11053 22070 16087 22072
rect 11053 22067 11119 22070
rect 16021 22067 16087 22070
rect 38193 21858 38259 21861
rect 39200 21858 39800 21888
rect 38193 21856 39800 21858
rect 38193 21800 38198 21856
rect 38254 21800 39800 21856
rect 38193 21798 39800 21800
rect 38193 21795 38259 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1761 21178 1827 21181
rect 200 21176 1827 21178
rect 200 21120 1766 21176
rect 1822 21120 1827 21176
rect 200 21118 1827 21120
rect 200 21088 800 21118
rect 1761 21115 1827 21118
rect 20529 20770 20595 20773
rect 20662 20770 20668 20772
rect 20529 20768 20668 20770
rect 20529 20712 20534 20768
rect 20590 20712 20668 20768
rect 20529 20710 20668 20712
rect 20529 20707 20595 20710
rect 20662 20708 20668 20710
rect 20732 20708 20738 20772
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 7833 20634 7899 20637
rect 14641 20634 14707 20637
rect 7833 20632 14707 20634
rect 7833 20576 7838 20632
rect 7894 20576 14646 20632
rect 14702 20576 14707 20632
rect 7833 20574 14707 20576
rect 7833 20571 7899 20574
rect 14641 20571 14707 20574
rect 1945 20498 2011 20501
rect 17401 20498 17467 20501
rect 1945 20496 17467 20498
rect 1945 20440 1950 20496
rect 2006 20440 17406 20496
rect 17462 20440 17467 20496
rect 1945 20438 17467 20440
rect 1945 20435 2011 20438
rect 17401 20435 17467 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 200 19818 800 19848
rect 1761 19818 1827 19821
rect 200 19816 1827 19818
rect 200 19760 1766 19816
rect 1822 19760 1827 19816
rect 200 19758 1827 19760
rect 200 19728 800 19758
rect 1761 19755 1827 19758
rect 6453 19818 6519 19821
rect 16113 19818 16179 19821
rect 6453 19816 16179 19818
rect 6453 19760 6458 19816
rect 6514 19760 16118 19816
rect 16174 19760 16179 19816
rect 6453 19758 16179 19760
rect 6453 19755 6519 19758
rect 16113 19755 16179 19758
rect 38285 19818 38351 19821
rect 39200 19818 39800 19848
rect 38285 19816 39800 19818
rect 38285 19760 38290 19816
rect 38346 19760 39800 19816
rect 38285 19758 39800 19760
rect 38285 19755 38351 19758
rect 39200 19728 39800 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 38285 18458 38351 18461
rect 39200 18458 39800 18488
rect 38285 18456 39800 18458
rect 38285 18400 38290 18456
rect 38346 18400 39800 18456
rect 38285 18398 39800 18400
rect 38285 18395 38351 18398
rect 39200 18368 39800 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1761 17778 1827 17781
rect 200 17776 1827 17778
rect 200 17720 1766 17776
rect 1822 17720 1827 17776
rect 200 17718 1827 17720
rect 200 17688 800 17718
rect 1761 17715 1827 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 38285 17098 38351 17101
rect 39200 17098 39800 17128
rect 38285 17096 39800 17098
rect 38285 17040 38290 17096
rect 38346 17040 39800 17096
rect 38285 17038 39800 17040
rect 38285 17035 38351 17038
rect 39200 17008 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 17401 16554 17467 16557
rect 20110 16554 20116 16556
rect 17401 16552 20116 16554
rect 17401 16496 17406 16552
rect 17462 16496 20116 16552
rect 17401 16494 20116 16496
rect 17401 16491 17467 16494
rect 20110 16492 20116 16494
rect 20180 16492 20186 16556
rect 20662 16492 20668 16556
rect 20732 16554 20738 16556
rect 33593 16554 33659 16557
rect 20732 16552 33659 16554
rect 20732 16496 33598 16552
rect 33654 16496 33659 16552
rect 20732 16494 33659 16496
rect 20732 16492 20738 16494
rect 33593 16491 33659 16494
rect 200 16418 800 16448
rect 1761 16418 1827 16421
rect 200 16416 1827 16418
rect 200 16360 1766 16416
rect 1822 16360 1827 16416
rect 200 16358 1827 16360
rect 200 16328 800 16358
rect 1761 16355 1827 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 38193 15058 38259 15061
rect 39200 15058 39800 15088
rect 38193 15056 39800 15058
rect 38193 15000 38198 15056
rect 38254 15000 39800 15056
rect 38193 14998 39800 15000
rect 38193 14995 38259 14998
rect 39200 14968 39800 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14408
rect 1577 14378 1643 14381
rect 200 14376 1643 14378
rect 200 14320 1582 14376
rect 1638 14320 1643 14376
rect 200 14318 1643 14320
rect 200 14288 800 14318
rect 1577 14315 1643 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 38285 13698 38351 13701
rect 39200 13698 39800 13728
rect 38285 13696 39800 13698
rect 38285 13640 38290 13696
rect 38346 13640 39800 13696
rect 38285 13638 39800 13640
rect 38285 13635 38351 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 12341 13290 12407 13293
rect 15653 13290 15719 13293
rect 12341 13288 15719 13290
rect 12341 13232 12346 13288
rect 12402 13232 15658 13288
rect 15714 13232 15719 13288
rect 12341 13230 15719 13232
rect 12341 13227 12407 13230
rect 15653 13227 15719 13230
rect 19570 13088 19886 13089
rect 200 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 1761 13018 1827 13021
rect 200 13016 1827 13018
rect 200 12960 1766 13016
rect 1822 12960 1827 13016
rect 200 12958 1827 12960
rect 200 12928 800 12958
rect 1761 12955 1827 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 38285 11658 38351 11661
rect 39200 11658 39800 11688
rect 38285 11656 39800 11658
rect 38285 11600 38290 11656
rect 38346 11600 39800 11656
rect 38285 11598 39800 11600
rect 38285 11595 38351 11598
rect 39200 11568 39800 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19425 11250 19491 11253
rect 19382 11248 19491 11250
rect 19382 11192 19430 11248
rect 19486 11192 19491 11248
rect 19382 11187 19491 11192
rect 200 10978 800 11008
rect 1577 10978 1643 10981
rect 200 10976 1643 10978
rect 200 10920 1582 10976
rect 1638 10920 1643 10976
rect 200 10918 1643 10920
rect 200 10888 800 10918
rect 1577 10915 1643 10918
rect 19382 10706 19442 11187
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 19517 10706 19583 10709
rect 19382 10704 19583 10706
rect 19382 10648 19522 10704
rect 19578 10648 19583 10704
rect 19382 10646 19583 10648
rect 19517 10643 19583 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 38285 10298 38351 10301
rect 39200 10298 39800 10328
rect 38285 10296 39800 10298
rect 38285 10240 38290 10296
rect 38346 10240 39800 10296
rect 38285 10238 39800 10240
rect 38285 10235 38351 10238
rect 39200 10208 39800 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9648
rect 1761 9618 1827 9621
rect 200 9616 1827 9618
rect 200 9560 1766 9616
rect 1822 9560 1827 9616
rect 200 9558 1827 9560
rect 200 9528 800 9558
rect 1761 9555 1827 9558
rect 10777 9618 10843 9621
rect 17217 9618 17283 9621
rect 10777 9616 17283 9618
rect 10777 9560 10782 9616
rect 10838 9560 17222 9616
rect 17278 9560 17283 9616
rect 10777 9558 17283 9560
rect 10777 9555 10843 9558
rect 17217 9555 17283 9558
rect 20621 9618 20687 9621
rect 27153 9618 27219 9621
rect 20621 9616 27219 9618
rect 20621 9560 20626 9616
rect 20682 9560 27158 9616
rect 27214 9560 27219 9616
rect 20621 9558 27219 9560
rect 20621 9555 20687 9558
rect 27153 9555 27219 9558
rect 15837 9346 15903 9349
rect 16757 9346 16823 9349
rect 15837 9344 16823 9346
rect 15837 9288 15842 9344
rect 15898 9288 16762 9344
rect 16818 9288 16823 9344
rect 15837 9286 16823 9288
rect 15837 9283 15903 9286
rect 16757 9283 16823 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 16021 9210 16087 9213
rect 18045 9210 18111 9213
rect 16021 9208 18111 9210
rect 16021 9152 16026 9208
rect 16082 9152 18050 9208
rect 18106 9152 18111 9208
rect 16021 9150 18111 9152
rect 16021 9147 16087 9150
rect 18045 9147 18111 9150
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 200 8258 800 8288
rect 1761 8258 1827 8261
rect 200 8256 1827 8258
rect 200 8200 1766 8256
rect 1822 8200 1827 8256
rect 200 8198 1827 8200
rect 200 8168 800 8198
rect 1761 8195 1827 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 5993 6898 6059 6901
rect 18873 6898 18939 6901
rect 5993 6896 18939 6898
rect 5993 6840 5998 6896
rect 6054 6840 18878 6896
rect 18934 6840 18939 6896
rect 5993 6838 18939 6840
rect 5993 6835 6059 6838
rect 18873 6835 18939 6838
rect 38193 6898 38259 6901
rect 39200 6898 39800 6928
rect 38193 6896 39800 6898
rect 38193 6840 38198 6896
rect 38254 6840 39800 6896
rect 38193 6838 39800 6840
rect 38193 6835 38259 6838
rect 39200 6808 39800 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 200 6218 800 6248
rect 1761 6218 1827 6221
rect 200 6216 1827 6218
rect 200 6160 1766 6216
rect 1822 6160 1827 6216
rect 200 6158 1827 6160
rect 200 6128 800 6158
rect 1761 6155 1827 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 5717 5674 5783 5677
rect 16573 5674 16639 5677
rect 5717 5672 16639 5674
rect 5717 5616 5722 5672
rect 5778 5616 16578 5672
rect 16634 5616 16639 5672
rect 5717 5614 16639 5616
rect 5717 5611 5783 5614
rect 16573 5611 16639 5614
rect 37181 5538 37247 5541
rect 39200 5538 39800 5568
rect 37181 5536 39800 5538
rect 37181 5480 37186 5536
rect 37242 5480 39800 5536
rect 37181 5478 39800 5480
rect 37181 5475 37247 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1761 4858 1827 4861
rect 200 4856 1827 4858
rect 200 4800 1766 4856
rect 1822 4800 1827 4856
rect 200 4798 1827 4800
rect 200 4768 800 4798
rect 1761 4795 1827 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 38193 3498 38259 3501
rect 39200 3498 39800 3528
rect 38193 3496 39800 3498
rect 38193 3440 38198 3496
rect 38254 3440 39800 3496
rect 38193 3438 39800 3440
rect 38193 3435 38259 3438
rect 39200 3408 39800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 200 2818 800 2848
rect 1761 2818 1827 2821
rect 200 2816 1827 2818
rect 200 2760 1766 2816
rect 1822 2760 1827 2816
rect 200 2758 1827 2760
rect 200 2728 800 2758
rect 1761 2755 1827 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 36905 2138 36971 2141
rect 39200 2138 39800 2168
rect 36905 2136 39800 2138
rect 36905 2080 36910 2136
rect 36966 2080 39800 2136
rect 36905 2078 39800 2080
rect 36905 2075 36971 2078
rect 39200 2048 39800 2078
rect 200 1458 800 1488
rect 2773 1458 2839 1461
rect 200 1456 2839 1458
rect 200 1400 2778 1456
rect 2834 1400 2839 1456
rect 200 1398 2839 1400
rect 200 1368 800 1398
rect 2773 1395 2839 1398
rect 38193 98 38259 101
rect 39200 98 39800 128
rect 38193 96 39800 98
rect 38193 40 38198 96
rect 38254 40 39800 96
rect 38193 38 39800 40
rect 38193 35 38259 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 2084 31724 2148 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 20116 25196 20180 25260
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 2084 23156 2148 23220
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 20668 20708 20732 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 20116 16492 20180 16556
rect 20668 16492 20732 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 2083 31788 2149 31789
rect 2083 31724 2084 31788
rect 2148 31724 2149 31788
rect 2083 31723 2149 31724
rect 2086 23221 2146 31723
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 2083 23220 2149 23221
rect 2083 23156 2084 23220
rect 2148 23156 2149 23220
rect 2083 23155 2149 23156
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 20115 25260 20181 25261
rect 20115 25196 20116 25260
rect 20180 25196 20181 25260
rect 20115 25195 20181 25196
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 20118 16557 20178 25195
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 20667 20772 20733 20773
rect 20667 20708 20668 20772
rect 20732 20708 20733 20772
rect 20667 20707 20733 20708
rect 20670 16557 20730 20707
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 20115 16556 20181 16557
rect 20115 16492 20116 16556
rect 20180 16492 20181 16556
rect 20115 16491 20181 16492
rect 20667 16556 20733 16557
rect 20667 16492 20668 16556
rect 20732 16492 20733 16556
rect 20667 16491 20733 16492
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 8648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform -1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 20332 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform 1 0 19780 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1667941163
transform 1 0 5520 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20
timestamp 1667941163
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71
timestamp 1667941163
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1667941163
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1667941163
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1667941163
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1667941163
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 1667941163
transform 1 0 14628 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_155
timestamp 1667941163
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1667941163
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_175
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1667941163
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1667941163
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_210
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_238
timestamp 1667941163
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1667941163
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 1667941163
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1667941163
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_322
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1667941163
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_342
timestamp 1667941163
transform 1 0 32568 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 1667941163
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1667941163
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 1667941163
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_399
timestamp 1667941163
transform 1 0 37812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_16
timestamp 1667941163
transform 1 0 2576 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_28
timestamp 1667941163
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_40
timestamp 1667941163
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1667941163
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_62
timestamp 1667941163
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_74
timestamp 1667941163
transform 1 0 7912 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1667941163
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_90
timestamp 1667941163
transform 1 0 9384 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_94
timestamp 1667941163
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1667941163
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_131
timestamp 1667941163
transform 1 0 13156 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_135
timestamp 1667941163
transform 1 0 13524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_147
timestamp 1667941163
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1667941163
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1667941163
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_194
timestamp 1667941163
transform 1 0 18952 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_206
timestamp 1667941163
transform 1 0 20056 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1667941163
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1667941163
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1667941163
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 1667941163
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_61
timestamp 1667941163
transform 1 0 6716 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1667941163
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1667941163
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_112
timestamp 1667941163
transform 1 0 11408 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_124
timestamp 1667941163
transform 1 0 12512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1667941163
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_185
timestamp 1667941163
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1667941163
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_123
timestamp 1667941163
transform 1 0 12420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_135
timestamp 1667941163
transform 1 0 13524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_147
timestamp 1667941163
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp 1667941163
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_174
timestamp 1667941163
transform 1 0 17112 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_186
timestamp 1667941163
transform 1 0 18216 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_198
timestamp 1667941163
transform 1 0 19320 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_210
timestamp 1667941163
transform 1 0 20424 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_112
timestamp 1667941163
transform 1 0 11408 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_116
timestamp 1667941163
transform 1 0 11776 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_120
timestamp 1667941163
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp 1667941163
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_183
timestamp 1667941163
transform 1 0 17940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_292
timestamp 1667941163
transform 1 0 27968 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1667941163
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1667941163
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1667941163
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1667941163
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_75
timestamp 1667941163
transform 1 0 8004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_87
timestamp 1667941163
transform 1 0 9108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_95
timestamp 1667941163
transform 1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1667941163
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_118
timestamp 1667941163
transform 1 0 11960 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_130
timestamp 1667941163
transform 1 0 13064 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_141
timestamp 1667941163
transform 1 0 14076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_153
timestamp 1667941163
transform 1 0 15180 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_157
timestamp 1667941163
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1667941163
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp 1667941163
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_342
timestamp 1667941163
transform 1 0 32568 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_354
timestamp 1667941163
transform 1 0 33672 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_366
timestamp 1667941163
transform 1 0 34776 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_378
timestamp 1667941163
transform 1 0 35880 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1667941163
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_36
timestamp 1667941163
transform 1 0 4416 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_43
timestamp 1667941163
transform 1 0 5060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_55
timestamp 1667941163
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_59
timestamp 1667941163
transform 1 0 6532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_68
timestamp 1667941163
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1667941163
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_124
timestamp 1667941163
transform 1 0 12512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1667941163
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_151
timestamp 1667941163
transform 1 0 14996 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_159
timestamp 1667941163
transform 1 0 15732 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1667941163
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_170
timestamp 1667941163
transform 1 0 16744 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_182
timestamp 1667941163
transform 1 0 17848 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_190
timestamp 1667941163
transform 1 0 18584 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_217
timestamp 1667941163
transform 1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_222
timestamp 1667941163
transform 1 0 21528 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_234
timestamp 1667941163
transform 1 0 22632 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_246
timestamp 1667941163
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_314
timestamp 1667941163
transform 1 0 29992 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_326
timestamp 1667941163
transform 1 0 31096 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_338
timestamp 1667941163
transform 1 0 32200 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_350
timestamp 1667941163
transform 1 0 33304 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1667941163
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_16
timestamp 1667941163
transform 1 0 2576 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_28
timestamp 1667941163
transform 1 0 3680 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_43
timestamp 1667941163
transform 1 0 5060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_63
timestamp 1667941163
transform 1 0 6900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_67
timestamp 1667941163
transform 1 0 7268 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_71
timestamp 1667941163
transform 1 0 7636 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1667941163
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_92
timestamp 1667941163
transform 1 0 9568 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_99
timestamp 1667941163
transform 1 0 10212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_122
timestamp 1667941163
transform 1 0 12328 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_128
timestamp 1667941163
transform 1 0 12880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_132
timestamp 1667941163
transform 1 0 13248 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_138
timestamp 1667941163
transform 1 0 13800 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_142
timestamp 1667941163
transform 1 0 14168 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1667941163
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_178
timestamp 1667941163
transform 1 0 17480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_182
timestamp 1667941163
transform 1 0 17848 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_201
timestamp 1667941163
transform 1 0 19596 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_212
timestamp 1667941163
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_241
timestamp 1667941163
transform 1 0 23276 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_245
timestamp 1667941163
transform 1 0 23644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_257
timestamp 1667941163
transform 1 0 24748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_265
timestamp 1667941163
transform 1 0 25484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_270
timestamp 1667941163
transform 1 0 25944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1667941163
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_37
timestamp 1667941163
transform 1 0 4508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_42
timestamp 1667941163
transform 1 0 4968 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_50
timestamp 1667941163
transform 1 0 5704 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_55
timestamp 1667941163
transform 1 0 6164 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_62
timestamp 1667941163
transform 1 0 6808 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_69
timestamp 1667941163
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1667941163
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_96
timestamp 1667941163
transform 1 0 9936 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_108
timestamp 1667941163
transform 1 0 11040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_114
timestamp 1667941163
transform 1 0 11592 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_123
timestamp 1667941163
transform 1 0 12420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1667941163
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_159
timestamp 1667941163
transform 1 0 15732 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_166
timestamp 1667941163
transform 1 0 16376 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1667941163
transform 1 0 17480 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_208
timestamp 1667941163
transform 1 0 20240 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_220
timestamp 1667941163
transform 1 0 21344 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_226
timestamp 1667941163
transform 1 0 21896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1667941163
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_242
timestamp 1667941163
transform 1 0 23368 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1667941163
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_259
timestamp 1667941163
transform 1 0 24932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_263
timestamp 1667941163
transform 1 0 25300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_275
timestamp 1667941163
transform 1 0 26404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_287
timestamp 1667941163
transform 1 0 27508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_299
timestamp 1667941163
transform 1 0 28612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_39
timestamp 1667941163
transform 1 0 4692 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_43
timestamp 1667941163
transform 1 0 5060 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_87
timestamp 1667941163
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_91
timestamp 1667941163
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1667941163
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_124
timestamp 1667941163
transform 1 0 12512 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_131
timestamp 1667941163
transform 1 0 13156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1667941163
transform 1 0 14260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_148
timestamp 1667941163
transform 1 0 14720 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1667941163
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1667941163
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp 1667941163
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_204
timestamp 1667941163
transform 1 0 19872 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1667941163
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_230
timestamp 1667941163
transform 1 0 22264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_241
timestamp 1667941163
transform 1 0 23276 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 1667941163
transform 1 0 23644 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_257
timestamp 1667941163
transform 1 0 24748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1667941163
transform 1 0 25852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1667941163
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_48
timestamp 1667941163
transform 1 0 5520 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_60
timestamp 1667941163
transform 1 0 6624 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_72
timestamp 1667941163
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1667941163
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_95
timestamp 1667941163
transform 1 0 9844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1667941163
transform 1 0 10488 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1667941163
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_129
timestamp 1667941163
transform 1 0 12972 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_160
timestamp 1667941163
transform 1 0 15824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_173
timestamp 1667941163
transform 1 0 17020 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1667941163
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_188
timestamp 1667941163
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1667941163
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_264
timestamp 1667941163
transform 1 0 25392 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1667941163
transform 1 0 26496 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_280
timestamp 1667941163
transform 1 0 26864 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_292
timestamp 1667941163
transform 1 0 27968 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 1667941163
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_9
timestamp 1667941163
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_21
timestamp 1667941163
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_33
timestamp 1667941163
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_45
timestamp 1667941163
transform 1 0 5244 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_62
timestamp 1667941163
transform 1 0 6808 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_74
timestamp 1667941163
transform 1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1667941163
transform 1 0 13156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1667941163
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1667941163
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_174
timestamp 1667941163
transform 1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_186
timestamp 1667941163
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_202
timestamp 1667941163
transform 1 0 19688 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp 1667941163
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1667941163
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_233
timestamp 1667941163
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_239
timestamp 1667941163
transform 1 0 23092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1667941163
transform 1 0 23460 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_247
timestamp 1667941163
transform 1 0 23828 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_259
timestamp 1667941163
transform 1 0 24932 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_269
timestamp 1667941163
transform 1 0 25852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1667941163
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_40
timestamp 1667941163
transform 1 0 4784 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_49
timestamp 1667941163
transform 1 0 5612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_56
timestamp 1667941163
transform 1 0 6256 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_63
timestamp 1667941163
transform 1 0 6900 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_71
timestamp 1667941163
transform 1 0 7636 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1667941163
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_156
timestamp 1667941163
transform 1 0 15456 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1667941163
transform 1 0 16100 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1667941163
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_190
timestamp 1667941163
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_216
timestamp 1667941163
transform 1 0 20976 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 1667941163
transform 1 0 21712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_235
timestamp 1667941163
transform 1 0 22724 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1667941163
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_261
timestamp 1667941163
transform 1 0 25116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_271
timestamp 1667941163
transform 1 0 26036 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_275
timestamp 1667941163
transform 1 0 26404 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_290
timestamp 1667941163
transform 1 0 27784 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1667941163
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_25
timestamp 1667941163
transform 1 0 3404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_29
timestamp 1667941163
transform 1 0 3772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1667941163
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_61
timestamp 1667941163
transform 1 0 6716 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_83
timestamp 1667941163
transform 1 0 8740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_138
timestamp 1667941163
transform 1 0 13800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1667941163
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_173
timestamp 1667941163
transform 1 0 17020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_183
timestamp 1667941163
transform 1 0 17940 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_190
timestamp 1667941163
transform 1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_197
timestamp 1667941163
transform 1 0 19228 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_204
timestamp 1667941163
transform 1 0 19872 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1667941163
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1667941163
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_234
timestamp 1667941163
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_238
timestamp 1667941163
transform 1 0 23000 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_246
timestamp 1667941163
transform 1 0 23736 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_257
timestamp 1667941163
transform 1 0 24748 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_264
timestamp 1667941163
transform 1 0 25392 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1667941163
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1667941163
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_301
timestamp 1667941163
transform 1 0 28796 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_306
timestamp 1667941163
transform 1 0 29256 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_318
timestamp 1667941163
transform 1 0 30360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1667941163
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_34
timestamp 1667941163
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1667941163
transform 1 0 5336 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_70
timestamp 1667941163
transform 1 0 7544 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1667941163
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_115
timestamp 1667941163
transform 1 0 11684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_127
timestamp 1667941163
transform 1 0 12788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_184
timestamp 1667941163
transform 1 0 18032 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1667941163
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_205
timestamp 1667941163
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_214
timestamp 1667941163
transform 1 0 20792 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_222
timestamp 1667941163
transform 1 0 21528 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_232
timestamp 1667941163
transform 1 0 22448 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_238
timestamp 1667941163
transform 1 0 23000 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_242
timestamp 1667941163
transform 1 0 23368 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1667941163
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_264
timestamp 1667941163
transform 1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_330
timestamp 1667941163
transform 1 0 31464 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_342
timestamp 1667941163
transform 1 0 32568 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_349
timestamp 1667941163
transform 1 0 33212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1667941163
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1667941163
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_63
timestamp 1667941163
transform 1 0 6900 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_85
timestamp 1667941163
transform 1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_97
timestamp 1667941163
transform 1 0 10028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1667941163
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_158
timestamp 1667941163
transform 1 0 15640 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_162
timestamp 1667941163
transform 1 0 16008 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1667941163
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_189
timestamp 1667941163
transform 1 0 18492 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_195
timestamp 1667941163
transform 1 0 19044 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_245
timestamp 1667941163
transform 1 0 23644 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_252
timestamp 1667941163
transform 1 0 24288 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_259
timestamp 1667941163
transform 1 0 24932 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_266
timestamp 1667941163
transform 1 0 25576 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1667941163
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_286
timestamp 1667941163
transform 1 0 27416 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_298
timestamp 1667941163
transform 1 0 28520 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_310
timestamp 1667941163
transform 1 0 29624 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_322
timestamp 1667941163
transform 1 0 30728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1667941163
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1667941163
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_401
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_63
timestamp 1667941163
transform 1 0 6900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1667941163
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_119
timestamp 1667941163
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1667941163
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1667941163
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1667941163
transform 1 0 15272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_161
timestamp 1667941163
transform 1 0 15916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_171
timestamp 1667941163
transform 1 0 16836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_186
timestamp 1667941163
transform 1 0 18216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1667941163
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_202
timestamp 1667941163
transform 1 0 19688 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1667941163
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_226
timestamp 1667941163
transform 1 0 21896 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_234
timestamp 1667941163
transform 1 0 22632 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_238
timestamp 1667941163
transform 1 0 23000 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_257
timestamp 1667941163
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_266
timestamp 1667941163
transform 1 0 25576 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_273
timestamp 1667941163
transform 1 0 26220 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_285
timestamp 1667941163
transform 1 0 27324 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_292
timestamp 1667941163
transform 1 0 27968 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1667941163
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_327
timestamp 1667941163
transform 1 0 31188 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_331
timestamp 1667941163
transform 1 0 31556 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_343
timestamp 1667941163
transform 1 0 32660 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_355
timestamp 1667941163
transform 1 0 33764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_75
timestamp 1667941163
transform 1 0 8004 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_96
timestamp 1667941163
transform 1 0 9936 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1667941163
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1667941163
transform 1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_140
timestamp 1667941163
transform 1 0 13984 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_146
timestamp 1667941163
transform 1 0 14536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp 1667941163
transform 1 0 14904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_157
timestamp 1667941163
transform 1 0 15548 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1667941163
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1667941163
transform 1 0 18492 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_202
timestamp 1667941163
transform 1 0 19688 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1667941163
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_248
timestamp 1667941163
transform 1 0 23920 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_260
timestamp 1667941163
transform 1 0 25024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_291
timestamp 1667941163
transform 1 0 27876 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_303
timestamp 1667941163
transform 1 0 28980 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_315
timestamp 1667941163
transform 1 0 30084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_327
timestamp 1667941163
transform 1 0 31188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_342
timestamp 1667941163
transform 1 0 32568 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_354
timestamp 1667941163
transform 1 0 33672 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_366
timestamp 1667941163
transform 1 0 34776 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_378
timestamp 1667941163
transform 1 0 35880 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1667941163
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_401
timestamp 1667941163
transform 1 0 37996 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_21
timestamp 1667941163
transform 1 0 3036 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1667941163
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_75
timestamp 1667941163
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_116
timestamp 1667941163
transform 1 0 11776 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_124
timestamp 1667941163
transform 1 0 12512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_128
timestamp 1667941163
transform 1 0 12880 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_134
timestamp 1667941163
transform 1 0 13432 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1667941163
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_170
timestamp 1667941163
transform 1 0 16744 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_179
timestamp 1667941163
transform 1 0 17572 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_185
timestamp 1667941163
transform 1 0 18124 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_205
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1667941163
transform 1 0 20884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1667941163
transform 1 0 21252 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_223
timestamp 1667941163
transform 1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_230
timestamp 1667941163
transform 1 0 22264 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1667941163
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_244
timestamp 1667941163
transform 1 0 23552 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_270
timestamp 1667941163
transform 1 0 25944 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_282
timestamp 1667941163
transform 1 0 27048 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_294
timestamp 1667941163
transform 1 0 28152 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1667941163
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_340
timestamp 1667941163
transform 1 0 32384 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_352
timestamp 1667941163
transform 1 0 33488 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_36
timestamp 1667941163
transform 1 0 4416 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1667941163
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1667941163
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_91
timestamp 1667941163
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1667941163
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp 1667941163
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_153
timestamp 1667941163
transform 1 0 15180 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1667941163
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1667941163
transform 1 0 18032 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_190
timestamp 1667941163
transform 1 0 18584 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_194
timestamp 1667941163
transform 1 0 18952 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_206
timestamp 1667941163
transform 1 0 20056 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_212
timestamp 1667941163
transform 1 0 20608 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_236
timestamp 1667941163
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_243
timestamp 1667941163
transform 1 0 23460 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_251
timestamp 1667941163
transform 1 0 24196 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_256
timestamp 1667941163
transform 1 0 24656 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_263
timestamp 1667941163
transform 1 0 25300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_270
timestamp 1667941163
transform 1 0 25944 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1667941163
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1667941163
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_9
timestamp 1667941163
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1667941163
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1667941163
transform 1 0 9660 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_115
timestamp 1667941163
transform 1 0 11684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_127
timestamp 1667941163
transform 1 0 12788 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_131
timestamp 1667941163
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1667941163
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_154
timestamp 1667941163
transform 1 0 15272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1667941163
transform 1 0 15640 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_162
timestamp 1667941163
transform 1 0 16008 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_174
timestamp 1667941163
transform 1 0 17112 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_182
timestamp 1667941163
transform 1 0 17848 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1667941163
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_207
timestamp 1667941163
transform 1 0 20148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_219
timestamp 1667941163
transform 1 0 21252 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_225
timestamp 1667941163
transform 1 0 21804 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1667941163
transform 1 0 22908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_241
timestamp 1667941163
transform 1 0 23276 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_260
timestamp 1667941163
transform 1 0 25024 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_272
timestamp 1667941163
transform 1 0 26128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_286
timestamp 1667941163
transform 1 0 27416 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_297
timestamp 1667941163
transform 1 0 28428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1667941163
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_315
timestamp 1667941163
transform 1 0 30084 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_327
timestamp 1667941163
transform 1 0 31188 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_339
timestamp 1667941163
transform 1 0 32292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_351
timestamp 1667941163
transform 1 0 33396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_37
timestamp 1667941163
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1667941163
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_157
timestamp 1667941163
transform 1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_182
timestamp 1667941163
transform 1 0 17848 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_190
timestamp 1667941163
transform 1 0 18584 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_201
timestamp 1667941163
transform 1 0 19596 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_208
timestamp 1667941163
transform 1 0 20240 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1667941163
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_250
timestamp 1667941163
transform 1 0 24104 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_257
timestamp 1667941163
transform 1 0 24748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_269
timestamp 1667941163
transform 1 0 25852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1667941163
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_286
timestamp 1667941163
transform 1 0 27416 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_294
timestamp 1667941163
transform 1 0 28152 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_298
timestamp 1667941163
transform 1 0 28520 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_310
timestamp 1667941163
transform 1 0 29624 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_322
timestamp 1667941163
transform 1 0 30728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1667941163
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_401
timestamp 1667941163
transform 1 0 37996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_15
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_35
timestamp 1667941163
transform 1 0 4324 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_61
timestamp 1667941163
transform 1 0 6716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1667941163
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1667941163
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 1667941163
transform 1 0 9292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_110
timestamp 1667941163
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_117
timestamp 1667941163
transform 1 0 11868 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_129
timestamp 1667941163
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1667941163
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 1667941163
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_151
timestamp 1667941163
transform 1 0 14996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_158
timestamp 1667941163
transform 1 0 15640 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_164
timestamp 1667941163
transform 1 0 16192 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_178
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1667941163
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_201
timestamp 1667941163
transform 1 0 19596 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_211
timestamp 1667941163
transform 1 0 20516 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1667941163
transform 1 0 21252 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1667941163
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1667941163
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_237
timestamp 1667941163
transform 1 0 22908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1667941163
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_269
timestamp 1667941163
transform 1 0 25852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_276
timestamp 1667941163
transform 1 0 26496 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_284
timestamp 1667941163
transform 1 0 27232 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_288
timestamp 1667941163
transform 1 0 27600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_300
timestamp 1667941163
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1667941163
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_31
timestamp 1667941163
transform 1 0 3956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_38
timestamp 1667941163
transform 1 0 4600 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1667941163
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1667941163
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_92
timestamp 1667941163
transform 1 0 9568 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1667941163
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_160
timestamp 1667941163
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_180
timestamp 1667941163
transform 1 0 17664 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_192
timestamp 1667941163
transform 1 0 18768 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_207
timestamp 1667941163
transform 1 0 20148 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1667941163
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_230
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_242
timestamp 1667941163
transform 1 0 23368 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_254
timestamp 1667941163
transform 1 0 24472 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_265
timestamp 1667941163
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1667941163
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_286
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_294
timestamp 1667941163
transform 1 0 28152 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_299
timestamp 1667941163
transform 1 0 28612 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_306
timestamp 1667941163
transform 1 0 29256 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_318
timestamp 1667941163
transform 1 0 30360 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1667941163
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_34
timestamp 1667941163
transform 1 0 4232 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_46
timestamp 1667941163
transform 1 0 5336 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_58
timestamp 1667941163
transform 1 0 6440 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_70
timestamp 1667941163
transform 1 0 7544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_105
timestamp 1667941163
transform 1 0 10764 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1667941163
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_146
timestamp 1667941163
transform 1 0 14536 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1667941163
transform 1 0 15640 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1667941163
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_169
timestamp 1667941163
transform 1 0 16652 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1667941163
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_185
timestamp 1667941163
transform 1 0 18124 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 1667941163
transform 1 0 19596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_211
timestamp 1667941163
transform 1 0 20516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_223
timestamp 1667941163
transform 1 0 21620 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_231
timestamp 1667941163
transform 1 0 22356 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_237
timestamp 1667941163
transform 1 0 22908 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_245
timestamp 1667941163
transform 1 0 23644 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_263
timestamp 1667941163
transform 1 0 25300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_283
timestamp 1667941163
transform 1 0 27140 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_293
timestamp 1667941163
transform 1 0 28060 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_300
timestamp 1667941163
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_314
timestamp 1667941163
transform 1 0 29992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_328
timestamp 1667941163
transform 1 0 31280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_335
timestamp 1667941163
transform 1 0 31924 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_342
timestamp 1667941163
transform 1 0 32568 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 1667941163
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1667941163
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_28
timestamp 1667941163
transform 1 0 3680 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_40
timestamp 1667941163
transform 1 0 4784 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1667941163
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1667941163
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_148
timestamp 1667941163
transform 1 0 14720 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1667941163
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp 1667941163
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1667941163
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_198
timestamp 1667941163
transform 1 0 19320 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_204
timestamp 1667941163
transform 1 0 19872 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_208
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1667941163
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_241
timestamp 1667941163
transform 1 0 23276 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_245
timestamp 1667941163
transform 1 0 23644 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1667941163
transform 1 0 24472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_268
timestamp 1667941163
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_8
timestamp 1667941163
transform 1 0 1840 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_20
timestamp 1667941163
transform 1 0 2944 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_49
timestamp 1667941163
transform 1 0 5612 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_73
timestamp 1667941163
transform 1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1667941163
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_120
timestamp 1667941163
transform 1 0 12144 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_126
timestamp 1667941163
transform 1 0 12696 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_130
timestamp 1667941163
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_157
timestamp 1667941163
transform 1 0 15548 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_170
timestamp 1667941163
transform 1 0 16744 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_182
timestamp 1667941163
transform 1 0 17848 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_186
timestamp 1667941163
transform 1 0 18216 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1667941163
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_215
timestamp 1667941163
transform 1 0 20884 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_219
timestamp 1667941163
transform 1 0 21252 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_231
timestamp 1667941163
transform 1 0 22356 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1667941163
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_262
timestamp 1667941163
transform 1 0 25208 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_268
timestamp 1667941163
transform 1 0 25760 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_272
timestamp 1667941163
transform 1 0 26128 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_279
timestamp 1667941163
transform 1 0 26772 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_286
timestamp 1667941163
transform 1 0 27416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_298
timestamp 1667941163
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1667941163
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_317
timestamp 1667941163
transform 1 0 30268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_327
timestamp 1667941163
transform 1 0 31188 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_335
timestamp 1667941163
transform 1 0 31924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_342
timestamp 1667941163
transform 1 0 32568 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_350
timestamp 1667941163
transform 1 0 33304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_355
timestamp 1667941163
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_65
timestamp 1667941163
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_89
timestamp 1667941163
transform 1 0 9292 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_101
timestamp 1667941163
transform 1 0 10396 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1667941163
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_131
timestamp 1667941163
transform 1 0 13156 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_153
timestamp 1667941163
transform 1 0 15180 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_179
timestamp 1667941163
transform 1 0 17572 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_188
timestamp 1667941163
transform 1 0 18400 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_201
timestamp 1667941163
transform 1 0 19596 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_213
timestamp 1667941163
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1667941163
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_241
timestamp 1667941163
transform 1 0 23276 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_253
timestamp 1667941163
transform 1 0 24380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_265
timestamp 1667941163
transform 1 0 25484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_298
timestamp 1667941163
transform 1 0 28520 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_310
timestamp 1667941163
transform 1 0 29624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_315
timestamp 1667941163
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_322
timestamp 1667941163
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1667941163
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_347
timestamp 1667941163
transform 1 0 33028 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_359
timestamp 1667941163
transform 1 0 34132 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_371
timestamp 1667941163
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_383
timestamp 1667941163
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_401
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_58
timestamp 1667941163
transform 1 0 6440 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_70
timestamp 1667941163
transform 1 0 7544 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_108
timestamp 1667941163
transform 1 0 11040 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_120
timestamp 1667941163
transform 1 0 12144 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1667941163
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_152
timestamp 1667941163
transform 1 0 15088 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_158
timestamp 1667941163
transform 1 0 15640 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_162
timestamp 1667941163
transform 1 0 16008 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_169
timestamp 1667941163
transform 1 0 16652 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1667941163
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_205
timestamp 1667941163
transform 1 0 19964 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_217
timestamp 1667941163
transform 1 0 21068 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_225
timestamp 1667941163
transform 1 0 21804 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1667941163
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_242
timestamp 1667941163
transform 1 0 23368 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1667941163
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_259
timestamp 1667941163
transform 1 0 24932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_263
timestamp 1667941163
transform 1 0 25300 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_271
timestamp 1667941163
transform 1 0 26036 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_280
timestamp 1667941163
transform 1 0 26864 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_288
timestamp 1667941163
transform 1 0 27600 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_297
timestamp 1667941163
transform 1 0 28428 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1667941163
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_314
timestamp 1667941163
transform 1 0 29992 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_326
timestamp 1667941163
transform 1 0 31096 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_338
timestamp 1667941163
transform 1 0 32200 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_350
timestamp 1667941163
transform 1 0 33304 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1667941163
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_8
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_12
timestamp 1667941163
transform 1 0 2208 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_34
timestamp 1667941163
transform 1 0 4232 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_46
timestamp 1667941163
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1667941163
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_148
timestamp 1667941163
transform 1 0 14720 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_160
timestamp 1667941163
transform 1 0 15824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_178
timestamp 1667941163
transform 1 0 17480 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_190
timestamp 1667941163
transform 1 0 18584 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_202
timestamp 1667941163
transform 1 0 19688 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_211
timestamp 1667941163
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp 1667941163
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_231
timestamp 1667941163
transform 1 0 22356 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_240
timestamp 1667941163
transform 1 0 23184 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_248
timestamp 1667941163
transform 1 0 23920 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1667941163
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1667941163
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_309
timestamp 1667941163
transform 1 0 29532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1667941163
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_320
timestamp 1667941163
transform 1 0 30544 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 1667941163
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_11
timestamp 1667941163
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_17
timestamp 1667941163
transform 1 0 2668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1667941163
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_55
timestamp 1667941163
transform 1 0 6164 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1667941163
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_123
timestamp 1667941163
transform 1 0 12420 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1667941163
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1667941163
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1667941163
transform 1 0 15272 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp 1667941163
transform 1 0 15916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_174
timestamp 1667941163
transform 1 0 17112 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1667941163
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_204
timestamp 1667941163
transform 1 0 19872 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_215
timestamp 1667941163
transform 1 0 20884 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_227
timestamp 1667941163
transform 1 0 21988 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_237
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1667941163
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_261
timestamp 1667941163
transform 1 0 25116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_267
timestamp 1667941163
transform 1 0 25668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_274
timestamp 1667941163
transform 1 0 26312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_281
timestamp 1667941163
transform 1 0 26956 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1667941163
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_299
timestamp 1667941163
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_319
timestamp 1667941163
transform 1 0 30452 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_331
timestamp 1667941163
transform 1 0 31556 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_343
timestamp 1667941163
transform 1 0 32660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_354
timestamp 1667941163
transform 1 0 33672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1667941163
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_405
timestamp 1667941163
transform 1 0 38364 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_11
timestamp 1667941163
transform 1 0 2116 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1667941163
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1667941163
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1667941163
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_124
timestamp 1667941163
transform 1 0 12512 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_130
timestamp 1667941163
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_154
timestamp 1667941163
transform 1 0 15272 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_174
timestamp 1667941163
transform 1 0 17112 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_186
timestamp 1667941163
transform 1 0 18216 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_194
timestamp 1667941163
transform 1 0 18952 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_211
timestamp 1667941163
transform 1 0 20516 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1667941163
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_234
timestamp 1667941163
transform 1 0 22632 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_246
timestamp 1667941163
transform 1 0 23736 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_258
timestamp 1667941163
transform 1 0 24840 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_265
timestamp 1667941163
transform 1 0 25484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1667941163
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_292
timestamp 1667941163
transform 1 0 27968 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_304
timestamp 1667941163
transform 1 0 29072 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_316
timestamp 1667941163
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1667941163
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_8
timestamp 1667941163
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1667941163
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1667941163
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_59
timestamp 1667941163
transform 1 0 6532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_74
timestamp 1667941163
transform 1 0 7912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_111
timestamp 1667941163
transform 1 0 11316 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_118
timestamp 1667941163
transform 1 0 11960 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_130
timestamp 1667941163
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_149
timestamp 1667941163
transform 1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_155
timestamp 1667941163
transform 1 0 15364 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_167
timestamp 1667941163
transform 1 0 16468 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_179
timestamp 1667941163
transform 1 0 17572 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_183
timestamp 1667941163
transform 1 0 17940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_225
timestamp 1667941163
transform 1 0 21804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_229
timestamp 1667941163
transform 1 0 22172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1667941163
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1667941163
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_263
timestamp 1667941163
transform 1 0 25300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1667941163
transform 1 0 25944 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_293
timestamp 1667941163
transform 1 0 28060 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_303
timestamp 1667941163
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_320
timestamp 1667941163
transform 1 0 30544 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_332
timestamp 1667941163
transform 1 0 31648 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_344
timestamp 1667941163
transform 1 0 32752 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1667941163
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1667941163
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_10
timestamp 1667941163
transform 1 0 2024 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_22
timestamp 1667941163
transform 1 0 3128 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_34
timestamp 1667941163
transform 1 0 4232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1667941163
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_65
timestamp 1667941163
transform 1 0 7084 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_90
timestamp 1667941163
transform 1 0 9384 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1667941163
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1667941163
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_159
timestamp 1667941163
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1667941163
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_187
timestamp 1667941163
transform 1 0 18308 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1667941163
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_212
timestamp 1667941163
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_238
timestamp 1667941163
transform 1 0 23000 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_247
timestamp 1667941163
transform 1 0 23828 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_259
timestamp 1667941163
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1667941163
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_292
timestamp 1667941163
transform 1 0 27968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_304
timestamp 1667941163
transform 1 0 29072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_309
timestamp 1667941163
transform 1 0 29532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_321
timestamp 1667941163
transform 1 0 30636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_328
timestamp 1667941163
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_343
timestamp 1667941163
transform 1 0 32660 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_348
timestamp 1667941163
transform 1 0 33120 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_360
timestamp 1667941163
transform 1 0 34224 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_372
timestamp 1667941163
transform 1 0 35328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_384
timestamp 1667941163
transform 1 0 36432 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1667941163
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_51
timestamp 1667941163
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_63
timestamp 1667941163
transform 1 0 6900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_75
timestamp 1667941163
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_120
timestamp 1667941163
transform 1 0 12144 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 1667941163
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1667941163
transform 1 0 15088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_159
timestamp 1667941163
transform 1 0 15732 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_166
timestamp 1667941163
transform 1 0 16376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_173
timestamp 1667941163
transform 1 0 17020 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_204
timestamp 1667941163
transform 1 0 19872 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_216
timestamp 1667941163
transform 1 0 20976 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_227
timestamp 1667941163
transform 1 0 21988 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_235
timestamp 1667941163
transform 1 0 22724 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_239
timestamp 1667941163
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1667941163
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_283
timestamp 1667941163
transform 1 0 27140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_287
timestamp 1667941163
transform 1 0 27508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_299
timestamp 1667941163
transform 1 0 28612 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_314
timestamp 1667941163
transform 1 0 29992 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_322
timestamp 1667941163
transform 1 0 30728 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_327
timestamp 1667941163
transform 1 0 31188 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_339
timestamp 1667941163
transform 1 0 32292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_351
timestamp 1667941163
transform 1 0 33396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1667941163
transform 1 0 1840 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_20
timestamp 1667941163
transform 1 0 2944 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_32
timestamp 1667941163
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_44
timestamp 1667941163
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_80
timestamp 1667941163
transform 1 0 8464 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_84
timestamp 1667941163
transform 1 0 8832 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_96
timestamp 1667941163
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1667941163
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_141
timestamp 1667941163
transform 1 0 14076 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_148
timestamp 1667941163
transform 1 0 14720 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1667941163
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_174
timestamp 1667941163
transform 1 0 17112 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_194
timestamp 1667941163
transform 1 0 18952 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_209
timestamp 1667941163
transform 1 0 20332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1667941163
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_254
timestamp 1667941163
transform 1 0 24472 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_266
timestamp 1667941163
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_298
timestamp 1667941163
transform 1 0 28520 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_310
timestamp 1667941163
transform 1 0 29624 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_322
timestamp 1667941163
transform 1 0 30728 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_326
timestamp 1667941163
transform 1 0 31096 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1667941163
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1667941163
transform 1 0 9476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_95
timestamp 1667941163
transform 1 0 9844 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_101
timestamp 1667941163
transform 1 0 10396 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_125
timestamp 1667941163
transform 1 0 12604 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_166
timestamp 1667941163
transform 1 0 16376 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_174
timestamp 1667941163
transform 1 0 17112 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1667941163
transform 1 0 17572 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1667941163
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1667941163
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_219
timestamp 1667941163
transform 1 0 21252 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_227
timestamp 1667941163
transform 1 0 21988 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1667941163
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_258
timestamp 1667941163
transform 1 0 24840 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_270
timestamp 1667941163
transform 1 0 25944 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_274
timestamp 1667941163
transform 1 0 26312 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_282
timestamp 1667941163
transform 1 0 27048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_286
timestamp 1667941163
transform 1 0 27416 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_294
timestamp 1667941163
transform 1 0 28152 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1667941163
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_318
timestamp 1667941163
transform 1 0 30360 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_330
timestamp 1667941163
transform 1 0 31464 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_342
timestamp 1667941163
transform 1 0 32568 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_354
timestamp 1667941163
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_7
timestamp 1667941163
transform 1 0 1748 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_17
timestamp 1667941163
transform 1 0 2668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_29
timestamp 1667941163
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_41
timestamp 1667941163
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1667941163
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_73
timestamp 1667941163
transform 1 0 7820 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_80
timestamp 1667941163
transform 1 0 8464 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_107
timestamp 1667941163
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_158
timestamp 1667941163
transform 1 0 15640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_162
timestamp 1667941163
transform 1 0 16008 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_175
timestamp 1667941163
transform 1 0 17204 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_185
timestamp 1667941163
transform 1 0 18124 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_197
timestamp 1667941163
transform 1 0 19228 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_204
timestamp 1667941163
transform 1 0 19872 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_216
timestamp 1667941163
transform 1 0 20976 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_255
timestamp 1667941163
transform 1 0 24564 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_265
timestamp 1667941163
transform 1 0 25484 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_272
timestamp 1667941163
transform 1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1667941163
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_299
timestamp 1667941163
transform 1 0 28612 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_311
timestamp 1667941163
transform 1 0 29716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_323
timestamp 1667941163
transform 1 0 30820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_9
timestamp 1667941163
transform 1 0 1932 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1667941163
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_51
timestamp 1667941163
transform 1 0 5796 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_63
timestamp 1667941163
transform 1 0 6900 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1667941163
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_111
timestamp 1667941163
transform 1 0 11316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1667941163
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_147
timestamp 1667941163
transform 1 0 14628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_151
timestamp 1667941163
transform 1 0 14996 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_158
timestamp 1667941163
transform 1 0 15640 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_164
timestamp 1667941163
transform 1 0 16192 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_174
timestamp 1667941163
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_181
timestamp 1667941163
transform 1 0 17756 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_188
timestamp 1667941163
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_201
timestamp 1667941163
transform 1 0 19596 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_205
timestamp 1667941163
transform 1 0 19964 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_215
timestamp 1667941163
transform 1 0 20884 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_227
timestamp 1667941163
transform 1 0 21988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1667941163
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1667941163
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_261
timestamp 1667941163
transform 1 0 25116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_267
timestamp 1667941163
transform 1 0 25668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_275
timestamp 1667941163
transform 1 0 26404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_280
timestamp 1667941163
transform 1 0 26864 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_284
timestamp 1667941163
transform 1 0 27232 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_293
timestamp 1667941163
transform 1 0 28060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_300
timestamp 1667941163
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_29
timestamp 1667941163
transform 1 0 3772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_41
timestamp 1667941163
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1667941163
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_68
timestamp 1667941163
transform 1 0 7360 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_75
timestamp 1667941163
transform 1 0 8004 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_87
timestamp 1667941163
transform 1 0 9108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_99
timestamp 1667941163
transform 1 0 10212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_131
timestamp 1667941163
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_153
timestamp 1667941163
transform 1 0 15180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1667941163
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_174
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_185
timestamp 1667941163
transform 1 0 18124 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_189
timestamp 1667941163
transform 1 0 18492 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_198
timestamp 1667941163
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_211
timestamp 1667941163
transform 1 0 20516 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1667941163
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_230
timestamp 1667941163
transform 1 0 22264 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_238
timestamp 1667941163
transform 1 0 23000 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_244
timestamp 1667941163
transform 1 0 23552 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_256
timestamp 1667941163
transform 1 0 24656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_262
timestamp 1667941163
transform 1 0 25208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_292
timestamp 1667941163
transform 1 0 27968 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_299
timestamp 1667941163
transform 1 0 28612 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_320
timestamp 1667941163
transform 1 0 30544 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1667941163
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_401
timestamp 1667941163
transform 1 0 37996 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1667941163
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_34
timestamp 1667941163
transform 1 0 4232 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_40
timestamp 1667941163
transform 1 0 4784 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_61
timestamp 1667941163
transform 1 0 6716 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_73
timestamp 1667941163
transform 1 0 7820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 1667941163
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_90
timestamp 1667941163
transform 1 0 9384 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_102
timestamp 1667941163
transform 1 0 10488 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_114
timestamp 1667941163
transform 1 0 11592 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_126
timestamp 1667941163
transform 1 0 12696 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1667941163
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_149
timestamp 1667941163
transform 1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_157
timestamp 1667941163
transform 1 0 15548 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_162
timestamp 1667941163
transform 1 0 16008 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_169
timestamp 1667941163
transform 1 0 16652 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_181
timestamp 1667941163
transform 1 0 17756 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1667941163
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_220
timestamp 1667941163
transform 1 0 21344 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_235
timestamp 1667941163
transform 1 0 22724 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_242
timestamp 1667941163
transform 1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1667941163
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_261
timestamp 1667941163
transform 1 0 25116 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_285
timestamp 1667941163
transform 1 0 27324 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_291
timestamp 1667941163
transform 1 0 27876 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_298
timestamp 1667941163
transform 1 0 28520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1667941163
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_28
timestamp 1667941163
transform 1 0 3680 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_40
timestamp 1667941163
transform 1 0 4784 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1667941163
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1667941163
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_133
timestamp 1667941163
transform 1 0 13340 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_154
timestamp 1667941163
transform 1 0 15272 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_162
timestamp 1667941163
transform 1 0 16008 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_182
timestamp 1667941163
transform 1 0 17848 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_194
timestamp 1667941163
transform 1 0 18952 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_213
timestamp 1667941163
transform 1 0 20700 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_233
timestamp 1667941163
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1667941163
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1667941163
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_299
timestamp 1667941163
transform 1 0 28612 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_306
timestamp 1667941163
transform 1 0 29256 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_314
timestamp 1667941163
transform 1 0 29992 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_324
timestamp 1667941163
transform 1 0 30912 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_12
timestamp 1667941163
transform 1 0 2208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_19
timestamp 1667941163
transform 1 0 2852 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1667941163
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_40
timestamp 1667941163
transform 1 0 4784 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_52
timestamp 1667941163
transform 1 0 5888 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_64
timestamp 1667941163
transform 1 0 6992 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_76
timestamp 1667941163
transform 1 0 8096 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1667941163
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_107
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_119
timestamp 1667941163
transform 1 0 12052 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_131
timestamp 1667941163
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_168
timestamp 1667941163
transform 1 0 16560 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_180
timestamp 1667941163
transform 1 0 17664 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1667941163
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1667941163
transform 1 0 20240 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_212
timestamp 1667941163
transform 1 0 20608 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_216
timestamp 1667941163
transform 1 0 20976 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_228
timestamp 1667941163
transform 1 0 22080 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_234
timestamp 1667941163
transform 1 0 22632 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1667941163
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_258
timestamp 1667941163
transform 1 0 24840 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_270
timestamp 1667941163
transform 1 0 25944 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_285
timestamp 1667941163
transform 1 0 27324 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_292
timestamp 1667941163
transform 1 0 27968 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1667941163
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_342
timestamp 1667941163
transform 1 0 32568 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_349
timestamp 1667941163
transform 1 0 33212 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1667941163
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1667941163
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_16
timestamp 1667941163
transform 1 0 2576 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1667941163
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_134
timestamp 1667941163
transform 1 0 13432 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_146
timestamp 1667941163
transform 1 0 14536 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_158
timestamp 1667941163
transform 1 0 15640 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1667941163
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_175
timestamp 1667941163
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_192
timestamp 1667941163
transform 1 0 18768 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_211
timestamp 1667941163
transform 1 0 20516 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_215
timestamp 1667941163
transform 1 0 20884 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_242
timestamp 1667941163
transform 1 0 23368 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_254
timestamp 1667941163
transform 1 0 24472 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_266
timestamp 1667941163
transform 1 0 25576 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_274
timestamp 1667941163
transform 1 0 26312 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1667941163
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_291
timestamp 1667941163
transform 1 0 27876 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_299
timestamp 1667941163
transform 1 0 28612 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_304
timestamp 1667941163
transform 1 0 29072 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_311
timestamp 1667941163
transform 1 0 29716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_323
timestamp 1667941163
transform 1 0 30820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_7
timestamp 1667941163
transform 1 0 1748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_16
timestamp 1667941163
transform 1 0 2576 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_23
timestamp 1667941163
transform 1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_47
timestamp 1667941163
transform 1 0 5428 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_50
timestamp 1667941163
transform 1 0 5704 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_75
timestamp 1667941163
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1667941163
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_113
timestamp 1667941163
transform 1 0 11500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1667941163
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_163
timestamp 1667941163
transform 1 0 16100 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_170
timestamp 1667941163
transform 1 0 16744 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_174
timestamp 1667941163
transform 1 0 17112 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_184
timestamp 1667941163
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_208
timestamp 1667941163
transform 1 0 20240 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_220
timestamp 1667941163
transform 1 0 21344 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_234
timestamp 1667941163
transform 1 0 22632 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1667941163
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_258
timestamp 1667941163
transform 1 0 24840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_270
timestamp 1667941163
transform 1 0 25944 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_276
timestamp 1667941163
transform 1 0 26496 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_288
timestamp 1667941163
transform 1 0 27600 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_299
timestamp 1667941163
transform 1 0 28612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1667941163
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_7
timestamp 1667941163
transform 1 0 1748 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_12
timestamp 1667941163
transform 1 0 2208 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_24
timestamp 1667941163
transform 1 0 3312 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_32
timestamp 1667941163
transform 1 0 4048 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_37
timestamp 1667941163
transform 1 0 4508 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1667941163
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_98
timestamp 1667941163
transform 1 0 10120 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_150
timestamp 1667941163
transform 1 0 14904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_162
timestamp 1667941163
transform 1 0 16008 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_175
timestamp 1667941163
transform 1 0 17204 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_179
timestamp 1667941163
transform 1 0 17572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_191
timestamp 1667941163
transform 1 0 18676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_197
timestamp 1667941163
transform 1 0 19228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_201
timestamp 1667941163
transform 1 0 19596 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_209
timestamp 1667941163
transform 1 0 20332 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_215
timestamp 1667941163
transform 1 0 20884 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1667941163
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_264
timestamp 1667941163
transform 1 0 25392 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1667941163
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_290
timestamp 1667941163
transform 1 0 27784 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_302
timestamp 1667941163
transform 1 0 28888 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_314
timestamp 1667941163
transform 1 0 29992 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_326
timestamp 1667941163
transform 1 0 31096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1667941163
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_401
timestamp 1667941163
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_8
timestamp 1667941163
transform 1 0 1840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1667941163
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_40
timestamp 1667941163
transform 1 0 4784 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_48
timestamp 1667941163
transform 1 0 5520 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_59
timestamp 1667941163
transform 1 0 6532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_71
timestamp 1667941163
transform 1 0 7636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_105
timestamp 1667941163
transform 1 0 10764 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_128
timestamp 1667941163
transform 1 0 12880 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_161
timestamp 1667941163
transform 1 0 15916 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1667941163
transform 1 0 16468 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1667941163
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_181
timestamp 1667941163
transform 1 0 17756 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_185
timestamp 1667941163
transform 1 0 18124 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_207
timestamp 1667941163
transform 1 0 20148 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_214
timestamp 1667941163
transform 1 0 20792 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_223
timestamp 1667941163
transform 1 0 21620 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_235
timestamp 1667941163
transform 1 0 22724 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_241
timestamp 1667941163
transform 1 0 23276 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1667941163
transform 1 0 24840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_272
timestamp 1667941163
transform 1 0 26128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_279
timestamp 1667941163
transform 1 0 26772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_285
timestamp 1667941163
transform 1 0 27324 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_7
timestamp 1667941163
transform 1 0 1748 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_11
timestamp 1667941163
transform 1 0 2116 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_19
timestamp 1667941163
transform 1 0 2852 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_29
timestamp 1667941163
transform 1 0 3772 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_42
timestamp 1667941163
transform 1 0 4968 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1667941163
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_62
timestamp 1667941163
transform 1 0 6808 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_74
timestamp 1667941163
transform 1 0 7912 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_86
timestamp 1667941163
transform 1 0 9016 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_98
timestamp 1667941163
transform 1 0 10120 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1667941163
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_140
timestamp 1667941163
transform 1 0 13984 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_148
timestamp 1667941163
transform 1 0 14720 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_152
timestamp 1667941163
transform 1 0 15088 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_159
timestamp 1667941163
transform 1 0 15732 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_179
timestamp 1667941163
transform 1 0 17572 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_183
timestamp 1667941163
transform 1 0 17940 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_197
timestamp 1667941163
transform 1 0 19228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_201
timestamp 1667941163
transform 1 0 19596 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_213
timestamp 1667941163
transform 1 0 20700 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_230
timestamp 1667941163
transform 1 0 22264 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_239
timestamp 1667941163
transform 1 0 23092 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_253
timestamp 1667941163
transform 1 0 24380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_259
timestamp 1667941163
transform 1 0 24932 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_268
timestamp 1667941163
transform 1 0 25760 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_10
timestamp 1667941163
transform 1 0 2024 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_22
timestamp 1667941163
transform 1 0 3128 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_37
timestamp 1667941163
transform 1 0 4508 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_42
timestamp 1667941163
transform 1 0 4968 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_49
timestamp 1667941163
transform 1 0 5612 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_61
timestamp 1667941163
transform 1 0 6716 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_73
timestamp 1667941163
transform 1 0 7820 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1667941163
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_96
timestamp 1667941163
transform 1 0 9936 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_105
timestamp 1667941163
transform 1 0 10764 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_117
timestamp 1667941163
transform 1 0 11868 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_129
timestamp 1667941163
transform 1 0 12972 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_137
timestamp 1667941163
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1667941163
transform 1 0 14444 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_155
timestamp 1667941163
transform 1 0 15364 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_167
timestamp 1667941163
transform 1 0 16468 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_174
timestamp 1667941163
transform 1 0 17112 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_186
timestamp 1667941163
transform 1 0 18216 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1667941163
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_217
timestamp 1667941163
transform 1 0 21068 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_228
timestamp 1667941163
transform 1 0 22080 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_240
timestamp 1667941163
transform 1 0 23184 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_260
timestamp 1667941163
transform 1 0 25024 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_272
timestamp 1667941163
transform 1 0 26128 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_284
timestamp 1667941163
transform 1 0 27232 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_296
timestamp 1667941163
transform 1 0 28336 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_20
timestamp 1667941163
transform 1 0 2944 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_32
timestamp 1667941163
transform 1 0 4048 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1667941163
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_63
timestamp 1667941163
transform 1 0 6900 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_72
timestamp 1667941163
transform 1 0 7728 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_84
timestamp 1667941163
transform 1 0 8832 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_92
timestamp 1667941163
transform 1 0 9568 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_96
timestamp 1667941163
transform 1 0 9936 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_100
timestamp 1667941163
transform 1 0 10304 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1667941163
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_121
timestamp 1667941163
transform 1 0 12236 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_154
timestamp 1667941163
transform 1 0 15272 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1667941163
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_189
timestamp 1667941163
transform 1 0 18492 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_200
timestamp 1667941163
transform 1 0 19504 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_212
timestamp 1667941163
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_241
timestamp 1667941163
transform 1 0 23276 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_245
timestamp 1667941163
transform 1 0 23644 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_257
timestamp 1667941163
transform 1 0 24748 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_264
timestamp 1667941163
transform 1 0 25392 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1667941163
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_321
timestamp 1667941163
transform 1 0 30636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_333
timestamp 1667941163
transform 1 0 31740 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_7
timestamp 1667941163
transform 1 0 1748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_11
timestamp 1667941163
transform 1 0 2116 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1667941163
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_34
timestamp 1667941163
transform 1 0 4232 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_46
timestamp 1667941163
transform 1 0 5336 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_54
timestamp 1667941163
transform 1 0 6072 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_58
timestamp 1667941163
transform 1 0 6440 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_72
timestamp 1667941163
transform 1 0 7728 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_95
timestamp 1667941163
transform 1 0 9844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_107
timestamp 1667941163
transform 1 0 10948 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_119
timestamp 1667941163
transform 1 0 12052 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_132
timestamp 1667941163
transform 1 0 13248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_146
timestamp 1667941163
transform 1 0 14536 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_158
timestamp 1667941163
transform 1 0 15640 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_170
timestamp 1667941163
transform 1 0 16744 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1667941163
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_207
timestamp 1667941163
transform 1 0 20148 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1667941163
transform 1 0 20700 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_217
timestamp 1667941163
transform 1 0 21068 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_229
timestamp 1667941163
transform 1 0 22172 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_237
timestamp 1667941163
transform 1 0 22908 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_241
timestamp 1667941163
transform 1 0 23276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1667941163
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_8
timestamp 1667941163
transform 1 0 1840 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_16
timestamp 1667941163
transform 1 0 2576 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_20
timestamp 1667941163
transform 1 0 2944 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_32
timestamp 1667941163
transform 1 0 4048 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1667941163
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_61
timestamp 1667941163
transform 1 0 6716 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_71
timestamp 1667941163
transform 1 0 7636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_83
timestamp 1667941163
transform 1 0 8740 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_87
timestamp 1667941163
transform 1 0 9108 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_91
timestamp 1667941163
transform 1 0 9476 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_103
timestamp 1667941163
transform 1 0 10580 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1667941163
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_124
timestamp 1667941163
transform 1 0 12512 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_130
timestamp 1667941163
transform 1 0 13064 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_134
timestamp 1667941163
transform 1 0 13432 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_141
timestamp 1667941163
transform 1 0 14076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_153
timestamp 1667941163
transform 1 0 15180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1667941163
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_180
timestamp 1667941163
transform 1 0 17664 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_187
timestamp 1667941163
transform 1 0 18308 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_199
timestamp 1667941163
transform 1 0 19412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_211
timestamp 1667941163
transform 1 0 20516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_230
timestamp 1667941163
transform 1 0 22264 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_242
timestamp 1667941163
transform 1 0 23368 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_254
timestamp 1667941163
transform 1 0 24472 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_266
timestamp 1667941163
transform 1 0 25576 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1667941163
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1667941163
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_353
timestamp 1667941163
transform 1 0 33580 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_362
timestamp 1667941163
transform 1 0 34408 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_374
timestamp 1667941163
transform 1 0 35512 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_386
timestamp 1667941163
transform 1 0 36616 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_12
timestamp 1667941163
transform 1 0 2208 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_19
timestamp 1667941163
transform 1 0 2852 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1667941163
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_35
timestamp 1667941163
transform 1 0 4324 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_47
timestamp 1667941163
transform 1 0 5428 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_55
timestamp 1667941163
transform 1 0 6164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_67
timestamp 1667941163
transform 1 0 7268 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_71
timestamp 1667941163
transform 1 0 7636 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_75
timestamp 1667941163
transform 1 0 8004 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_91
timestamp 1667941163
transform 1 0 9476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_98
timestamp 1667941163
transform 1 0 10120 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_102
timestamp 1667941163
transform 1 0 10488 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_106
timestamp 1667941163
transform 1 0 10856 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_119
timestamp 1667941163
transform 1 0 12052 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_131
timestamp 1667941163
transform 1 0 13156 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_136
timestamp 1667941163
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_171
timestamp 1667941163
transform 1 0 16836 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_175
timestamp 1667941163
transform 1 0 17204 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_187
timestamp 1667941163
transform 1 0 18308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_203
timestamp 1667941163
transform 1 0 19780 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_210
timestamp 1667941163
transform 1 0 20424 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_217
timestamp 1667941163
transform 1 0 21068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_229
timestamp 1667941163
transform 1 0 22172 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_238
timestamp 1667941163
transform 1 0 23000 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1667941163
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_298
timestamp 1667941163
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1667941163
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_12
timestamp 1667941163
transform 1 0 2208 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_24
timestamp 1667941163
transform 1 0 3312 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_36
timestamp 1667941163
transform 1 0 4416 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1667941163
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1667941163
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_62
timestamp 1667941163
transform 1 0 6808 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_76
timestamp 1667941163
transform 1 0 8096 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_80
timestamp 1667941163
transform 1 0 8464 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_84
timestamp 1667941163
transform 1 0 8832 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_97
timestamp 1667941163
transform 1 0 10028 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_101
timestamp 1667941163
transform 1 0 10396 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_124
timestamp 1667941163
transform 1 0 12512 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_132
timestamp 1667941163
transform 1 0 13248 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_144
timestamp 1667941163
transform 1 0 14352 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_153
timestamp 1667941163
transform 1 0 15180 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_165
timestamp 1667941163
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_180
timestamp 1667941163
transform 1 0 17664 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_192
timestamp 1667941163
transform 1 0 18768 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_200
timestamp 1667941163
transform 1 0 19504 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_206
timestamp 1667941163
transform 1 0 20056 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_212
timestamp 1667941163
transform 1 0 20608 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1667941163
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_229
timestamp 1667941163
transform 1 0 22172 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_233
timestamp 1667941163
transform 1 0 22540 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_240
timestamp 1667941163
transform 1 0 23184 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_252
timestamp 1667941163
transform 1 0 24288 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_264
timestamp 1667941163
transform 1 0 25392 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1667941163
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_13
timestamp 1667941163
transform 1 0 2300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_20
timestamp 1667941163
transform 1 0 2944 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_46
timestamp 1667941163
transform 1 0 5336 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_58
timestamp 1667941163
transform 1 0 6440 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_70
timestamp 1667941163
transform 1 0 7544 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1667941163
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_96
timestamp 1667941163
transform 1 0 9936 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_108
timestamp 1667941163
transform 1 0 11040 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_112
timestamp 1667941163
transform 1 0 11408 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_116
timestamp 1667941163
transform 1 0 11776 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_123
timestamp 1667941163
transform 1 0 12420 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_135
timestamp 1667941163
transform 1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_152
timestamp 1667941163
transform 1 0 15088 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_164
timestamp 1667941163
transform 1 0 16192 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_169
timestamp 1667941163
transform 1 0 16652 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_178
timestamp 1667941163
transform 1 0 17480 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1667941163
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_272
timestamp 1667941163
transform 1 0 26128 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_284
timestamp 1667941163
transform 1 0 27232 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_296
timestamp 1667941163
transform 1 0 28336 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_7
timestamp 1667941163
transform 1 0 1748 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_11
timestamp 1667941163
transform 1 0 2116 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_23
timestamp 1667941163
transform 1 0 3220 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_35
timestamp 1667941163
transform 1 0 4324 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_40
timestamp 1667941163
transform 1 0 4784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_44
timestamp 1667941163
transform 1 0 5152 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_67
timestamp 1667941163
transform 1 0 7268 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_74
timestamp 1667941163
transform 1 0 7912 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_86
timestamp 1667941163
transform 1 0 9016 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_101
timestamp 1667941163
transform 1 0 10396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_109
timestamp 1667941163
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_123
timestamp 1667941163
transform 1 0 12420 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_131
timestamp 1667941163
transform 1 0 13156 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_136
timestamp 1667941163
transform 1 0 13616 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_143
timestamp 1667941163
transform 1 0 14260 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_147
timestamp 1667941163
transform 1 0 14628 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_151
timestamp 1667941163
transform 1 0 14996 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_157
timestamp 1667941163
transform 1 0 15548 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1667941163
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_174
timestamp 1667941163
transform 1 0 17112 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_186
timestamp 1667941163
transform 1 0 18216 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_197
timestamp 1667941163
transform 1 0 19228 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_204
timestamp 1667941163
transform 1 0 19872 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_216
timestamp 1667941163
transform 1 0 20976 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_287
timestamp 1667941163
transform 1 0 27508 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_291
timestamp 1667941163
transform 1 0 27876 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_303
timestamp 1667941163
transform 1 0 28980 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_315
timestamp 1667941163
transform 1 0 30084 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_327
timestamp 1667941163
transform 1 0 31188 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_8
timestamp 1667941163
transform 1 0 1840 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_16
timestamp 1667941163
transform 1 0 2576 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_22
timestamp 1667941163
transform 1 0 3128 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_34
timestamp 1667941163
transform 1 0 4232 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_46
timestamp 1667941163
transform 1 0 5336 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_58
timestamp 1667941163
transform 1 0 6440 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_70
timestamp 1667941163
transform 1 0 7544 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1667941163
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_90
timestamp 1667941163
transform 1 0 9384 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_102
timestamp 1667941163
transform 1 0 10488 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_114
timestamp 1667941163
transform 1 0 11592 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_126
timestamp 1667941163
transform 1 0 12696 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_147
timestamp 1667941163
transform 1 0 14628 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_151
timestamp 1667941163
transform 1 0 14996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_158
timestamp 1667941163
transform 1 0 15640 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_242
timestamp 1667941163
transform 1 0 23368 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1667941163
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_7
timestamp 1667941163
transform 1 0 1748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_11
timestamp 1667941163
transform 1 0 2116 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_18
timestamp 1667941163
transform 1 0 2760 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_30
timestamp 1667941163
transform 1 0 3864 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_42
timestamp 1667941163
transform 1 0 4968 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1667941163
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_118
timestamp 1667941163
transform 1 0 11960 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_130
timestamp 1667941163
transform 1 0 13064 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_134
timestamp 1667941163
transform 1 0 13432 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_143
timestamp 1667941163
transform 1 0 14260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_155
timestamp 1667941163
transform 1 0 15364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_178
timestamp 1667941163
transform 1 0 17480 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_190
timestamp 1667941163
transform 1 0 18584 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_202
timestamp 1667941163
transform 1 0 19688 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_214
timestamp 1667941163
transform 1 0 20792 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1667941163
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_244
timestamp 1667941163
transform 1 0 23552 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_256
timestamp 1667941163
transform 1 0 24656 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_268
timestamp 1667941163
transform 1 0 25760 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_401
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_8
timestamp 1667941163
transform 1 0 1840 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_20
timestamp 1667941163
transform 1 0 2944 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_128
timestamp 1667941163
transform 1 0 12880 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_135
timestamp 1667941163
transform 1 0 13524 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_146
timestamp 1667941163
transform 1 0 14536 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_158
timestamp 1667941163
transform 1 0 15640 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_170
timestamp 1667941163
transform 1 0 16744 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_182
timestamp 1667941163
transform 1 0 17848 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1667941163
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_370
timestamp 1667941163
transform 1 0 35144 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_382
timestamp 1667941163
transform 1 0 36248 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_394
timestamp 1667941163
transform 1 0 37352 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1667941163
transform 1 0 38456 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_10
timestamp 1667941163
transform 1 0 2024 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_22
timestamp 1667941163
transform 1 0 3128 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_34
timestamp 1667941163
transform 1 0 4232 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_46
timestamp 1667941163
transform 1 0 5336 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1667941163
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_153
timestamp 1667941163
transform 1 0 15180 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_157
timestamp 1667941163
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_165
timestamp 1667941163
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_398
timestamp 1667941163
transform 1 0 37720 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_406
timestamp 1667941163
transform 1 0 38456 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_353
timestamp 1667941163
transform 1 0 33580 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_365
timestamp 1667941163
transform 1 0 34684 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_377
timestamp 1667941163
transform 1 0 35788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_389
timestamp 1667941163
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_20
timestamp 1667941163
transform 1 0 2944 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_320
timestamp 1667941163
transform 1 0 30544 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_332
timestamp 1667941163
transform 1 0 31648 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_344
timestamp 1667941163
transform 1 0 32752 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_356
timestamp 1667941163
transform 1 0 33856 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_21
timestamp 1667941163
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_33
timestamp 1667941163
transform 1 0 4140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_45
timestamp 1667941163
transform 1 0 5244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1667941163
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_357
timestamp 1667941163
transform 1 0 33948 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_362
timestamp 1667941163
transform 1 0 34408 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_374
timestamp 1667941163
transform 1 0 35512 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_386
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_16
timestamp 1667941163
transform 1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1667941163
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_65
timestamp 1667941163
transform 1 0 7084 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_69
timestamp 1667941163
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1667941163
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_104
timestamp 1667941163
transform 1 0 10672 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_118
timestamp 1667941163
transform 1 0 11960 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_149
timestamp 1667941163
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1667941163
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_174
timestamp 1667941163
transform 1 0 17112 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_182
timestamp 1667941163
transform 1 0 17848 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_203
timestamp 1667941163
transform 1 0 19780 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_211
timestamp 1667941163
transform 1 0 20516 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_217
timestamp 1667941163
transform 1 0 21068 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1667941163
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_233
timestamp 1667941163
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_272
timestamp 1667941163
transform 1 0 26128 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1667941163
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_342
timestamp 1667941163
transform 1 0 32568 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_356
timestamp 1667941163
transform 1 0 33856 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_382
timestamp 1667941163
transform 1 0 36248 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0404_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0405_
timestamp 1667941163
transform 1 0 19596 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0406_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18584 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0407_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0408_
timestamp 1667941163
transform 1 0 4692 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0409_
timestamp 1667941163
transform 1 0 5336 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0410_
timestamp 1667941163
transform 1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0411_
timestamp 1667941163
transform 1 0 23184 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_
timestamp 1667941163
transform 1 0 23184 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0413_
timestamp 1667941163
transform 1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0414_
timestamp 1667941163
transform 1 0 17112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1667941163
transform 1 0 17756 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0416_
timestamp 1667941163
transform 1 0 21988 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 23000 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_
timestamp 1667941163
transform 1 0 22816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 23368 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 22264 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 15732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 17480 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 17204 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform 1 0 18584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 18124 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 9844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 9200 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 10488 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform 1 0 18216 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 18676 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 7636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 6808 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 6164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 11500 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 19596 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 16100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 16836 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 16008 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 19872 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 16468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 26220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1667941163
transform 1 0 15824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 23552 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform 1 0 28336 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 27324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform 1 0 28244 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 29256 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 12972 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 16100 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 3220 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 2576 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform 1 0 1932 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform 1 0 2024 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform 1 0 2668 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 23368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0480_
timestamp 1667941163
transform 1 0 23736 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1667941163
transform 1 0 23368 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 11684 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 6532 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0486_
timestamp 1667941163
transform 1 0 4968 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1667941163
transform 1 0 5060 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0488_
timestamp 1667941163
transform 1 0 13248 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1667941163
transform 1 0 12604 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 20976 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1667941163
transform 1 0 24196 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0493_
timestamp 1667941163
transform 1 0 24564 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1667941163
transform 1 0 21344 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0495_
timestamp 1667941163
transform 1 0 21804 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 20056 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1667941163
transform 1 0 19596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0499_
timestamp 1667941163
transform 1 0 19688 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0500_
timestamp 1667941163
transform 1 0 24472 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0501_
timestamp 1667941163
transform 1 0 24748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 26496 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1667941163
transform 1 0 27784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0505_
timestamp 1667941163
transform 1 0 27140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 20700 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0509_
timestamp 1667941163
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0510_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 21620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 26680 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1667941163
transform 1 0 25668 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0514_
timestamp 1667941163
transform 1 0 25944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0515_
timestamp 1667941163
transform 1 0 21988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform 1 0 21528 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 21344 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1667941163
transform 1 0 23092 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 25024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 25208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0522_
timestamp 1667941163
transform 1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0523_
timestamp 1667941163
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0524_
timestamp 1667941163
transform 1 0 26036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform 1 0 25392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 25668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1667941163
transform 1 0 26312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 2576 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1667941163
transform 1 0 19964 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0532_
timestamp 1667941163
transform 1 0 20056 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0533_
timestamp 1667941163
transform 1 0 15732 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 16376 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform 1 0 18032 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1667941163
transform 1 0 17940 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 27140 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 28980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0540_
timestamp 1667941163
transform 1 0 27048 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0541_
timestamp 1667941163
transform 1 0 26404 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0542_
timestamp 1667941163
transform 1 0 26036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 21252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform 1 0 25208 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1667941163
transform 1 0 24932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 28980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 28244 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 27232 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0550_
timestamp 1667941163
transform 1 0 27692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1667941163
transform 1 0 28336 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1667941163
transform 1 0 28336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 27600 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform 1 0 28244 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 18032 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 13800 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0558_
timestamp 1667941163
transform 1 0 14996 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1667941163
transform 1 0 19320 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 19596 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 20332 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0564_
timestamp 1667941163
transform 1 0 22356 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 10580 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 2668 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform 1 0 8372 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0568_
timestamp 1667941163
transform 1 0 7728 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0569_
timestamp 1667941163
transform 1 0 12144 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1667941163
transform 1 0 13432 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 13156 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 13984 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform 1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 16376 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 3220 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1667941163
transform 1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0577_
timestamp 1667941163
transform 1 0 10120 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1667941163
transform 1 0 16836 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 17204 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform 1 0 14720 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1667941163
transform 1 0 15364 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 17664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1667941163
transform 1 0 7176 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0586_
timestamp 1667941163
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0587_
timestamp 1667941163
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1667941163
transform 1 0 15272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0590_
timestamp 1667941163
transform 1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1667941163
transform 1 0 15456 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1667941163
transform 1 0 27140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0595_
timestamp 1667941163
transform 1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0596_
timestamp 1667941163
transform 1 0 28980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1667941163
transform 1 0 30360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 30452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1667941163
transform 1 0 28980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1667941163
transform 1 0 29808 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 21988 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1667941163
transform 1 0 25484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0604_
timestamp 1667941163
transform 1 0 24932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0605_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1667941163
transform 1 0 22632 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 24380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1667941163
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0609_
timestamp 1667941163
transform 1 0 23368 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 27784 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 27140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1667941163
transform 1 0 26036 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0613_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1667941163
transform 1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 30268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1667941163
transform 1 0 20976 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0622_
timestamp 1667941163
transform 1 0 20976 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0623_
timestamp 1667941163
transform 1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1667941163
transform 1 0 17204 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 3312 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1667941163
transform 1 0 20608 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1667941163
transform 1 0 19688 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 16100 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 18124 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 1667941163
transform 1 0 17848 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0632_
timestamp 1667941163
transform 1 0 15456 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1667941163
transform 1 0 16836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 6624 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1667941163
transform 1 0 16468 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1667941163
transform 1 0 16192 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 23092 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1667941163
transform 1 0 20700 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0640_
timestamp 1667941163
transform 1 0 20792 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0641_
timestamp 1667941163
transform 1 0 25392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 26220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1667941163
transform 1 0 25576 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1667941163
transform 1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 22264 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 22632 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1667941163
transform 1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0649_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1667941163
transform 1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 25208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1667941163
transform 1 0 24748 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 22724 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 23460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform 1 0 25668 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1667941163
transform 1 0 25024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0659_
timestamp 1667941163
transform 1 0 25300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 24656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1667941163
transform 1 0 25208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 10488 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 9200 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1667941163
transform 1 0 12328 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0667_
timestamp 1667941163
transform 1 0 12236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0668_
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 7728 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1667941163
transform 1 0 15640 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1667941163
transform 1 0 14996 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 18032 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 19320 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0675_
timestamp 1667941163
transform 1 0 16928 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0676_
timestamp 1667941163
transform 1 0 17112 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 4232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1667941163
transform 1 0 19320 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0679_
timestamp 1667941163
transform 1 0 20516 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1667941163
transform 1 0 19504 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1667941163
transform 1 0 20148 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 22632 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0685_
timestamp 1667941163
transform 1 0 22356 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0686_
timestamp 1667941163
transform 1 0 23092 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1667941163
transform 1 0 28336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1667941163
transform 1 0 27784 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 27416 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 30360 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 28980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 5152 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 18676 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 4692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 27508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 33304 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 27600 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 33304 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 5336 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0706_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 33396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 9660 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0710_
timestamp 1667941163
transform 1 0 32752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 1840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 32108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 21252 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 30084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 17296 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 31004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0718_
timestamp 1667941163
transform 1 0 32200 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0719_
timestamp 1667941163
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 1932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 19596 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0725_
timestamp 1667941163
transform 1 0 3956 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 14260 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 31464 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 31648 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 31188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 28796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 28244 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 20792 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 1840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 13248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 31004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 29440 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 17572 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 26496 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 27508 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 31280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 1840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 22724 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 33488 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 15272 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 9108 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0751_
timestamp 1667941163
transform 1 0 4416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0752_
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 25668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 29716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 1840 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0756_
timestamp 1667941163
transform 1 0 1840 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 25024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 32292 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 29808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 28704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 4784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 18584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 4784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 14076 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 7636 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 18308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 14720 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 3956 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 19780 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 23736 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 26312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 3956 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 26128 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0783_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10120 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0784_
timestamp 1667941163
transform 1 0 15732 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 13156 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 12236 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 13340 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 16100 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 16008 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 15456 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 16928 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 12880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0795_
timestamp 1667941163
transform 1 0 15824 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 13524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 14444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 16376 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 14720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 15640 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 15272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0806_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16376 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 6624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 7544 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 14996 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 7452 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 7728 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 9568 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0817_
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 15732 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 15364 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 14536 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 15272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 14996 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 14628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0828_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 9200 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 16376 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 12788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 17480 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 15088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 8188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 8372 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 11592 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 15732 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0839_
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 14720 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 15824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 13800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 15364 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0850_
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1667941163
transform 1 0 4324 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 9568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 3220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 5336 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 3128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1667941163
transform 1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1667941163
transform 1 0 4968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 13064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0865_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0866_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5888 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0867_
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0868_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10948 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0869_
timestamp 1667941163
transform 1 0 9108 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0870_
timestamp 1667941163
transform 1 0 9384 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0871_
timestamp 1667941163
transform 1 0 14168 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0872_
timestamp 1667941163
transform 1 0 10304 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0873_
timestamp 1667941163
transform 1 0 13432 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0874_
timestamp 1667941163
transform 1 0 10948 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0875_
timestamp 1667941163
transform 1 0 9476 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0876_
timestamp 1667941163
transform 1 0 14260 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0878_
timestamp 1667941163
transform 1 0 10488 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0879_
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0880_
timestamp 1667941163
transform 1 0 8004 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0881_
timestamp 1667941163
transform 1 0 2576 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0882_
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0883_
timestamp 1667941163
transform 1 0 9384 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0884_
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0885_
timestamp 1667941163
transform -1 0 13616 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0886_
timestamp 1667941163
transform 1 0 5428 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0887_
timestamp 1667941163
transform 1 0 3956 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0888_
timestamp 1667941163
transform 1 0 11684 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0889_
timestamp 1667941163
transform 1 0 6532 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0890_
timestamp 1667941163
transform 1 0 1840 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0891_
timestamp 1667941163
transform 1 0 1748 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0892_
timestamp 1667941163
transform 1 0 6532 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0893_
timestamp 1667941163
transform 1 0 10304 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0894_
timestamp 1667941163
transform 1 0 13156 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0895_
timestamp 1667941163
transform 1 0 3956 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0896_
timestamp 1667941163
transform 1 0 8832 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0897_
timestamp 1667941163
transform 1 0 12972 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0898_
timestamp 1667941163
transform 1 0 11500 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0899_
timestamp 1667941163
transform 1 0 2208 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0900_
timestamp 1667941163
transform 1 0 7268 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0901_
timestamp 1667941163
transform 1 0 12880 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0902_
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0903_
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0904_
timestamp 1667941163
transform 1 0 13064 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0905_
timestamp 1667941163
transform 1 0 6072 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0906_
timestamp 1667941163
transform 1 0 4324 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0907_
timestamp 1667941163
transform 1 0 12880 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 10304 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0909_
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0910_
timestamp 1667941163
transform 1 0 12880 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0911_
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 1932 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0913_
timestamp 1667941163
transform 1 0 6900 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0914_
timestamp 1667941163
transform 1 0 13248 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0915_
timestamp 1667941163
transform 1 0 3956 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0916_
timestamp 1667941163
transform 1 0 1564 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0917_
timestamp 1667941163
transform 1 0 3864 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0918_
timestamp 1667941163
transform 1 0 4416 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0919_
timestamp 1667941163
transform 1 0 8924 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0920_
timestamp 1667941163
transform 1 0 4968 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0921_
timestamp 1667941163
transform 1 0 13800 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 8096 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0923_
timestamp 1667941163
transform 1 0 9844 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 1564 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0925_
timestamp 1667941163
transform 1 0 9752 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0926_
timestamp 1667941163
transform 1 0 6808 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0927_
timestamp 1667941163
transform 1 0 3956 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 4324 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0929_
timestamp 1667941163
transform 1 0 2300 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0930_
timestamp 1667941163
transform 1 0 7360 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0931_
timestamp 1667941163
transform 1 0 5888 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0932_
timestamp 1667941163
transform 1 0 6992 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0933_
timestamp 1667941163
transform 1 0 6532 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0934_
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 13248 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0936_
timestamp 1667941163
transform 1 0 9108 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0937_
timestamp 1667941163
transform 1 0 9108 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform 1 0 10212 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _0976_
timestamp 1667941163
transform 1 0 32292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1667941163
transform 1 0 31464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0978_
timestamp 1667941163
transform 1 0 32936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 1667941163
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1667941163
transform 1 0 1748 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0981_
timestamp 1667941163
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0982_
timestamp 1667941163
transform 1 0 17204 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1667941163
transform 1 0 23276 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1667941163
transform 1 0 31188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1667941163
transform 1 0 1748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1667941163
transform 1 0 32292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1667941163
transform 1 0 13800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1667941163
transform 1 0 34132 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1667941163
transform 1 0 34132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1667941163
transform 1 0 32292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1667941163
transform 1 0 11500 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 20792 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 37444 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1667941163
transform 1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1667941163
transform 1 0 2852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 18952 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1667941163
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1667941163
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1667941163
transform 1 0 4140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 1748 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 30912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 32936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 34868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 23092 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 30268 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 4784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1014_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27140 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1015_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1015__100 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1016_
timestamp 1667941163
transform 1 0 23276 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1017_
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1018_
timestamp 1667941163
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1019_
timestamp 1667941163
transform 1 0 29532 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1020_
timestamp 1667941163
transform 1 0 19412 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1021_
timestamp 1667941163
transform 1 0 18032 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1021__101
timestamp 1667941163
transform 1 0 18216 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1022_
timestamp 1667941163
transform 1 0 16836 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1023_
timestamp 1667941163
transform 1 0 18768 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1024_
timestamp 1667941163
transform 1 0 3956 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1025_
timestamp 1667941163
transform 1 0 19596 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1026_
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1027__102
timestamp 1667941163
transform 1 0 11684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1027_
timestamp 1667941163
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1028_
timestamp 1667941163
transform 1 0 11316 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1029_
timestamp 1667941163
transform 1 0 10396 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1030_
timestamp 1667941163
transform 1 0 8372 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1031_
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1032_
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1033_
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1033__103
timestamp 1667941163
transform 1 0 25116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1034_
timestamp 1667941163
transform 1 0 22172 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1035_
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1036_
timestamp 1667941163
transform 1 0 24656 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1037_
timestamp 1667941163
transform 1 0 23092 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1038_
timestamp 1667941163
transform 1 0 24564 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1039__104
timestamp 1667941163
transform 1 0 23368 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1039_
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1040_
timestamp 1667941163
transform 1 0 21252 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1041_
timestamp 1667941163
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1042_
timestamp 1667941163
transform 1 0 25024 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1043_
timestamp 1667941163
transform 1 0 22540 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1044_
timestamp 1667941163
transform 1 0 25576 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1045__105
timestamp 1667941163
transform 1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1045_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1046_
timestamp 1667941163
transform 1 0 20608 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1047_
timestamp 1667941163
transform 1 0 21896 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1048_
timestamp 1667941163
transform 1 0 24748 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1049_
timestamp 1667941163
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1050_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17572 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1051__106
timestamp 1667941163
transform 1 0 17296 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 17204 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1052_
timestamp 1667941163
transform 1 0 17940 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1053_
timestamp 1667941163
transform 1 0 17756 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1054_
timestamp 1667941163
transform 1 0 9108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1055_
timestamp 1667941163
transform 1 0 18584 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1056_
timestamp 1667941163
transform 1 0 17296 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1057_
timestamp 1667941163
transform 1 0 19136 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1057__107
timestamp 1667941163
transform 1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1058_
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1059_
timestamp 1667941163
transform 1 0 18768 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1060_
timestamp 1667941163
transform 1 0 3956 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1061_
timestamp 1667941163
transform 1 0 19780 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1062_
timestamp 1667941163
transform 1 0 30452 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1063_
timestamp 1667941163
transform 1 0 29716 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1063__108
timestamp 1667941163
transform 1 0 29624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1064_
timestamp 1667941163
transform 1 0 26680 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1065_
timestamp 1667941163
transform 1 0 28428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1066_
timestamp 1667941163
transform 1 0 29900 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1067_
timestamp 1667941163
transform 1 0 27140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1068_
timestamp 1667941163
transform 1 0 19688 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1069__109
timestamp 1667941163
transform 1 0 22632 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1069_
timestamp 1667941163
transform 1 0 23184 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1070_
timestamp 1667941163
transform 1 0 22540 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1071_
timestamp 1667941163
transform 1 0 20240 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1072_
timestamp 1667941163
transform 1 0 24840 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1073_
timestamp 1667941163
transform 1 0 22448 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1074_
timestamp 1667941163
transform 1 0 30452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1075__110
timestamp 1667941163
transform 1 0 30912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1075_
timestamp 1667941163
transform 1 0 30360 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 26128 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1077_
timestamp 1667941163
transform 1 0 26404 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1078_
timestamp 1667941163
transform 1 0 32292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1079_
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1080_
timestamp 1667941163
transform 1 0 17112 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1081__111
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1081_
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1082_
timestamp 1667941163
transform 1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1083_
timestamp 1667941163
transform 1 0 11684 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1084_
timestamp 1667941163
transform 1 0 17020 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1085_
timestamp 1667941163
transform 1 0 18124 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1086_
timestamp 1667941163
transform 1 0 16836 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1087__112
timestamp 1667941163
transform 1 0 16008 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1087_
timestamp 1667941163
transform 1 0 15640 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1088_
timestamp 1667941163
transform 1 0 9200 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1089_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1090_
timestamp 1667941163
transform 1 0 12788 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1091_
timestamp 1667941163
transform 1 0 4140 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1092_
timestamp 1667941163
transform 1 0 14352 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1093_
timestamp 1667941163
transform 1 0 15548 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1093__113
timestamp 1667941163
transform 1 0 14904 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1094_
timestamp 1667941163
transform 1 0 7360 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1095_
timestamp 1667941163
transform 1 0 11224 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1096_
timestamp 1667941163
transform 1 0 12972 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1097_
timestamp 1667941163
transform 1 0 3312 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1098_
timestamp 1667941163
transform 1 0 19136 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1099_
timestamp 1667941163
transform 1 0 20608 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1099__114
timestamp 1667941163
transform 1 0 20608 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1100_
timestamp 1667941163
transform 1 0 14536 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1101_
timestamp 1667941163
transform 1 0 17480 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1102_
timestamp 1667941163
transform 1 0 18216 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1103_
timestamp 1667941163
transform 1 0 13156 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1104_
timestamp 1667941163
transform 1 0 29716 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1105__115
timestamp 1667941163
transform 1 0 28428 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1105_
timestamp 1667941163
transform 1 0 27324 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1106_
timestamp 1667941163
transform 1 0 27876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1107_
timestamp 1667941163
transform 1 0 30084 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1108_
timestamp 1667941163
transform 1 0 28520 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1109_
timestamp 1667941163
transform 1 0 28888 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1110_
timestamp 1667941163
transform 1 0 24656 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1111__116
timestamp 1667941163
transform 1 0 23276 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1111_
timestamp 1667941163
transform 1 0 23276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1112_
timestamp 1667941163
transform 1 0 27140 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1113_
timestamp 1667941163
transform 1 0 27140 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1114_
timestamp 1667941163
transform 1 0 22172 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 27876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1116_
timestamp 1667941163
transform 1 0 15916 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1117_
timestamp 1667941163
transform 1 0 16928 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1117__117
timestamp 1667941163
transform 1 0 17204 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1118_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1119_
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1120_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1121_
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1122_
timestamp 1667941163
transform 1 0 24104 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1123__118
timestamp 1667941163
transform 1 0 22632 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1123_
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1124_
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1125_
timestamp 1667941163
transform 1 0 25300 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1126_
timestamp 1667941163
transform 1 0 23736 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1127_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1128_
timestamp 1667941163
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1129__119
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1129_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1130_
timestamp 1667941163
transform 1 0 25392 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1131_
timestamp 1667941163
transform 1 0 20424 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1132_
timestamp 1667941163
transform 1 0 20148 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1133_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1134_
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1135__120
timestamp 1667941163
transform 1 0 18952 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1135_
timestamp 1667941163
transform 1 0 19596 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1136_
timestamp 1667941163
transform 1 0 25760 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1137_
timestamp 1667941163
transform 1 0 17664 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1138_
timestamp 1667941163
transform 1 0 20056 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1139_
timestamp 1667941163
transform 1 0 25852 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1140_
timestamp 1667941163
transform 1 0 23276 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1140__121
timestamp 1667941163
transform 1 0 23368 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1141_
timestamp 1667941163
transform 1 0 20148 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1142_
timestamp 1667941163
transform 1 0 19688 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1143_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1144__122
timestamp 1667941163
transform 1 0 21160 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1144_
timestamp 1667941163
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1145_
timestamp 1667941163
transform 1 0 20516 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1146_
timestamp 1667941163
transform 1 0 21896 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1147_
timestamp 1667941163
transform 1 0 20608 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1148__123
timestamp 1667941163
transform 1 0 14260 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1148_
timestamp 1667941163
transform 1 0 13524 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1149_
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1150_
timestamp 1667941163
transform 1 0 11684 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1151_
timestamp 1667941163
transform 1 0 6532 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1152_
timestamp 1667941163
transform 1 0 14352 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1152__124
timestamp 1667941163
transform 1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1153_
timestamp 1667941163
transform 1 0 22632 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1154_
timestamp 1667941163
transform 1 0 15548 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1155_
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1156__125
timestamp 1667941163
transform 1 0 4416 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 2668 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1157_
timestamp 1667941163
transform 1 0 1840 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1158_
timestamp 1667941163
transform 1 0 2944 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1159_
timestamp 1667941163
transform 1 0 1840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1160__126
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1160_
timestamp 1667941163
transform 1 0 11684 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1161_
timestamp 1667941163
transform 1 0 19044 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1162_
timestamp 1667941163
transform 1 0 14260 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1163_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1164__127
timestamp 1667941163
transform 1 0 28336 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1164_
timestamp 1667941163
transform 1 0 28244 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1165_
timestamp 1667941163
transform 1 0 27968 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 28152 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1167_
timestamp 1667941163
transform 1 0 28336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1168__128
timestamp 1667941163
transform 1 0 22724 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 23092 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1169_
timestamp 1667941163
transform 1 0 11684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1170_
timestamp 1667941163
transform 1 0 21896 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1171_
timestamp 1667941163
transform 1 0 20608 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1172__129
timestamp 1667941163
transform 1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1172_
timestamp 1667941163
transform 1 0 16192 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1173_
timestamp 1667941163
transform 1 0 21712 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1174_
timestamp 1667941163
transform 1 0 17756 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 17480 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1176_
timestamp 1667941163
transform 1 0 18492 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1176__130
timestamp 1667941163
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1177_
timestamp 1667941163
transform 1 0 15732 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1178_
timestamp 1667941163
transform 1 0 19136 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1179_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1180__131
timestamp 1667941163
transform 1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1180_
timestamp 1667941163
transform 1 0 9108 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1181_
timestamp 1667941163
transform 1 0 6440 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 2668 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1183_
timestamp 1667941163
transform 1 0 6808 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1184__132
timestamp 1667941163
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 18768 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1185_
timestamp 1667941163
transform 1 0 12420 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 18124 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1187_
timestamp 1667941163
transform 1 0 11776 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1188_
timestamp 1667941163
transform 1 0 17204 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1188__133
timestamp 1667941163
transform 1 0 17296 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1189_
timestamp 1667941163
transform 1 0 17020 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1190_
timestamp 1667941163
transform 1 0 17020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 18492 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1192_
timestamp 1667941163
transform 1 0 20700 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1192__134
timestamp 1667941163
transform 1 0 20700 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform 1 0 23644 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1194_
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1195_
timestamp 1667941163
transform 1 0 23368 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1196__135
timestamp 1667941163
transform 1 0 17020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1197_
timestamp 1667941163
transform 1 0 22080 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1198_
timestamp 1667941163
transform 1 0 17664 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1199_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1200_
timestamp 1667941163
transform 1 0 5704 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1200__136
timestamp 1667941163
transform 1 0 6532 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1201_
timestamp 1667941163
transform 1 0 19136 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 17296 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1203_
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 38088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 38088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 38088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 2944 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 36708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 38088 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 14904 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 38088 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform 1 0 1564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 38088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 38088 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 1564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 5244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 38088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 1564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 31004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 38088 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 38088 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 2300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 38088 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 20700 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 12972 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 1564 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 18584 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 1564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 36616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 35880 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 7820 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 0 nsew signal input
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 1 nsew signal input
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 2 nsew signal input
flabel metal3 s 39200 11568 39800 11688 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 3 nsew signal input
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 4 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 5 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 6 nsew signal input
flabel metal2 s 15474 200 15530 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 7 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 8 nsew signal input
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 9 nsew signal input
flabel metal3 s 39200 31288 39800 31408 0 FreeSans 480 0 0 0 ccff_head
port 10 nsew signal input
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 ccff_tail
port 11 nsew signal tristate
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_right_in[0]
port 12 nsew signal input
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 13 nsew signal input
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chanx_right_in[11]
port 14 nsew signal input
flabel metal3 s 39200 19728 39800 19848 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 15 nsew signal input
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chanx_right_in[13]
port 16 nsew signal input
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 17 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 18 nsew signal input
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 chanx_right_in[16]
port 19 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 20 nsew signal input
flabel metal3 s 39200 34688 39800 34808 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 21 nsew signal input
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 22 nsew signal input
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chanx_right_in[2]
port 23 nsew signal input
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 24 nsew signal input
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_right_in[4]
port 25 nsew signal input
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_right_in[5]
port 26 nsew signal input
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 27 nsew signal input
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 28 nsew signal input
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 29 nsew signal input
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 30 nsew signal input
flabel metal3 s 39200 36728 39800 36848 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 31 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 32 nsew signal tristate
flabel metal2 s 23846 39200 23902 39800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 33 nsew signal tristate
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_right_out[12]
port 34 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 35 nsew signal tristate
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 36 nsew signal tristate
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 37 nsew signal tristate
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 38 nsew signal tristate
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chanx_right_out[17]
port 39 nsew signal tristate
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 40 nsew signal tristate
flabel metal2 s 20626 39200 20682 39800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 41 nsew signal tristate
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 42 nsew signal tristate
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 43 nsew signal tristate
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 44 nsew signal tristate
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 45 nsew signal tristate
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 46 nsew signal tristate
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 47 nsew signal tristate
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 48 nsew signal tristate
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 49 nsew signal tristate
flabel metal3 s 200 2728 800 2848 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 50 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chany_bottom_in[10]
port 51 nsew signal input
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 52 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 53 nsew signal input
flabel metal2 s 34794 39200 34850 39800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 54 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 55 nsew signal input
flabel metal2 s 2594 200 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 56 nsew signal input
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 57 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 58 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[18]
port 59 nsew signal input
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 60 nsew signal input
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 61 nsew signal input
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 62 nsew signal input
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 63 nsew signal input
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 64 nsew signal input
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 65 nsew signal input
flabel metal3 s 200 16328 800 16448 0 FreeSans 480 0 0 0 chany_bottom_in[7]
port 66 nsew signal input
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 67 nsew signal input
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 chany_bottom_in[9]
port 68 nsew signal input
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 69 nsew signal tristate
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 70 nsew signal tristate
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 71 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 72 nsew signal tristate
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 73 nsew signal tristate
flabel metal3 s 200 8168 800 8288 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 74 nsew signal tristate
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 75 nsew signal tristate
flabel metal3 s 200 12928 800 13048 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 76 nsew signal tristate
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 77 nsew signal tristate
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 78 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal2 s 7746 200 7802 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal2 s 12254 200 12310 800 0 FreeSans 224 90 0 0 pReset
port 88 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 prog_clk
port 89 nsew signal input
flabel metal3 s 39200 23128 39800 23248 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 90 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 91 nsew signal input
flabel metal2 s 31574 39200 31630 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 92 nsew signal input
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 93 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 94 nsew signal input
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 95 nsew signal input
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
port 96 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
port 97 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
port 98 nsew signal input
flabel metal3 s 39200 18368 39800 18488 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
port 99 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 16100 24718 16100 24718 0 _0000_
rlabel metal1 14628 24038 14628 24038 0 _0001_
rlabel metal1 15594 22950 15594 22950 0 _0002_
rlabel metal2 13478 20638 13478 20638 0 _0003_
rlabel metal2 14950 18088 14950 18088 0 _0004_
rlabel metal2 15410 16320 15410 16320 0 _0005_
rlabel metal1 15180 13158 15180 13158 0 _0006_
rlabel metal1 14681 12886 14681 12886 0 _0007_
rlabel metal1 8471 12138 8471 12138 0 _0008_
rlabel metal1 6033 17578 6033 17578 0 _0009_
rlabel metal1 14352 15674 14352 15674 0 _0010_
rlabel metal1 12381 16490 12381 16490 0 _0011_
rlabel metal1 16284 27370 16284 27370 0 _0012_
rlabel metal2 15226 20230 15226 20230 0 _0013_
rlabel metal1 3871 21930 3871 21930 0 _0014_
rlabel metal1 6992 25126 6992 25126 0 _0015_
rlabel metal1 11362 14518 11362 14518 0 _0016_
rlabel metal2 15870 17374 15870 17374 0 _0017_
rlabel metal1 8379 23018 8379 23018 0 _0018_
rlabel metal1 3135 9962 3135 9962 0 _0019_
rlabel metal2 6026 9180 6026 9180 0 _0020_
rlabel metal2 13938 20672 13938 20672 0 _0021_
rlabel metal2 11362 15368 11362 15368 0 _0022_
rlabel via2 16606 5627 16606 5627 0 _0023_
rlabel metal1 14299 10710 14299 10710 0 _0024_
rlabel metal2 15318 10302 15318 10302 0 _0025_
rlabel metal1 14168 6358 14168 6358 0 _0026_
rlabel metal2 3818 8806 3818 8806 0 _0027_
rlabel metal1 7498 15130 7498 15130 0 _0028_
rlabel metal1 9384 8058 9384 8058 0 _0029_
rlabel metal1 4048 14586 4048 14586 0 _0030_
rlabel metal2 4094 16966 4094 16966 0 _0031_
rlabel metal1 4002 10234 4002 10234 0 _0032_
rlabel metal1 7038 8058 7038 8058 0 _0033_
rlabel metal1 5888 16422 5888 16422 0 _0034_
rlabel metal2 7590 9792 7590 9792 0 _0035_
rlabel metal1 4508 14518 4508 14518 0 _0036_
rlabel metal2 3266 12648 3266 12648 0 _0037_
rlabel metal1 14674 8425 14674 8425 0 _0038_
rlabel metal2 5106 16388 5106 16388 0 _0039_
rlabel metal2 13202 8704 13202 8704 0 _0040_
rlabel metal2 13018 9282 13018 9282 0 _0041_
rlabel metal1 14168 26010 14168 26010 0 _0042_
rlabel metal1 10396 24718 10396 24718 0 _0043_
rlabel metal2 13110 29189 13110 29189 0 _0044_
rlabel metal1 12696 32198 12696 32198 0 _0045_
rlabel metal2 14858 25976 14858 25976 0 _0046_
rlabel metal2 13846 28934 13846 28934 0 _0047_
rlabel metal2 14950 10846 14950 10846 0 _0048_
rlabel metal1 13846 18700 13846 18700 0 _0049_
rlabel metal1 16560 25670 16560 25670 0 _0050_
rlabel metal1 12926 13498 12926 13498 0 _0051_
rlabel metal1 11093 19754 11093 19754 0 _0052_
rlabel metal2 14582 21794 14582 21794 0 _0053_
rlabel metal1 11461 24106 11461 24106 0 _0054_
rlabel metal1 13478 21964 13478 21964 0 _0055_
rlabel metal1 6355 14382 6355 14382 0 _0056_
rlabel metal2 10994 26214 10994 26214 0 _0057_
rlabel metal1 9936 11322 9936 11322 0 _0058_
rlabel metal2 16238 12138 16238 12138 0 _0059_
rlabel metal1 14950 11798 14950 11798 0 _0060_
rlabel metal1 15923 15062 15923 15062 0 _0061_
rlabel metal1 9016 8534 9016 8534 0 _0062_
rlabel metal1 6348 5882 6348 5882 0 _0063_
rlabel metal2 6762 10472 6762 10472 0 _0064_
rlabel metal1 9890 5610 9890 5610 0 _0065_
rlabel metal1 7636 22406 7636 22406 0 _0066_
rlabel metal2 15134 12580 15134 12580 0 _0067_
rlabel metal1 5389 24786 5389 24786 0 _0068_
rlabel metal2 7866 22712 7866 22712 0 _0069_
rlabel metal2 9706 21352 9706 21352 0 _0070_
rlabel metal1 13478 19448 13478 19448 0 _0071_
rlabel metal1 14812 24378 14812 24378 0 _0072_
rlabel metal1 12933 22678 12933 22678 0 _0073_
rlabel metal1 19044 10234 19044 10234 0 _0074_
rlabel metal1 5474 28050 5474 28050 0 _0075_
rlabel metal1 23138 20026 23138 20026 0 _0076_
rlabel metal1 17572 9146 17572 9146 0 _0077_
rlabel metal2 23598 27642 23598 27642 0 _0078_
rlabel metal1 23138 31348 23138 31348 0 _0079_
rlabel metal1 17112 18258 17112 18258 0 _0080_
rlabel metal2 17710 10982 17710 10982 0 _0081_
rlabel metal1 9982 30906 9982 30906 0 _0082_
rlabel metal1 18584 12410 18584 12410 0 _0083_
rlabel metal2 6394 29818 6394 29818 0 _0084_
rlabel metal1 13294 5610 13294 5610 0 _0085_
rlabel metal2 16882 28934 16882 28934 0 _0086_
rlabel metal1 20056 15130 20056 15130 0 _0087_
rlabel metal1 19642 8432 19642 8432 0 _0088_
rlabel metal1 18354 7956 18354 7956 0 _0089_
rlabel metal1 27876 25262 27876 25262 0 _0090_
rlabel metal1 12696 5678 12696 5678 0 _0091_
rlabel metal1 23782 8432 23782 8432 0 _0092_
rlabel metal2 28474 14076 28474 14076 0 _0093_
rlabel metal1 29624 20570 29624 20570 0 _0094_
rlabel metal1 20562 6324 20562 6324 0 _0095_
rlabel metal2 12098 5338 12098 5338 0 _0096_
rlabel metal2 1978 31110 1978 31110 0 _0097_
rlabel metal1 2898 31824 2898 31824 0 _0098_
rlabel metal2 23782 6460 23782 6460 0 _0099_
rlabel metal2 15686 6596 15686 6596 0 _0100_
rlabel metal1 5152 31450 5152 31450 0 _0101_
rlabel metal1 13064 33966 13064 33966 0 _0102_
rlabel metal2 24242 21828 24242 21828 0 _0103_
rlabel metal1 21712 27642 21712 27642 0 _0104_
rlabel metal1 19826 22746 19826 22746 0 _0105_
rlabel metal2 24978 13668 24978 13668 0 _0106_
rlabel metal1 27600 9554 27600 9554 0 _0107_
rlabel metal2 16882 3638 16882 3638 0 _0108_
rlabel metal1 22448 7378 22448 7378 0 _0109_
rlabel metal2 26174 11594 26174 11594 0 _0110_
rlabel metal1 21896 12410 21896 12410 0 _0111_
rlabel metal1 23690 10030 23690 10030 0 _0112_
rlabel metal1 21804 14382 21804 14382 0 _0113_
rlabel metal1 25852 18734 25852 18734 0 _0114_
rlabel metal1 25967 19958 25967 19958 0 _0115_
rlabel metal1 20148 25466 20148 25466 0 _0116_
rlabel metal1 16606 15504 16606 15504 0 _0117_
rlabel metal2 18170 13770 18170 13770 0 _0118_
rlabel metal2 27094 25670 27094 25670 0 _0119_
rlabel metal2 26082 22406 26082 22406 0 _0120_
rlabel metal2 25162 23868 25162 23868 0 _0121_
rlabel metal2 27922 20604 27922 20604 0 _0122_
rlabel metal2 28382 24310 28382 24310 0 _0123_
rlabel metal1 28474 24208 28474 24208 0 _0124_
rlabel metal2 15042 28492 15042 28492 0 _0125_
rlabel metal1 19596 20910 19596 20910 0 _0126_
rlabel metal2 22586 19516 22586 19516 0 _0127_
rlabel metal1 8188 30702 8188 30702 0 _0128_
rlabel metal1 12926 31926 12926 31926 0 _0129_
rlabel metal1 14536 31790 14536 31790 0 _0130_
rlabel metal1 10626 32402 10626 32402 0 _0131_
rlabel metal2 17434 31994 17434 31994 0 _0132_
rlabel metal1 15594 32912 15594 32912 0 _0133_
rlabel metal2 7222 6460 7222 6460 0 _0134_
rlabel metal1 14306 7378 14306 7378 0 _0135_
rlabel metal1 15686 20944 15686 20944 0 _0136_
rlabel metal1 26151 16558 26151 16558 0 _0137_
rlabel metal1 29808 15130 29808 15130 0 _0138_
rlabel metal1 29532 17170 29532 17170 0 _0139_
rlabel metal2 25530 16388 25530 16388 0 _0140_
rlabel metal2 22862 14586 22862 14586 0 _0141_
rlabel metal2 23598 11594 23598 11594 0 _0142_
rlabel metal1 27370 13974 27370 13974 0 _0143_
rlabel metal1 29026 13260 29026 13260 0 _0144_
rlabel metal2 29946 17850 29946 17850 0 _0145_
rlabel metal2 21022 16388 21022 16388 0 _0146_
rlabel metal1 17664 15470 17664 15470 0 _0147_
rlabel metal1 20286 24786 20286 24786 0 _0148_
rlabel metal2 18078 23868 18078 23868 0 _0149_
rlabel metal2 17066 27676 17066 27676 0 _0150_
rlabel metal2 16514 26962 16514 26962 0 _0151_
rlabel metal2 21022 24956 21022 24956 0 _0152_
rlabel metal1 25829 22950 25829 22950 0 _0153_
rlabel metal2 25622 14756 25622 14756 0 _0154_
rlabel metal2 21942 20230 21942 20230 0 _0155_
rlabel metal2 24610 26894 24610 26894 0 _0156_
rlabel metal2 24978 28730 24978 28730 0 _0157_
rlabel metal1 25484 12818 25484 12818 0 _0158_
rlabel metal2 25346 9996 25346 9996 0 _0159_
rlabel metal2 25254 8636 25254 8636 0 _0160_
rlabel metal2 12374 29750 12374 29750 0 _0161_
rlabel metal1 8694 29138 8694 29138 0 _0162_
rlabel metal1 15226 18768 15226 18768 0 _0163_
rlabel metal2 17342 30090 17342 30090 0 _0164_
rlabel metal1 20056 27098 20056 27098 0 _0165_
rlabel metal1 20378 30668 20378 30668 0 _0166_
rlabel metal2 22402 25670 22402 25670 0 _0167_
rlabel metal1 28198 15130 28198 15130 0 _0168_
rlabel metal1 11684 5270 11684 5270 0 _0169_
rlabel metal1 13524 12206 13524 12206 0 _0170_
rlabel metal1 16146 11764 16146 11764 0 _0171_
rlabel metal2 6854 8704 6854 8704 0 _0172_
rlabel metal1 14858 11730 14858 11730 0 _0173_
rlabel metal1 15134 19788 15134 19788 0 _0174_
rlabel metal2 16882 6289 16882 6289 0 _0175_
rlabel metal2 5382 8398 5382 8398 0 _0176_
rlabel metal1 27554 23766 27554 23766 0 _0177_
rlabel metal1 28198 15674 28198 15674 0 _0178_
rlabel metal2 23506 25228 23506 25228 0 _0179_
rlabel metal2 25346 24990 25346 24990 0 _0180_
rlabel metal1 23184 24650 23184 24650 0 _0181_
rlabel metal2 29854 15844 29854 15844 0 _0182_
rlabel metal1 19918 29682 19918 29682 0 _0183_
rlabel metal2 20562 27846 20562 27846 0 _0184_
rlabel metal1 17112 28050 17112 28050 0 _0185_
rlabel metal2 18998 29580 18998 29580 0 _0186_
rlabel metal2 4370 27234 4370 27234 0 _0187_
rlabel metal2 19458 28322 19458 28322 0 _0188_
rlabel metal1 6808 23766 6808 23766 0 _0189_
rlabel metal1 14214 18870 14214 18870 0 _0190_
rlabel metal2 11546 29852 11546 29852 0 _0191_
rlabel metal2 10626 28968 10626 28968 0 _0192_
rlabel metal2 7866 6120 7866 6120 0 _0193_
rlabel metal2 9338 29852 9338 29852 0 _0194_
rlabel metal1 24702 9486 24702 9486 0 _0195_
rlabel metal1 25806 8364 25806 8364 0 _0196_
rlabel metal1 24472 12682 24472 12682 0 _0197_
rlabel metal1 23000 10642 23000 10642 0 _0198_
rlabel metal2 24886 10268 24886 10268 0 _0199_
rlabel metal1 23460 20434 23460 20434 0 _0200_
rlabel metal2 24794 27166 24794 27166 0 _0201_
rlabel metal1 24518 28730 24518 28730 0 _0202_
rlabel metal1 21758 20570 21758 20570 0 _0203_
rlabel metal1 23506 21896 23506 21896 0 _0204_
rlabel metal1 25300 27642 25300 27642 0 _0205_
rlabel metal2 22770 15844 22770 15844 0 _0206_
rlabel metal2 26634 23528 26634 23528 0 _0207_
rlabel metal2 25898 15300 25898 15300 0 _0208_
rlabel metal2 20838 24412 20838 24412 0 _0209_
rlabel metal2 22126 23970 22126 23970 0 _0210_
rlabel metal2 26358 14756 26358 14756 0 _0211_
rlabel metal2 22310 23834 22310 23834 0 _0212_
rlabel metal1 17342 25942 17342 25942 0 _0213_
rlabel metal1 16836 26282 16836 26282 0 _0214_
rlabel metal1 18032 22066 18032 22066 0 _0215_
rlabel metal1 17986 20808 17986 20808 0 _0216_
rlabel metal1 8786 28458 8786 28458 0 _0217_
rlabel metal1 18538 23290 18538 23290 0 _0218_
rlabel metal2 17250 15912 17250 15912 0 _0219_
rlabel metal1 19550 24922 19550 24922 0 _0220_
rlabel metal2 21022 16932 21022 16932 0 _0221_
rlabel metal1 18722 16762 18722 16762 0 _0222_
rlabel metal1 4186 25160 4186 25160 0 _0223_
rlabel metal1 20516 18190 20516 18190 0 _0224_
rlabel metal1 30682 13260 30682 13260 0 _0225_
rlabel metal1 29808 17850 29808 17850 0 _0226_
rlabel metal1 27048 13362 27048 13362 0 _0227_
rlabel metal1 28290 12818 28290 12818 0 _0228_
rlabel metal2 30406 20196 30406 20196 0 _0229_
rlabel metal1 27324 11730 27324 11730 0 _0230_
rlabel metal1 19918 14280 19918 14280 0 _0231_
rlabel metal2 23414 11492 23414 11492 0 _0232_
rlabel metal1 23782 17034 23782 17034 0 _0233_
rlabel metal1 20838 17306 20838 17306 0 _0234_
rlabel metal1 25024 11186 25024 11186 0 _0235_
rlabel metal1 22356 17850 22356 17850 0 _0236_
rlabel metal1 30544 15674 30544 15674 0 _0237_
rlabel metal1 30222 17306 30222 17306 0 _0238_
rlabel metal1 26128 16422 26128 16422 0 _0239_
rlabel metal1 26956 15130 26956 15130 0 _0240_
rlabel metal1 31556 17170 31556 17170 0 _0241_
rlabel metal1 27600 17306 27600 17306 0 _0242_
rlabel metal2 17434 8432 17434 8432 0 _0243_
rlabel metal2 16514 19720 16514 19720 0 _0244_
rlabel metal2 7406 5678 7406 5678 0 _0245_
rlabel metal1 11132 7446 11132 7446 0 _0246_
rlabel metal1 17526 20026 17526 20026 0 _0247_
rlabel metal2 18354 3774 18354 3774 0 _0248_
rlabel metal2 17250 31518 17250 31518 0 _0249_
rlabel metal1 15870 32436 15870 32436 0 _0250_
rlabel metal1 9798 31382 9798 31382 0 _0251_
rlabel metal1 16652 31790 16652 31790 0 _0252_
rlabel metal1 13248 30906 13248 30906 0 _0253_
rlabel metal1 3588 25466 3588 25466 0 _0254_
rlabel metal2 14582 30906 14582 30906 0 _0255_
rlabel metal1 15318 31926 15318 31926 0 _0256_
rlabel metal2 7774 31076 7774 31076 0 _0257_
rlabel metal1 11454 30600 11454 30600 0 _0258_
rlabel metal2 13202 29580 13202 29580 0 _0259_
rlabel metal1 3174 30226 3174 30226 0 _0260_
rlabel metal2 19366 20638 19366 20638 0 _0261_
rlabel metal1 22402 19244 22402 19244 0 _0262_
rlabel metal2 14858 28322 14858 28322 0 _0263_
rlabel metal1 17848 18666 17848 18666 0 _0264_
rlabel metal2 20470 21012 20470 21012 0 _0265_
rlabel metal1 13662 28118 13662 28118 0 _0266_
rlabel metal2 29946 24174 29946 24174 0 _0267_
rlabel metal1 27922 23086 27922 23086 0 _0268_
rlabel metal1 27922 20570 27922 20570 0 _0269_
rlabel metal1 30176 24854 30176 24854 0 _0270_
rlabel metal2 29026 24820 29026 24820 0 _0271_
rlabel metal1 28750 21522 28750 21522 0 _0272_
rlabel metal1 24886 22712 24886 22712 0 _0273_
rlabel metal1 24242 23154 24242 23154 0 _0274_
rlabel metal1 27370 25772 27370 25772 0 _0275_
rlabel metal1 27324 22202 27324 22202 0 _0276_
rlabel metal2 21390 22916 21390 22916 0 _0277_
rlabel metal1 28612 26418 28612 26418 0 _0278_
rlabel metal2 16422 16082 16422 16082 0 _0279_
rlabel metal2 17986 14212 17986 14212 0 _0280_
rlabel metal2 19642 26520 19642 26520 0 _0281_
rlabel metal1 16376 22746 16376 22746 0 _0282_
rlabel metal1 16652 17170 16652 17170 0 _0283_
rlabel metal1 2392 22678 2392 22678 0 _0284_
rlabel metal2 24334 18462 24334 18462 0 _0285_
rlabel metal1 22862 17748 22862 17748 0 _0286_
rlabel metal2 21390 15028 21390 15028 0 _0287_
rlabel metal1 25346 17850 25346 17850 0 _0288_
rlabel metal2 23966 15844 23966 15844 0 _0289_
rlabel metal2 25346 19652 25346 19652 0 _0290_
rlabel metal2 20930 13022 20930 13022 0 _0291_
rlabel metal2 23138 11730 23138 11730 0 _0292_
rlabel metal2 25990 11560 25990 11560 0 _0293_
rlabel metal1 20838 11050 20838 11050 0 _0294_
rlabel metal1 20930 12274 20930 12274 0 _0295_
rlabel metal1 27094 18938 27094 18938 0 _0296_
rlabel metal1 16928 3978 16928 3978 0 _0297_
rlabel metal2 22034 8262 22034 8262 0 _0298_
rlabel metal1 26726 9690 26726 9690 0 _0299_
rlabel metal1 17756 7174 17756 7174 0 _0300_
rlabel metal2 20838 9486 20838 9486 0 _0301_
rlabel metal1 26358 17238 26358 17238 0 _0302_
rlabel metal1 24150 13498 24150 13498 0 _0303_
rlabel metal1 20056 23154 20056 23154 0 _0304_
rlabel metal2 21022 15232 21022 15232 0 _0305_
rlabel metal2 20194 21828 20194 21828 0 _0306_
rlabel metal1 21436 28050 21436 28050 0 _0307_
rlabel metal1 22218 22032 22218 22032 0 _0308_
rlabel metal2 22126 26180 22126 26180 0 _0309_
rlabel metal2 20838 26588 20838 26588 0 _0310_
rlabel metal1 13754 33524 13754 33524 0 _0311_
rlabel metal1 5290 31994 5290 31994 0 _0312_
rlabel metal1 11868 32402 11868 32402 0 _0313_
rlabel metal1 6716 31450 6716 31450 0 _0314_
rlabel metal2 15502 7344 15502 7344 0 _0315_
rlabel metal2 23414 6596 23414 6596 0 _0316_
rlabel metal1 15686 8330 15686 8330 0 _0317_
rlabel metal1 23874 7378 23874 7378 0 _0318_
rlabel metal1 2806 31926 2806 31926 0 _0319_
rlabel metal1 2300 26418 2300 26418 0 _0320_
rlabel metal2 3174 29342 3174 29342 0 _0321_
rlabel metal1 2254 25874 2254 25874 0 _0322_
rlabel metal2 11914 4284 11914 4284 0 _0323_
rlabel metal1 19826 7446 19826 7446 0 _0324_
rlabel metal2 14490 5916 14490 5916 0 _0325_
rlabel metal1 16652 20502 16652 20502 0 _0326_
rlabel metal1 29118 21114 29118 21114 0 _0327_
rlabel metal2 28290 14212 28290 14212 0 _0328_
rlabel metal1 28428 18938 28428 18938 0 _0329_
rlabel metal1 27876 18938 27876 18938 0 _0330_
rlabel metal2 23598 8738 23598 8738 0 _0331_
rlabel metal2 12282 6324 12282 6324 0 _0332_
rlabel metal2 22126 9112 22126 9112 0 _0333_
rlabel metal2 20746 9418 20746 9418 0 _0334_
rlabel metal1 17365 7718 17365 7718 0 _0335_
rlabel metal1 20700 8602 20700 8602 0 _0336_
rlabel metal1 17284 8874 17284 8874 0 _0337_
rlabel metal1 17710 8364 17710 8364 0 _0338_
rlabel metal1 19366 16150 19366 16150 0 _0339_
rlabel metal1 16008 28594 16008 28594 0 _0340_
rlabel metal1 19550 18938 19550 18938 0 _0341_
rlabel metal1 18814 27438 18814 27438 0 _0342_
rlabel metal2 13570 6256 13570 6256 0 _0343_
rlabel metal1 6440 29818 6440 29818 0 _0344_
rlabel metal1 6716 19686 6716 19686 0 _0345_
rlabel metal2 6946 30056 6946 30056 0 _0346_
rlabel metal1 18860 12954 18860 12954 0 _0347_
rlabel metal1 12650 29512 12650 29512 0 _0348_
rlabel metal1 18308 17306 18308 17306 0 _0349_
rlabel metal1 11592 27030 11592 27030 0 _0350_
rlabel metal1 18032 12886 18032 12886 0 _0351_
rlabel metal2 17250 17884 17250 17884 0 _0352_
rlabel metal1 16560 13498 16560 13498 0 _0353_
rlabel metal2 18722 22780 18722 22780 0 _0354_
rlabel metal2 22954 31620 22954 31620 0 _0355_
rlabel metal1 23644 27574 23644 27574 0 _0356_
rlabel metal2 21666 29852 21666 29852 0 _0357_
rlabel metal1 23368 29818 23368 29818 0 _0358_
rlabel metal1 17710 10234 17710 10234 0 _0359_
rlabel metal2 22862 21352 22862 21352 0 _0360_
rlabel metal1 18308 10778 18308 10778 0 _0361_
rlabel metal1 22770 12886 22770 12886 0 _0362_
rlabel metal2 5934 27608 5934 27608 0 _0363_
rlabel metal2 19366 10846 19366 10846 0 _0364_
rlabel metal1 17250 21658 17250 21658 0 _0365_
rlabel metal1 19872 9622 19872 9622 0 _0366_
rlabel metal1 7268 37230 7268 37230 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 4048 37230 4048 37230 0 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1234 27948 1234 27948 0 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 38318 11679 38318 11679 0 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel via2 38318 25245 38318 25245 0 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 22724 37230 22724 37230 0 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 10350 1588 10350 1588 0 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 15502 1588 15502 1588 0 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 32246 1588 32246 1588 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal3 1740 1428 1740 1428 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 38134 31569 38134 31569 0 ccff_head
rlabel metal2 4554 1520 4554 1520 0 ccff_tail
rlabel metal2 34178 1588 34178 1588 0 chanx_right_in[0]
rlabel metal3 1234 32708 1234 32708 0 chanx_right_in[10]
rlabel metal1 33672 37230 33672 37230 0 chanx_right_in[11]
rlabel via2 38318 19805 38318 19805 0 chanx_right_in[12]
rlabel metal1 11776 37230 11776 37230 0 chanx_right_in[13]
rlabel metal3 1924 37468 1924 37468 0 chanx_right_in[14]
rlabel metal2 3174 26129 3174 26129 0 chanx_right_in[15]
rlabel metal2 38686 1554 38686 1554 0 chanx_right_in[16]
rlabel metal3 1234 17748 1234 17748 0 chanx_right_in[17]
rlabel metal2 38318 34901 38318 34901 0 chanx_right_in[18]
rlabel metal1 37352 5678 37352 5678 0 chanx_right_in[1]
rlabel metal1 25944 37230 25944 37230 0 chanx_right_in[2]
rlabel metal3 1234 21148 1234 21148 0 chanx_right_in[3]
rlabel metal1 14996 37230 14996 37230 0 chanx_right_in[4]
rlabel metal2 16146 38226 16146 38226 0 chanx_right_in[5]
rlabel metal1 29486 37230 29486 37230 0 chanx_right_in[6]
rlabel metal3 1234 29308 1234 29308 0 chanx_right_in[7]
rlabel metal2 37490 37723 37490 37723 0 chanx_right_in[8]
rlabel metal2 38318 33439 38318 33439 0 chanx_right_in[9]
rlabel metal2 38226 36567 38226 36567 0 chanx_right_out[0]
rlabel metal2 38226 8857 38226 8857 0 chanx_right_out[10]
rlabel metal1 24334 37094 24334 37094 0 chanx_right_out[11]
rlabel metal1 18216 37094 18216 37094 0 chanx_right_out[12]
rlabel metal3 1234 4828 1234 4828 0 chanx_right_out[13]
rlabel metal1 1794 37128 1794 37128 0 chanx_right_out[14]
rlabel metal2 9062 1520 9062 1520 0 chanx_right_out[15]
rlabel metal2 38226 28815 38226 28815 0 chanx_right_out[16]
rlabel metal2 37398 1520 37398 1520 0 chanx_right_out[17]
rlabel metal2 38226 15181 38226 15181 0 chanx_right_out[18]
rlabel metal1 20838 37094 20838 37094 0 chanx_right_out[1]
rlabel metal1 13064 37094 13064 37094 0 chanx_right_out[2]
rlabel metal2 38226 1445 38226 1445 0 chanx_right_out[3]
rlabel via2 38226 30005 38226 30005 0 chanx_right_out[4]
rlabel metal1 38134 36890 38134 36890 0 chanx_right_out[5]
rlabel metal3 1234 6188 1234 6188 0 chanx_right_out[6]
rlabel metal2 13570 1520 13570 1520 0 chanx_right_out[7]
rlabel metal3 38740 6868 38740 6868 0 chanx_right_out[8]
rlabel metal3 1234 22508 1234 22508 0 chanx_right_out[9]
rlabel metal3 1234 2788 1234 2788 0 chany_bottom_in[0]
rlabel metal3 1234 30668 1234 30668 0 chany_bottom_in[10]
rlabel metal1 10488 37230 10488 37230 0 chany_bottom_in[11]
rlabel metal2 29026 1588 29026 1588 0 chany_bottom_in[12]
rlabel metal1 34960 37230 34960 37230 0 chany_bottom_in[13]
rlabel metal2 24518 1588 24518 1588 0 chany_bottom_in[14]
rlabel metal2 2622 1588 2622 1588 0 chany_bottom_in[15]
rlabel metal3 1234 19788 1234 19788 0 chany_bottom_in[16]
rlabel metal2 35466 1588 35466 1588 0 chany_bottom_in[17]
rlabel metal2 38318 17119 38318 17119 0 chany_bottom_in[18]
rlabel metal2 38318 10455 38318 10455 0 chany_bottom_in[1]
rlabel metal2 27738 1588 27738 1588 0 chany_bottom_in[2]
rlabel metal3 1234 34068 1234 34068 0 chany_bottom_in[3]
rlabel metal2 36938 2567 36938 2567 0 chany_bottom_in[4]
rlabel metal1 5336 37230 5336 37230 0 chany_bottom_in[5]
rlabel metal2 38318 13787 38318 13787 0 chany_bottom_in[6]
rlabel metal3 1234 16388 1234 16388 0 chany_bottom_in[7]
rlabel metal2 30958 1588 30958 1588 0 chany_bottom_in[8]
rlabel metal2 38318 26775 38318 26775 0 chany_bottom_in[9]
rlabel metal2 18722 1520 18722 1520 0 chany_bottom_out[0]
rlabel metal2 1794 24463 1794 24463 0 chany_bottom_out[10]
rlabel metal2 20010 1520 20010 1520 0 chany_bottom_out[11]
rlabel metal2 46 1792 46 1792 0 chany_bottom_out[12]
rlabel metal2 23230 1520 23230 1520 0 chany_bottom_out[13]
rlabel metal3 1234 8228 1234 8228 0 chany_bottom_out[14]
rlabel metal1 19504 37094 19504 37094 0 chany_bottom_out[15]
rlabel metal3 1234 12988 1234 12988 0 chany_bottom_out[16]
rlabel metal1 1242 36890 1242 36890 0 chany_bottom_out[17]
rlabel metal2 5842 1520 5842 1520 0 chany_bottom_out[18]
rlabel metal2 1334 1520 1334 1520 0 chany_bottom_out[1]
rlabel metal1 36800 37094 36800 37094 0 chany_bottom_out[2]
rlabel metal1 27232 37094 27232 37094 0 chany_bottom_out[3]
rlabel metal2 16790 1520 16790 1520 0 chany_bottom_out[4]
rlabel metal1 37720 37434 37720 37434 0 chany_bottom_out[5]
rlabel metal2 38226 3417 38226 3417 0 chany_bottom_out[6]
rlabel metal3 1234 9588 1234 9588 0 chany_bottom_out[7]
rlabel via2 38226 21845 38226 21845 0 chany_bottom_out[8]
rlabel metal2 7774 1520 7774 1520 0 chany_bottom_out[9]
rlabel metal2 1886 9282 1886 9282 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal2 3358 8874 3358 8874 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal2 17710 8058 17710 8058 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal1 18170 20434 18170 20434 0 mem_bottom_track_11.DFFR_0_.D
rlabel metal1 22218 23800 22218 23800 0 mem_bottom_track_11.DFFR_0_.Q
rlabel metal2 28566 23052 28566 23052 0 mem_bottom_track_11.DFFR_1_.Q
rlabel metal2 25438 23358 25438 23358 0 mem_bottom_track_13.DFFR_0_.Q
rlabel metal2 23598 21794 23598 21794 0 mem_bottom_track_13.DFFR_1_.Q
rlabel metal2 2530 22270 2530 22270 0 mem_bottom_track_15.DFFR_0_.Q
rlabel metal1 1886 16184 1886 16184 0 mem_bottom_track_15.DFFR_1_.Q
rlabel metal1 25576 19346 25576 19346 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal2 25070 17850 25070 17850 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal1 25990 12206 25990 12206 0 mem_bottom_track_19.DFFR_0_.Q
rlabel metal1 22218 12172 22218 12172 0 mem_bottom_track_19.DFFR_1_.Q
rlabel metal1 9338 9350 9338 9350 0 mem_bottom_track_23.DFFR_0_.Q
rlabel metal1 18952 18734 18952 18734 0 mem_bottom_track_23.DFFR_1_.Q
rlabel metal1 5191 21114 5191 21114 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal1 9844 12206 9844 12206 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal1 9200 17306 9200 17306 0 mem_bottom_track_27.DFFR_0_.Q
rlabel metal2 18354 11084 18354 11084 0 mem_bottom_track_27.DFFR_1_.Q
rlabel metal1 16514 18258 16514 18258 0 mem_bottom_track_29.DFFR_0_.Q
rlabel metal1 7636 16422 7636 16422 0 mem_bottom_track_29.DFFR_1_.Q
rlabel via2 16790 9333 16790 9333 0 mem_bottom_track_3.DFFR_0_.Q
rlabel metal1 5658 11866 5658 11866 0 mem_bottom_track_3.DFFR_1_.Q
rlabel metal2 23046 28832 23046 28832 0 mem_bottom_track_31.DFFR_0_.Q
rlabel metal2 22494 30770 22494 30770 0 mem_bottom_track_31.DFFR_1_.Q
rlabel metal1 22770 16762 22770 16762 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal1 17434 8942 17434 8942 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal1 18814 10098 18814 10098 0 mem_bottom_track_35.DFFR_0_.Q
rlabel metal1 10994 9622 10994 9622 0 mem_bottom_track_35.DFFR_1_.Q
rlabel metal2 6854 10336 6854 10336 0 mem_bottom_track_37.DFFR_0_.Q
rlabel metal1 11132 32402 11132 32402 0 mem_bottom_track_5.DFFR_0_.Q
rlabel metal2 16422 32096 16422 32096 0 mem_bottom_track_5.DFFR_1_.Q
rlabel metal1 2346 24718 2346 24718 0 mem_bottom_track_7.DFFR_0_.Q
rlabel metal1 12834 19244 12834 19244 0 mem_bottom_track_7.DFFR_1_.Q
rlabel metal2 22770 20094 22770 20094 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal1 22816 24786 22816 24786 0 mem_right_track_0.DFFR_0_.Q
rlabel metal1 24564 25262 24564 25262 0 mem_right_track_0.DFFR_1_.Q
rlabel metal2 22356 24174 22356 24174 0 mem_right_track_10.DFFR_0_.D
rlabel metal1 23138 24208 23138 24208 0 mem_right_track_10.DFFR_0_.Q
rlabel metal1 25622 23052 25622 23052 0 mem_right_track_10.DFFR_1_.Q
rlabel metal2 12558 21760 12558 21760 0 mem_right_track_12.DFFR_0_.Q
rlabel metal1 8326 27064 8326 27064 0 mem_right_track_12.DFFR_1_.Q
rlabel metal1 21068 16082 21068 16082 0 mem_right_track_14.DFFR_0_.Q
rlabel metal2 18078 15266 18078 15266 0 mem_right_track_14.DFFR_1_.Q
rlabel metal1 28658 18258 28658 18258 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 28382 13362 28382 13362 0 mem_right_track_16.DFFR_1_.Q
rlabel metal1 25254 16082 25254 16082 0 mem_right_track_18.DFFR_0_.Q
rlabel metal2 21114 16932 21114 16932 0 mem_right_track_18.DFFR_1_.Q
rlabel metal1 19688 28050 19688 28050 0 mem_right_track_2.DFFR_0_.Q
rlabel metal1 16882 30702 16882 30702 0 mem_right_track_2.DFFR_1_.Q
rlabel metal1 13248 16150 13248 16150 0 mem_right_track_20.DFFR_0_.Q
rlabel metal2 24702 14416 24702 14416 0 mem_right_track_20.DFFR_1_.Q
rlabel metal1 24426 21454 24426 21454 0 mem_right_track_22.DFFR_0_.Q
rlabel metal1 14352 23834 14352 23834 0 mem_right_track_22.DFFR_1_.Q
rlabel metal2 3726 22848 3726 22848 0 mem_right_track_24.DFFR_0_.Q
rlabel metal1 11960 33490 11960 33490 0 mem_right_track_24.DFFR_1_.Q
rlabel metal1 23736 6766 23736 6766 0 mem_right_track_26.DFFR_0_.Q
rlabel metal1 3266 9996 3266 9996 0 mem_right_track_26.DFFR_1_.Q
rlabel metal1 4186 10166 4186 10166 0 mem_right_track_28.DFFR_0_.Q
rlabel metal1 2530 31790 2530 31790 0 mem_right_track_28.DFFR_1_.Q
rlabel metal1 17618 6664 17618 6664 0 mem_right_track_30.DFFR_0_.Q
rlabel metal1 5428 11050 5428 11050 0 mem_right_track_30.DFFR_1_.Q
rlabel metal1 8004 11254 8004 11254 0 mem_right_track_32.DFFR_0_.Q
rlabel metal1 28934 18734 28934 18734 0 mem_right_track_32.DFFR_1_.Q
rlabel metal1 13662 5746 13662 5746 0 mem_right_track_34.DFFR_0_.Q
rlabel metal2 6394 9792 6394 9792 0 mem_right_track_34.DFFR_1_.Q
rlabel metal2 17618 12036 17618 12036 0 mem_right_track_36.DFFR_0_.Q
rlabel metal1 8142 5678 8142 5678 0 mem_right_track_4.DFFR_0_.Q
rlabel metal1 10764 18666 10764 18666 0 mem_right_track_4.DFFR_1_.Q
rlabel metal1 24150 20910 24150 20910 0 mem_right_track_6.DFFR_0_.Q
rlabel metal1 22724 11118 22724 11118 0 mem_right_track_6.DFFR_1_.Q
rlabel metal1 22356 19822 22356 19822 0 mem_right_track_8.DFFR_0_.Q
rlabel metal2 2438 5950 2438 5950 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 23828 9962 23828 9962 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 20286 8534 20286 8534 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17388 3026 17388 3026 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 17618 3332 17618 3332 0 mux_bottom_track_1.out
rlabel metal1 30130 21454 30130 21454 0 mux_bottom_track_11.INVTX1_0_.out
rlabel metal1 27968 20978 27968 20978 0 mux_bottom_track_11.INVTX1_1_.out
rlabel metal1 23690 27948 23690 27948 0 mux_bottom_track_11.INVTX1_2_.out
rlabel metal2 29578 23188 29578 23188 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 29854 23460 29854 23460 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 30498 24242 30498 24242 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 33074 30294 33074 30294 0 mux_bottom_track_11.out
rlabel metal2 27922 28492 27922 28492 0 mux_bottom_track_13.INVTX1_0_.out
rlabel metal2 22218 22372 22218 22372 0 mux_bottom_track_13.INVTX1_2_.out
rlabel metal2 27646 24106 27646 24106 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23276 23222 23276 23222 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 27738 21505 27738 21505 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 33166 10234 33166 10234 0 mux_bottom_track_13.out
rlabel metal1 2070 22542 2070 22542 0 mux_bottom_track_15.INVTX1_0_.out
rlabel metal2 16698 5031 16698 5031 0 mux_bottom_track_15.INVTX1_2_.out
rlabel metal1 16422 23188 16422 23188 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17526 16048 17526 16048 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15916 9078 15916 9078 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 4738 8976 4738 8976 0 mux_bottom_track_15.out
rlabel metal1 24610 19958 24610 19958 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal1 18906 6222 18906 6222 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal2 25438 18938 25438 18938 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23782 17510 23782 17510 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25714 18156 25714 18156 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 31142 20740 31142 20740 0 mux_bottom_track_17.out
rlabel metal1 26956 27302 26956 27302 0 mux_bottom_track_19.INVTX1_0_.out
rlabel metal2 25806 11458 25806 11458 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 20838 12954 20838 12954 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 21206 7242 21206 7242 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 11086 3196 11086 3196 0 mux_bottom_track_19.out
rlabel metal2 20838 27676 20838 27676 0 mux_bottom_track_23.INVTX1_0_.out
rlabel metal1 15732 28594 15732 28594 0 mux_bottom_track_23.INVTX1_1_.out
rlabel metal1 19366 19278 19366 19278 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18814 6290 18814 6290 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 18906 5882 18906 5882 0 mux_bottom_track_23.out
rlabel metal2 11086 30668 11086 30668 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal2 7774 32062 7774 32062 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal1 5152 21318 5152 21318 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 4140 7378 4140 7378 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 4508 5678 4508 5678 0 mux_bottom_track_25.out
rlabel metal1 14490 32198 14490 32198 0 mux_bottom_track_27.INVTX1_0_.out
rlabel metal2 13018 28832 13018 28832 0 mux_bottom_track_27.INVTX1_1_.out
rlabel metal1 15364 17782 15364 17782 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 19320 11084 19320 11084 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 20562 8092 20562 8092 0 mux_bottom_track_27.out
rlabel metal2 13938 19040 13938 19040 0 mux_bottom_track_29.INVTX1_0_.out
rlabel metal1 18308 17850 18308 17850 0 mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 5842 8500 5842 8500 0 mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 6348 8466 6348 8466 0 mux_bottom_track_29.out
rlabel metal2 27830 3706 27830 3706 0 mux_bottom_track_3.INVTX1_0_.out
rlabel metal2 7314 4148 7314 4148 0 mux_bottom_track_3.INVTX1_1_.out
rlabel metal1 9982 5134 9982 5134 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17158 9452 17158 9452 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 5658 6324 5658 6324 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 5014 6256 5014 6256 0 mux_bottom_track_3.out
rlabel metal2 23874 30294 23874 30294 0 mux_bottom_track_31.INVTX1_0_.out
rlabel metal2 24058 29376 24058 29376 0 mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21620 29818 21620 29818 0 mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 19320 32402 19320 32402 0 mux_bottom_track_31.out
rlabel metal1 22126 12920 22126 12920 0 mux_bottom_track_33.INVTX1_0_.out
rlabel metal1 22448 21454 22448 21454 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18032 11050 18032 11050 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 2898 6800 2898 6800 0 mux_bottom_track_33.out
rlabel metal2 25070 10336 25070 10336 0 mux_bottom_track_35.INVTX1_0_.out
rlabel metal1 19964 11730 19964 11730 0 mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 5106 32878 5106 32878 0 mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 3082 32912 3082 32912 0 mux_bottom_track_35.out
rlabel metal2 25990 21998 25990 21998 0 mux_bottom_track_37.INVTX1_0_.out
rlabel metal2 17802 6426 17802 6426 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19872 8806 19872 8806 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 18262 6698 18262 6698 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 6670 4250 6670 4250 0 mux_bottom_track_37.out
rlabel metal2 3542 26690 3542 26690 0 mux_bottom_track_5.INVTX1_0_.out
rlabel metal1 14674 30226 14674 30226 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16054 32096 16054 32096 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 21758 31926 21758 31926 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30176 36142 30176 36142 0 mux_bottom_track_5.out
rlabel metal1 3772 30158 3772 30158 0 mux_bottom_track_7.INVTX1_0_.out
rlabel metal1 6624 31110 6624 31110 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 14490 29954 14490 29954 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 19504 32334 19504 32334 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 21528 32538 21528 32538 0 mux_bottom_track_7.out
rlabel metal1 13846 27982 13846 27982 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 16698 18598 16698 18598 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 19274 19924 19274 19924 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17066 7480 17066 7480 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 16192 7174 16192 7174 0 mux_bottom_track_9.out
rlabel metal1 24058 18326 24058 18326 0 mux_right_track_0.INVTX1_0_.out
rlabel metal1 23368 24718 23368 24718 0 mux_right_track_0.INVTX1_1_.out
rlabel metal1 29348 9622 29348 9622 0 mux_right_track_0.INVTX1_2_.out
rlabel metal1 24012 24922 24012 24922 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 28704 23562 28704 23562 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 27968 23766 27968 23766 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 36478 31926 36478 31926 0 mux_right_track_0.out
rlabel metal1 2438 33286 2438 33286 0 mux_right_track_10.INVTX1_0_.out
rlabel metal1 17710 23630 17710 23630 0 mux_right_track_10.INVTX1_1_.out
rlabel metal1 24794 14892 24794 14892 0 mux_right_track_10.INVTX1_2_.out
rlabel metal2 21390 23936 21390 23936 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 25484 23630 25484 23630 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 27462 24242 27462 24242 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 33902 35802 33902 35802 0 mux_right_track_10.out
rlabel metal1 28428 19346 28428 19346 0 mux_right_track_12.INVTX1_1_.out
rlabel metal1 9522 31858 9522 31858 0 mux_right_track_12.INVTX1_2_.out
rlabel metal1 18538 21862 18538 21862 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17618 27540 17618 27540 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 6026 6817 6026 6817 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 6026 7174 6026 7174 0 mux_right_track_12.out
rlabel metal1 23138 17272 23138 17272 0 mux_right_track_14.INVTX1_1_.out
rlabel metal2 3358 26588 3358 26588 0 mux_right_track_14.INVTX1_2_.out
rlabel metal2 20654 17612 20654 17612 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal3 18791 16524 18791 16524 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 18446 6051 18446 6051 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 14030 5168 14030 5168 0 mux_right_track_14.out
rlabel metal1 24426 17136 24426 17136 0 mux_right_track_16.INVTX1_1_.out
rlabel metal1 30084 20434 30084 20434 0 mux_right_track_16.INVTX1_2_.out
rlabel metal1 28290 12750 28290 12750 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 30452 18938 30452 18938 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 30866 13192 30866 13192 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 32522 11900 32522 11900 0 mux_right_track_16.out
rlabel metal1 24886 11084 24886 11084 0 mux_right_track_18.INVTX1_2_.out
rlabel metal1 22678 18054 22678 18054 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23322 11594 23322 11594 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 20884 17782 20884 17782 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel via2 1978 20451 1978 20451 0 mux_right_track_18.out
rlabel metal1 18492 29682 18492 29682 0 mux_right_track_2.INVTX1_1_.out
rlabel metal2 4094 25874 4094 25874 0 mux_right_track_2.INVTX1_2_.out
rlabel metal2 20102 29104 20102 29104 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16882 28084 16882 28084 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 19182 28594 19182 28594 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 19642 29818 19642 29818 0 mux_right_track_2.out
rlabel metal3 2047 31756 2047 31756 0 mux_right_track_20.INVTX1_1_.out
rlabel metal1 20056 15538 20056 15538 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24058 14008 24058 14008 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 31418 10506 31418 10506 0 mux_right_track_20.out
rlabel metal2 33626 16473 33626 16473 0 mux_right_track_22.INVTX1_1_.out
rlabel metal1 21252 22066 21252 22066 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22770 29444 22770 29444 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 22862 32198 22862 32198 0 mux_right_track_22.out
rlabel metal2 23138 20128 23138 20128 0 mux_right_track_24.INVTX1_0_.out
rlabel metal1 5014 32334 5014 32334 0 mux_right_track_24.INVTX1_1_.out
rlabel metal1 9476 32470 9476 32470 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 13938 32912 13938 32912 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 17434 34000 17434 34000 0 mux_right_track_24.out
rlabel metal1 24932 6426 24932 6426 0 mux_right_track_26.INVTX1_0_.out
rlabel metal1 22678 6732 22678 6732 0 mux_right_track_26.INVTX1_1_.out
rlabel metal1 23414 6630 23414 6630 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13524 6154 13524 6154 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 6762 6596 6762 6596 0 mux_right_track_26.out
rlabel metal2 1886 26588 1886 26588 0 mux_right_track_28.INVTX1_1_.out
rlabel metal2 3082 27268 3082 27268 0 mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 2484 33422 2484 33422 0 mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 1978 34102 1978 34102 0 mux_right_track_28.out
rlabel metal1 22908 6834 22908 6834 0 mux_right_track_30.INVTX1_1_.out
rlabel metal2 19366 6290 19366 6290 0 mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12052 5202 12052 5202 0 mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 9706 3060 9706 3060 0 mux_right_track_30.out
rlabel metal2 29946 13974 29946 13974 0 mux_right_track_32.INVTX1_1_.out
rlabel metal1 28842 19346 28842 19346 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 28934 23664 28934 23664 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 32798 25262 32798 25262 0 mux_right_track_32.out
rlabel metal1 7314 5780 7314 5780 0 mux_right_track_34.INVTX1_1_.out
rlabel metal1 21528 8874 21528 8874 0 mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23506 9044 23506 9044 0 mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 30268 7718 30268 7718 0 mux_right_track_34.out
rlabel metal2 32430 16932 32430 16932 0 mux_right_track_36.INVTX1_2_.out
rlabel metal1 27462 17782 27462 17782 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 31050 17408 31050 17408 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 31050 15538 31050 15538 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 32522 15436 32522 15436 0 mux_right_track_36.out
rlabel metal2 5842 6426 5842 6426 0 mux_right_track_4.INVTX1_2_.out
rlabel metal2 10534 29274 10534 29274 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 10626 6222 10626 6222 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 10764 29070 10764 29070 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 11316 31790 11316 31790 0 mux_right_track_4.out
rlabel metal1 24334 8058 24334 8058 0 mux_right_track_6.INVTX1_2_.out
rlabel metal1 23184 20230 23184 20230 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 25438 9894 25438 9894 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 24150 9690 24150 9690 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 31418 5270 31418 5270 0 mux_right_track_6.out
rlabel metal2 25070 30124 25070 30124 0 mux_right_track_8.INVTX1_2_.out
rlabel metal2 23230 20281 23230 20281 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 25208 28186 25208 28186 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 24104 22066 24104 22066 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 33902 30226 33902 30226 0 mux_right_track_8.out
rlabel metal1 7912 31314 7912 31314 0 net1
rlabel metal1 6578 2992 6578 2992 0 net10
rlabel metal2 28474 15776 28474 15776 0 net100
rlabel metal1 18216 27506 18216 27506 0 net101
rlabel metal2 11822 19550 11822 19550 0 net102
rlabel metal2 25162 8160 25162 8160 0 net103
rlabel metal1 23736 29070 23736 29070 0 net104
rlabel metal2 24610 15776 24610 15776 0 net105
rlabel metal2 17342 26656 17342 26656 0 net106
rlabel metal1 18860 25330 18860 25330 0 net107
rlabel metal2 29670 18564 29670 18564 0 net108
rlabel metal2 23230 11900 23230 11900 0 net109
rlabel metal1 24702 26520 24702 26520 0 net11
rlabel metal1 30682 17714 30682 17714 0 net110
rlabel metal1 16652 18802 16652 18802 0 net111
rlabel metal2 15686 32572 15686 32572 0 net112
rlabel metal2 15594 31008 15594 31008 0 net113
rlabel metal2 20654 19040 20654 19040 0 net114
rlabel metal1 27922 23154 27922 23154 0 net115
rlabel metal2 23322 23392 23322 23392 0 net116
rlabel metal1 17112 14450 17112 14450 0 net117
rlabel metal2 22678 18156 22678 18156 0 net118
rlabel metal1 19734 13362 19734 13362 0 net119
rlabel metal2 26174 5644 26174 5644 0 net12
rlabel metal1 19320 9010 19320 9010 0 net120
rlabel metal2 23414 13600 23414 13600 0 net121
rlabel metal2 20838 28220 20838 28220 0 net122
rlabel metal2 13570 33660 13570 33660 0 net123
rlabel metal2 14490 7650 14490 7650 0 net124
rlabel metal2 2806 29886 2806 29886 0 net125
rlabel metal1 11454 4114 11454 4114 0 net126
rlabel metal2 28382 22304 28382 22304 0 net127
rlabel metal2 23230 9248 23230 9248 0 net128
rlabel metal1 15962 7786 15962 7786 0 net129
rlabel metal2 1886 31178 1886 31178 0 net13
rlabel metal2 18722 15776 18722 15776 0 net130
rlabel metal2 9246 7072 9246 7072 0 net131
rlabel metal2 18906 14110 18906 14110 0 net132
rlabel metal2 17342 12512 17342 12512 0 net133
rlabel metal2 20746 31620 20746 31620 0 net134
rlabel metal2 17526 11424 17526 11424 0 net135
rlabel metal2 5842 27744 5842 27744 0 net136
rlabel metal1 33028 37094 33028 37094 0 net14
rlabel metal2 33074 20774 33074 20774 0 net15
rlabel metal2 14306 29852 14306 29852 0 net16
rlabel metal1 3450 37094 3450 37094 0 net17
rlabel metal1 1978 25296 1978 25296 0 net18
rlabel metal2 35650 3604 35650 3604 0 net19
rlabel metal1 5428 37162 5428 37162 0 net2
rlabel metal1 1978 18054 1978 18054 0 net20
rlabel metal2 37306 30940 37306 30940 0 net21
rlabel metal1 32062 5746 32062 5746 0 net22
rlabel metal1 24840 37162 24840 37162 0 net23
rlabel metal2 2438 20026 2438 20026 0 net24
rlabel metal1 14858 37094 14858 37094 0 net25
rlabel metal1 16744 37094 16744 37094 0 net26
rlabel metal2 29762 32606 29762 32606 0 net27
rlabel metal2 1978 28730 1978 28730 0 net28
rlabel metal2 37766 32334 37766 32334 0 net29
rlabel metal2 4002 28594 4002 28594 0 net3
rlabel metal2 29486 29580 29486 29580 0 net30
rlabel metal1 2208 3706 2208 3706 0 net31
rlabel metal1 1748 28050 1748 28050 0 net32
rlabel metal1 10074 31790 10074 31790 0 net33
rlabel metal1 28750 11118 28750 11118 0 net34
rlabel metal1 34776 37094 34776 37094 0 net35
rlabel metal1 24242 2618 24242 2618 0 net36
rlabel metal1 3726 2618 3726 2618 0 net37
rlabel metal1 2254 20026 2254 20026 0 net38
rlabel metal1 34316 2618 34316 2618 0 net39
rlabel metal2 32430 13668 32430 13668 0 net4
rlabel metal1 37030 16966 37030 16966 0 net40
rlabel metal1 37536 10778 37536 10778 0 net41
rlabel metal1 27692 2618 27692 2618 0 net42
rlabel metal1 1794 26962 1794 26962 0 net43
rlabel metal2 36754 4420 36754 4420 0 net44
rlabel metal1 4968 37094 4968 37094 0 net45
rlabel metal1 37628 14042 37628 14042 0 net46
rlabel metal1 1564 16422 1564 16422 0 net47
rlabel metal1 29486 2550 29486 2550 0 net48
rlabel metal1 37720 26758 37720 26758 0 net49
rlabel metal2 38134 25636 38134 25636 0 net5
rlabel metal2 10166 3876 10166 3876 0 net50
rlabel metal2 36478 21964 36478 21964 0 net51
rlabel metal1 21666 2618 21666 2618 0 net52
rlabel metal1 29900 37162 29900 37162 0 net53
rlabel metal1 24610 27506 24610 27506 0 net54
rlabel metal2 2346 33116 2346 33116 0 net55
rlabel metal2 9154 34986 9154 34986 0 net56
rlabel metal2 27186 4454 27186 4454 0 net57
rlabel metal1 1794 11186 1794 11186 0 net58
rlabel metal1 2576 36006 2576 36006 0 net59
rlabel metal1 21850 37094 21850 37094 0 net6
rlabel metal1 37007 18598 37007 18598 0 net60
rlabel metal1 4646 2448 4646 2448 0 net61
rlabel metal1 37766 34714 37766 34714 0 net62
rlabel metal2 32890 9418 32890 9418 0 net63
rlabel metal1 23966 37230 23966 37230 0 net64
rlabel metal1 17710 37230 17710 37230 0 net65
rlabel metal1 6532 6630 6532 6630 0 net66
rlabel metal1 1702 34714 1702 34714 0 net67
rlabel metal2 9154 2618 9154 2618 0 net68
rlabel metal1 37352 29138 37352 29138 0 net69
rlabel metal1 10810 2618 10810 2618 0 net7
rlabel metal1 37490 2448 37490 2448 0 net70
rlabel metal1 36961 15470 36961 15470 0 net71
rlabel metal1 20792 37230 20792 37230 0 net72
rlabel metal1 12512 37230 12512 37230 0 net73
rlabel metal1 38042 3060 38042 3060 0 net74
rlabel metal1 36961 30226 36961 30226 0 net75
rlabel metal1 36961 36754 36961 36754 0 net76
rlabel metal1 3588 6358 3588 6358 0 net77
rlabel metal2 14306 3706 14306 3706 0 net78
rlabel metal2 34086 9452 34086 9452 0 net79
rlabel metal2 17158 4454 17158 4454 0 net8
rlabel metal1 1702 20570 1702 20570 0 net80
rlabel metal2 18630 2890 18630 2890 0 net81
rlabel metal1 1794 24174 1794 24174 0 net82
rlabel metal2 20102 3978 20102 3978 0 net83
rlabel metal1 1610 3060 1610 3060 0 net84
rlabel metal1 22172 6630 22172 6630 0 net85
rlabel metal1 1610 8534 1610 8534 0 net86
rlabel metal1 19228 37230 19228 37230 0 net87
rlabel metal1 2162 13294 2162 13294 0 net88
rlabel metal1 2254 36754 2254 36754 0 net89
rlabel metal1 29762 10574 29762 10574 0 net9
rlabel metal2 6578 2890 6578 2890 0 net90
rlabel metal1 1610 2482 1610 2482 0 net91
rlabel metal2 36662 36788 36662 36788 0 net92
rlabel metal1 25162 33082 25162 33082 0 net93
rlabel metal2 16790 4522 16790 4522 0 net94
rlabel metal1 35696 37230 35696 37230 0 net95
rlabel metal2 38042 6698 38042 6698 0 net96
rlabel metal1 4600 9146 4600 9146 0 net97
rlabel metal2 30958 21556 30958 21556 0 net98
rlabel metal1 8096 2414 8096 2414 0 net99
rlabel metal2 12282 1588 12282 1588 0 pReset
rlabel metal1 1978 18190 1978 18190 0 prog_clk
rlabel metal2 38318 23443 38318 23443 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 21298 1588 21298 1588 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 32154 37230 32154 37230 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 30498 37230 30498 37230 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 2254 37230 2254 37230 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 8878 37230 8878 37230 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 26450 1588 26450 1588 0 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal3 1142 10948 1142 10948 0 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal3 1234 36108 1234 36108 0 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 38318 18581 38318 18581 0 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
