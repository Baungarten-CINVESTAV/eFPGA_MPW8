magic
tech sky130A
magscale 1 2
timestamp 1672417252
<< viali >>
rect 7205 37281 7239 37315
rect 1593 37213 1627 37247
rect 2513 37213 2547 37247
rect 3157 37213 3191 37247
rect 3985 37213 4019 37247
rect 5273 37213 5307 37247
rect 7481 37213 7515 37247
rect 9321 37213 9355 37247
rect 10609 37213 10643 37247
rect 11897 37213 11931 37247
rect 13185 37213 13219 37247
rect 14933 37213 14967 37247
rect 16865 37213 16899 37247
rect 18153 37213 18187 37247
rect 19441 37213 19475 37247
rect 20913 37213 20947 37247
rect 22845 37213 22879 37247
rect 24593 37213 24627 37247
rect 25881 37213 25915 37247
rect 27353 37213 27387 37247
rect 29745 37213 29779 37247
rect 30665 37213 30699 37247
rect 32505 37213 32539 37247
rect 33793 37213 33827 37247
rect 35081 37213 35115 37247
rect 36921 37213 36955 37247
rect 38025 37213 38059 37247
rect 1777 37077 1811 37111
rect 2329 37077 2363 37111
rect 2973 37077 3007 37111
rect 4169 37077 4203 37111
rect 5457 37077 5491 37111
rect 9137 37077 9171 37111
rect 10425 37077 10459 37111
rect 11713 37077 11747 37111
rect 13001 37077 13035 37111
rect 15117 37077 15151 37111
rect 17049 37077 17083 37111
rect 18337 37077 18371 37111
rect 19625 37077 19659 37111
rect 20729 37077 20763 37111
rect 22661 37077 22695 37111
rect 24777 37077 24811 37111
rect 26065 37077 26099 37111
rect 27169 37077 27203 37111
rect 29929 37077 29963 37111
rect 30481 37077 30515 37111
rect 32321 37077 32355 37111
rect 33609 37077 33643 37111
rect 34897 37077 34931 37111
rect 36737 37077 36771 37111
rect 38209 37077 38243 37111
rect 1777 36873 1811 36907
rect 2329 36873 2363 36907
rect 38209 36873 38243 36907
rect 1593 36737 1627 36771
rect 2513 36737 2547 36771
rect 36921 36737 36955 36771
rect 38025 36737 38059 36771
rect 36737 36533 36771 36567
rect 1777 36125 1811 36159
rect 38301 36125 38335 36159
rect 1593 35989 1627 36023
rect 38117 35989 38151 36023
rect 2513 35785 2547 35819
rect 2421 35649 2455 35683
rect 5733 35241 5767 35275
rect 15117 35241 15151 35275
rect 16497 35241 16531 35275
rect 17417 35241 17451 35275
rect 21097 35241 21131 35275
rect 23213 35241 23247 35275
rect 5917 35037 5951 35071
rect 12081 35037 12115 35071
rect 15301 35037 15335 35071
rect 16681 35037 16715 35071
rect 17601 35037 17635 35071
rect 21281 35037 21315 35071
rect 23397 35037 23431 35071
rect 30481 35037 30515 35071
rect 38025 35037 38059 35071
rect 12173 34901 12207 34935
rect 30573 34901 30607 34935
rect 38209 34901 38243 34935
rect 7941 34697 7975 34731
rect 18337 34697 18371 34731
rect 27169 34697 27203 34731
rect 1593 34561 1627 34595
rect 8125 34561 8159 34595
rect 11989 34561 12023 34595
rect 18521 34561 18555 34595
rect 19901 34561 19935 34595
rect 27353 34561 27387 34595
rect 33241 34561 33275 34595
rect 12081 34493 12115 34527
rect 19993 34493 20027 34527
rect 33333 34493 33367 34527
rect 1777 34357 1811 34391
rect 7205 34153 7239 34187
rect 25973 34153 26007 34187
rect 34897 34153 34931 34187
rect 7113 33949 7147 33983
rect 21741 33949 21775 33983
rect 25881 33949 25915 33983
rect 29745 33949 29779 33983
rect 35081 33949 35115 33983
rect 21833 33813 21867 33847
rect 29837 33813 29871 33847
rect 10793 33473 10827 33507
rect 38025 33473 38059 33507
rect 38209 33337 38243 33371
rect 10885 33269 10919 33303
rect 1777 32861 1811 32895
rect 1593 32725 1627 32759
rect 34713 32521 34747 32555
rect 6561 32385 6595 32419
rect 23213 32385 23247 32419
rect 34897 32385 34931 32419
rect 6653 32181 6687 32215
rect 23305 32181 23339 32215
rect 9873 31977 9907 32011
rect 26065 31909 26099 31943
rect 38117 31909 38151 31943
rect 29837 31841 29871 31875
rect 8401 31773 8435 31807
rect 8493 31773 8527 31807
rect 9137 31773 9171 31807
rect 9229 31773 9263 31807
rect 9781 31773 9815 31807
rect 25145 31773 25179 31807
rect 25237 31773 25271 31807
rect 25973 31773 26007 31807
rect 29745 31773 29779 31807
rect 38301 31773 38335 31807
rect 30757 31297 30791 31331
rect 30849 31093 30883 31127
rect 4169 30889 4203 30923
rect 17325 30889 17359 30923
rect 34897 30889 34931 30923
rect 1777 30685 1811 30719
rect 4353 30685 4387 30719
rect 17233 30685 17267 30719
rect 35081 30685 35115 30719
rect 1593 30549 1627 30583
rect 15669 30277 15703 30311
rect 15577 30209 15611 30243
rect 38301 30209 38335 30243
rect 38117 30005 38151 30039
rect 6101 29801 6135 29835
rect 17233 29801 17267 29835
rect 19533 29801 19567 29835
rect 22017 29801 22051 29835
rect 34897 29801 34931 29835
rect 1593 29597 1627 29631
rect 3985 29597 4019 29631
rect 6009 29597 6043 29631
rect 17141 29597 17175 29631
rect 19441 29597 19475 29631
rect 21925 29597 21959 29631
rect 35081 29597 35115 29631
rect 1777 29461 1811 29495
rect 4077 29461 4111 29495
rect 18061 29257 18095 29291
rect 29193 29257 29227 29291
rect 17969 29121 18003 29155
rect 29101 29121 29135 29155
rect 38025 29121 38059 29155
rect 38209 28985 38243 29019
rect 29837 28713 29871 28747
rect 6929 28509 6963 28543
rect 29745 28509 29779 28543
rect 7021 28373 7055 28407
rect 1777 28033 1811 28067
rect 32321 28033 32355 28067
rect 1593 27829 1627 27863
rect 32413 27829 32447 27863
rect 7481 27421 7515 27455
rect 34161 27421 34195 27455
rect 7573 27285 7607 27319
rect 34253 27285 34287 27319
rect 38025 26945 38059 26979
rect 38209 26741 38243 26775
rect 29837 26537 29871 26571
rect 1593 26469 1627 26503
rect 1777 26333 1811 26367
rect 29745 26333 29779 26367
rect 4077 25993 4111 26027
rect 4261 25857 4295 25891
rect 28825 25449 28859 25483
rect 28733 25245 28767 25279
rect 38301 25245 38335 25279
rect 38117 25109 38151 25143
rect 1593 24769 1627 24803
rect 19073 24769 19107 24803
rect 34989 24769 35023 24803
rect 17141 24701 17175 24735
rect 19257 24701 19291 24735
rect 20177 24701 20211 24735
rect 34805 24633 34839 24667
rect 1777 24565 1811 24599
rect 19441 24565 19475 24599
rect 18153 24361 18187 24395
rect 19993 24225 20027 24259
rect 20637 24225 20671 24259
rect 16865 24157 16899 24191
rect 17325 24157 17359 24191
rect 18061 24157 18095 24191
rect 18889 24157 18923 24191
rect 20085 24089 20119 24123
rect 16681 24021 16715 24055
rect 17417 24021 17451 24055
rect 18705 24021 18739 24055
rect 16129 23817 16163 23851
rect 18337 23817 18371 23851
rect 34805 23817 34839 23851
rect 17141 23749 17175 23783
rect 17233 23749 17267 23783
rect 19073 23749 19107 23783
rect 19809 23749 19843 23783
rect 20361 23749 20395 23783
rect 7757 23681 7791 23715
rect 13185 23681 13219 23715
rect 15485 23681 15519 23715
rect 16313 23681 16347 23715
rect 18521 23681 18555 23715
rect 18981 23681 19015 23715
rect 34989 23681 35023 23715
rect 38301 23681 38335 23715
rect 17417 23613 17451 23647
rect 19717 23613 19751 23647
rect 7849 23477 7883 23511
rect 13001 23477 13035 23511
rect 15301 23477 15335 23511
rect 38117 23477 38151 23511
rect 19809 23273 19843 23307
rect 17969 23205 18003 23239
rect 18705 23205 18739 23239
rect 21097 23205 21131 23239
rect 19625 23137 19659 23171
rect 20729 23137 20763 23171
rect 11989 23069 12023 23103
rect 12909 23069 12943 23103
rect 13369 23069 13403 23103
rect 14565 23069 14599 23103
rect 15209 23069 15243 23103
rect 15853 23069 15887 23103
rect 16865 23069 16899 23103
rect 18889 23069 18923 23103
rect 19441 23069 19475 23103
rect 20913 23069 20947 23103
rect 17417 23001 17451 23035
rect 17509 23001 17543 23035
rect 12081 22933 12115 22967
rect 12725 22933 12759 22967
rect 13461 22933 13495 22967
rect 14381 22933 14415 22967
rect 15025 22933 15059 22967
rect 15669 22933 15703 22967
rect 16681 22933 16715 22967
rect 5457 22729 5491 22763
rect 19901 22729 19935 22763
rect 21097 22729 21131 22763
rect 14289 22661 14323 22695
rect 15669 22661 15703 22695
rect 17049 22661 17083 22695
rect 17601 22661 17635 22695
rect 1777 22593 1811 22627
rect 5641 22593 5675 22627
rect 11897 22593 11931 22627
rect 12081 22593 12115 22627
rect 13553 22593 13587 22627
rect 14197 22593 14231 22627
rect 15025 22593 15059 22627
rect 18705 22593 18739 22627
rect 19809 22593 19843 22627
rect 20453 22593 20487 22627
rect 15577 22525 15611 22559
rect 16957 22525 16991 22559
rect 19165 22525 19199 22559
rect 20637 22525 20671 22559
rect 16129 22457 16163 22491
rect 1593 22389 1627 22423
rect 12541 22389 12575 22423
rect 13645 22389 13679 22423
rect 14841 22389 14875 22423
rect 18521 22389 18555 22423
rect 13277 22185 13311 22219
rect 18613 22185 18647 22219
rect 20545 22185 20579 22219
rect 4445 22049 4479 22083
rect 12357 22049 12391 22083
rect 13093 22049 13127 22083
rect 14381 22049 14415 22083
rect 15025 22049 15059 22083
rect 16589 22049 16623 22083
rect 18245 22049 18279 22083
rect 18429 22049 18463 22083
rect 28365 22049 28399 22083
rect 4353 21981 4387 22015
rect 10057 21981 10091 22015
rect 11161 21981 11195 22015
rect 11805 21981 11839 22015
rect 12265 21981 12299 22015
rect 12909 21981 12943 22015
rect 17785 21981 17819 22015
rect 19441 21981 19475 22015
rect 20729 21981 20763 22015
rect 21373 21981 21407 22015
rect 28273 21981 28307 22015
rect 38301 21981 38335 22015
rect 14473 21913 14507 21947
rect 16129 21913 16163 21947
rect 16221 21913 16255 21947
rect 10149 21845 10183 21879
rect 10977 21845 11011 21879
rect 11621 21845 11655 21879
rect 17601 21845 17635 21879
rect 19533 21845 19567 21879
rect 21189 21845 21223 21879
rect 38117 21845 38151 21879
rect 10333 21641 10367 21675
rect 14933 21641 14967 21675
rect 20177 21641 20211 21675
rect 20637 21573 20671 21607
rect 1593 21505 1627 21539
rect 5089 21505 5123 21539
rect 8125 21505 8159 21539
rect 9689 21505 9723 21539
rect 10517 21505 10551 21539
rect 10977 21505 11011 21539
rect 11713 21505 11747 21539
rect 13185 21505 13219 21539
rect 13369 21505 13403 21539
rect 15117 21505 15151 21539
rect 15761 21505 15795 21539
rect 17325 21505 17359 21539
rect 17785 21505 17819 21539
rect 18429 21505 18463 21539
rect 19717 21505 19751 21539
rect 31401 21505 31435 21539
rect 34621 21505 34655 21539
rect 8769 21437 8803 21471
rect 11069 21437 11103 21471
rect 11897 21437 11931 21471
rect 14289 21437 14323 21471
rect 15577 21437 15611 21471
rect 18613 21437 18647 21471
rect 19533 21437 19567 21471
rect 22569 21437 22603 21471
rect 5181 21369 5215 21403
rect 13829 21369 13863 21403
rect 15945 21369 15979 21403
rect 18797 21369 18831 21403
rect 1777 21301 1811 21335
rect 8217 21301 8251 21335
rect 9781 21301 9815 21335
rect 12081 21301 12115 21335
rect 17141 21301 17175 21335
rect 17877 21301 17911 21335
rect 31493 21301 31527 21335
rect 34713 21301 34747 21335
rect 9965 21097 9999 21131
rect 15209 21097 15243 21131
rect 16129 21097 16163 21131
rect 18705 21097 18739 21131
rect 19809 21097 19843 21131
rect 28917 21097 28951 21131
rect 7757 21029 7791 21063
rect 11621 21029 11655 21063
rect 9597 20961 9631 20995
rect 9781 20961 9815 20995
rect 11437 20961 11471 20995
rect 13001 20961 13035 20995
rect 14841 20961 14875 20995
rect 16957 20961 16991 20995
rect 17693 20961 17727 20995
rect 19441 20961 19475 20995
rect 19625 20961 19659 20995
rect 22569 20961 22603 20995
rect 23213 20961 23247 20995
rect 7941 20893 7975 20927
rect 8585 20893 8619 20927
rect 11253 20893 11287 20927
rect 12909 20893 12943 20927
rect 13737 20893 13771 20927
rect 14657 20893 14691 20927
rect 15761 20893 15795 20927
rect 15945 20893 15979 20927
rect 16865 20893 16899 20927
rect 17509 20893 17543 20927
rect 18889 20893 18923 20927
rect 20545 20893 20579 20927
rect 22017 20893 22051 20927
rect 28825 20893 28859 20927
rect 18153 20825 18187 20859
rect 22661 20825 22695 20859
rect 8401 20757 8435 20791
rect 13553 20757 13587 20791
rect 20637 20757 20671 20791
rect 21833 20757 21867 20791
rect 5273 20553 5307 20587
rect 14473 20553 14507 20587
rect 18061 20553 18095 20587
rect 18797 20553 18831 20587
rect 23581 20553 23615 20587
rect 20821 20485 20855 20519
rect 24225 20485 24259 20519
rect 5457 20417 5491 20451
rect 8769 20417 8803 20451
rect 8953 20417 8987 20451
rect 10149 20417 10183 20451
rect 10333 20417 10367 20451
rect 11897 20417 11931 20451
rect 12357 20417 12391 20451
rect 13921 20417 13955 20451
rect 14381 20417 14415 20451
rect 15025 20417 15059 20451
rect 15853 20417 15887 20451
rect 17601 20417 17635 20451
rect 18981 20417 19015 20451
rect 19533 20417 19567 20451
rect 22477 20417 22511 20451
rect 23765 20417 23799 20451
rect 8125 20349 8159 20383
rect 12541 20349 12575 20383
rect 15669 20349 15703 20383
rect 17417 20349 17451 20383
rect 19717 20349 19751 20383
rect 20729 20349 20763 20383
rect 21373 20349 21407 20383
rect 22661 20349 22695 20383
rect 9137 20281 9171 20315
rect 11713 20281 11747 20315
rect 13001 20281 13035 20315
rect 15117 20281 15151 20315
rect 10609 20213 10643 20247
rect 13737 20213 13771 20247
rect 16037 20213 16071 20247
rect 20177 20213 20211 20247
rect 22845 20213 22879 20247
rect 10977 20009 11011 20043
rect 14473 20009 14507 20043
rect 16129 20009 16163 20043
rect 22201 20009 22235 20043
rect 24593 20009 24627 20043
rect 8401 19941 8435 19975
rect 9229 19941 9263 19975
rect 17693 19941 17727 19975
rect 18705 19941 18739 19975
rect 20085 19941 20119 19975
rect 23949 19941 23983 19975
rect 10057 19873 10091 19907
rect 15945 19873 15979 19907
rect 21741 19873 21775 19907
rect 23213 19873 23247 19907
rect 1777 19805 1811 19839
rect 7941 19805 7975 19839
rect 8585 19805 8619 19839
rect 9413 19805 9447 19839
rect 9873 19805 9907 19839
rect 11161 19805 11195 19839
rect 11621 19805 11655 19839
rect 12449 19805 12483 19839
rect 14657 19805 14691 19839
rect 15301 19805 15335 19839
rect 15761 19805 15795 19839
rect 18889 19805 18923 19839
rect 20821 19805 20855 19839
rect 21557 19805 21591 19839
rect 23857 19805 23891 19839
rect 24777 19805 24811 19839
rect 25421 19805 25455 19839
rect 38301 19805 38335 19839
rect 11713 19737 11747 19771
rect 12909 19737 12943 19771
rect 17141 19737 17175 19771
rect 17233 19737 17267 19771
rect 19533 19737 19567 19771
rect 19625 19737 19659 19771
rect 22753 19737 22787 19771
rect 22845 19737 22879 19771
rect 1593 19669 1627 19703
rect 7757 19669 7791 19703
rect 10517 19669 10551 19703
rect 12265 19669 12299 19703
rect 13553 19669 13587 19703
rect 15117 19669 15151 19703
rect 20637 19669 20671 19703
rect 25237 19669 25271 19703
rect 38117 19669 38151 19703
rect 7757 19465 7791 19499
rect 12725 19465 12759 19499
rect 14749 19465 14783 19499
rect 16037 19465 16071 19499
rect 16865 19465 16899 19499
rect 17509 19465 17543 19499
rect 18153 19465 18187 19499
rect 22569 19465 22603 19499
rect 24501 19465 24535 19499
rect 8677 19397 8711 19431
rect 11161 19397 11195 19431
rect 13369 19397 13403 19431
rect 20085 19397 20119 19431
rect 23397 19397 23431 19431
rect 23489 19397 23523 19431
rect 7665 19329 7699 19363
rect 8585 19329 8619 19363
rect 9229 19329 9263 19363
rect 9321 19329 9355 19363
rect 12081 19329 12115 19363
rect 14933 19329 14967 19363
rect 17049 19329 17083 19363
rect 17693 19329 17727 19363
rect 18797 19329 18831 19363
rect 19441 19329 19475 19363
rect 21097 19329 21131 19363
rect 22477 19329 22511 19363
rect 24685 19329 24719 19363
rect 9873 19261 9907 19295
rect 10517 19261 10551 19295
rect 10701 19261 10735 19295
rect 12265 19261 12299 19295
rect 13277 19261 13311 19295
rect 13921 19261 13955 19295
rect 15393 19261 15427 19295
rect 15577 19261 15611 19295
rect 18981 19261 19015 19295
rect 19993 19261 20027 19295
rect 24041 19261 24075 19295
rect 20545 19193 20579 19227
rect 21189 19125 21223 19159
rect 16773 18921 16807 18955
rect 17417 18921 17451 18955
rect 22293 18921 22327 18955
rect 10149 18853 10183 18887
rect 11805 18853 11839 18887
rect 18889 18853 18923 18887
rect 20453 18853 20487 18887
rect 8493 18785 8527 18819
rect 9689 18785 9723 18819
rect 11621 18785 11655 18819
rect 12725 18785 12759 18819
rect 13737 18785 13771 18819
rect 14289 18785 14323 18819
rect 14473 18785 14507 18819
rect 16221 18785 16255 18819
rect 18429 18785 18463 18819
rect 19901 18785 19935 18819
rect 21005 18785 21039 18819
rect 21189 18785 21223 18819
rect 23673 18785 23707 18819
rect 8401 18717 8435 18751
rect 9505 18717 9539 18751
rect 10977 18717 11011 18751
rect 11437 18717 11471 18751
rect 15669 18717 15703 18751
rect 16129 18717 16163 18751
rect 16957 18717 16991 18751
rect 17601 18717 17635 18751
rect 18245 18717 18279 18751
rect 22477 18717 22511 18751
rect 33057 18717 33091 18751
rect 38301 18717 38335 18751
rect 12817 18649 12851 18683
rect 19993 18649 20027 18683
rect 23029 18649 23063 18683
rect 23121 18649 23155 18683
rect 7205 18581 7239 18615
rect 10793 18581 10827 18615
rect 14933 18581 14967 18615
rect 15485 18581 15519 18615
rect 21649 18581 21683 18615
rect 33149 18581 33183 18615
rect 38117 18581 38151 18615
rect 9045 18377 9079 18411
rect 9689 18377 9723 18411
rect 14197 18377 14231 18411
rect 18337 18377 18371 18411
rect 21189 18377 21223 18411
rect 23673 18377 23707 18411
rect 7113 18309 7147 18343
rect 7205 18309 7239 18343
rect 7757 18309 7791 18343
rect 11897 18309 11931 18343
rect 15669 18309 15703 18343
rect 17049 18309 17083 18343
rect 1777 18241 1811 18275
rect 8585 18241 8619 18275
rect 9229 18241 9263 18275
rect 10517 18241 10551 18275
rect 11161 18241 11195 18275
rect 11805 18241 11839 18275
rect 12633 18241 12667 18275
rect 14381 18241 14415 18275
rect 15025 18241 15059 18275
rect 18245 18241 18279 18275
rect 18889 18241 18923 18275
rect 22477 18241 22511 18275
rect 23581 18241 23615 18275
rect 24409 18241 24443 18275
rect 13093 18173 13127 18207
rect 13277 18173 13311 18207
rect 15577 18173 15611 18207
rect 16957 18173 16991 18207
rect 17417 18173 17451 18207
rect 19073 18173 19107 18207
rect 20545 18173 20579 18207
rect 20729 18173 20763 18207
rect 22661 18173 22695 18207
rect 10977 18105 11011 18139
rect 12449 18105 12483 18139
rect 16129 18105 16163 18139
rect 1593 18037 1627 18071
rect 8401 18037 8435 18071
rect 10333 18037 10367 18071
rect 13737 18037 13771 18071
rect 14841 18037 14875 18071
rect 19533 18037 19567 18071
rect 22845 18037 22879 18071
rect 24225 18037 24259 18071
rect 7113 17833 7147 17867
rect 9505 17833 9539 17867
rect 13737 17833 13771 17867
rect 16957 17833 16991 17867
rect 18705 17833 18739 17867
rect 20913 17833 20947 17867
rect 21557 17833 21591 17867
rect 23397 17833 23431 17867
rect 11897 17765 11931 17799
rect 14657 17765 14691 17799
rect 22753 17765 22787 17799
rect 10885 17697 10919 17731
rect 13093 17697 13127 17731
rect 15393 17697 15427 17731
rect 16037 17697 16071 17731
rect 17601 17697 17635 17731
rect 19809 17697 19843 17731
rect 20453 17697 20487 17731
rect 22201 17697 22235 17731
rect 22385 17697 22419 17731
rect 1961 17629 1995 17663
rect 2421 17629 2455 17663
rect 3249 17629 3283 17663
rect 5181 17629 5215 17663
rect 6653 17629 6687 17663
rect 7297 17629 7331 17663
rect 7757 17629 7791 17663
rect 8585 17629 8619 17663
rect 9689 17629 9723 17663
rect 11805 17629 11839 17663
rect 12633 17629 12667 17663
rect 13277 17629 13311 17663
rect 14841 17629 14875 17663
rect 16497 17629 16531 17663
rect 16681 17629 16715 17663
rect 17785 17629 17819 17663
rect 18889 17629 18923 17663
rect 21097 17629 21131 17663
rect 21741 17629 21775 17663
rect 23305 17629 23339 17663
rect 31493 17629 31527 17663
rect 33149 17629 33183 17663
rect 10241 17561 10275 17595
rect 10333 17561 10367 17595
rect 15485 17561 15519 17595
rect 19901 17561 19935 17595
rect 1777 17493 1811 17527
rect 2513 17493 2547 17527
rect 3065 17493 3099 17527
rect 4997 17493 5031 17527
rect 6469 17493 6503 17527
rect 7849 17493 7883 17527
rect 8401 17493 8435 17527
rect 12449 17493 12483 17527
rect 18245 17493 18279 17527
rect 31585 17493 31619 17527
rect 33241 17493 33275 17527
rect 8585 17289 8619 17323
rect 10333 17289 10367 17323
rect 11069 17289 11103 17323
rect 12909 17289 12943 17323
rect 13553 17289 13587 17323
rect 17509 17289 17543 17323
rect 19993 17289 20027 17323
rect 21005 17289 21039 17323
rect 22661 17289 22695 17323
rect 23121 17289 23155 17323
rect 4721 17221 4755 17255
rect 14841 17221 14875 17255
rect 15485 17221 15519 17255
rect 18889 17221 18923 17255
rect 1869 17153 1903 17187
rect 2605 17153 2639 17187
rect 3249 17153 3283 17187
rect 5825 17153 5859 17187
rect 8769 17153 8803 17187
rect 9413 17153 9447 17187
rect 10977 17153 11011 17187
rect 12449 17153 12483 17187
rect 13093 17153 13127 17187
rect 16313 17153 16347 17187
rect 16865 17153 16899 17187
rect 18245 17153 18279 17187
rect 21189 17153 21223 17187
rect 23305 17153 23339 17187
rect 23949 17153 23983 17187
rect 24593 17153 24627 17187
rect 38025 17153 38059 17187
rect 4629 17085 4663 17119
rect 4905 17085 4939 17119
rect 6745 17085 6779 17119
rect 7389 17085 7423 17119
rect 7573 17085 7607 17119
rect 9229 17085 9263 17119
rect 14197 17085 14231 17119
rect 14381 17085 14415 17119
rect 17049 17085 17083 17119
rect 18429 17085 18463 17119
rect 19349 17085 19383 17119
rect 19533 17085 19567 17119
rect 22017 17085 22051 17119
rect 22201 17085 22235 17119
rect 3341 17017 3375 17051
rect 24409 17017 24443 17051
rect 38209 17017 38243 17051
rect 1961 16949 1995 16983
rect 2697 16949 2731 16983
rect 5917 16949 5951 16983
rect 7757 16949 7791 16983
rect 9689 16949 9723 16983
rect 12265 16949 12299 16983
rect 16129 16949 16163 16983
rect 23765 16949 23799 16983
rect 11621 16745 11655 16779
rect 12909 16745 12943 16779
rect 16773 16745 16807 16779
rect 22845 16745 22879 16779
rect 8493 16677 8527 16711
rect 10977 16677 11011 16711
rect 16037 16677 16071 16711
rect 20085 16677 20119 16711
rect 23489 16677 23523 16711
rect 4721 16609 4755 16643
rect 6285 16609 6319 16643
rect 6469 16609 6503 16643
rect 7941 16609 7975 16643
rect 9321 16609 9355 16643
rect 15485 16609 15519 16643
rect 19533 16609 19567 16643
rect 20637 16609 20671 16643
rect 20821 16609 20855 16643
rect 21741 16609 21775 16643
rect 1593 16541 1627 16575
rect 2329 16541 2363 16575
rect 2973 16541 3007 16575
rect 3985 16541 4019 16575
rect 5641 16541 5675 16575
rect 9137 16541 9171 16575
rect 10517 16541 10551 16575
rect 11161 16541 11195 16575
rect 11805 16541 11839 16575
rect 12449 16541 12483 16575
rect 13093 16541 13127 16575
rect 13737 16541 13771 16575
rect 14933 16541 14967 16575
rect 16957 16541 16991 16575
rect 17601 16541 17635 16575
rect 18245 16541 18279 16575
rect 18705 16541 18739 16575
rect 21925 16541 21959 16575
rect 23029 16541 23063 16575
rect 23673 16541 23707 16575
rect 3065 16473 3099 16507
rect 8033 16473 8067 16507
rect 15577 16473 15611 16507
rect 19625 16473 19659 16507
rect 1777 16405 1811 16439
rect 2421 16405 2455 16439
rect 4077 16405 4111 16439
rect 5733 16405 5767 16439
rect 6929 16405 6963 16439
rect 9781 16405 9815 16439
rect 10333 16405 10367 16439
rect 12265 16405 12299 16439
rect 13553 16405 13587 16439
rect 14749 16405 14783 16439
rect 17417 16405 17451 16439
rect 18061 16405 18095 16439
rect 21281 16405 21315 16439
rect 22385 16405 22419 16439
rect 5365 16201 5399 16235
rect 9689 16201 9723 16235
rect 12725 16201 12759 16235
rect 21189 16201 21223 16235
rect 22753 16201 22787 16235
rect 23213 16201 23247 16235
rect 7757 16133 7791 16167
rect 8493 16133 8527 16167
rect 10609 16133 10643 16167
rect 11161 16133 11195 16167
rect 14933 16133 14967 16167
rect 18705 16133 18739 16167
rect 19625 16133 19659 16167
rect 1961 16065 1995 16099
rect 2513 16065 2547 16099
rect 3157 16065 3191 16099
rect 4445 16065 4479 16099
rect 5549 16065 5583 16099
rect 7205 16065 7239 16099
rect 7665 16065 7699 16099
rect 9873 16065 9907 16099
rect 12357 16065 12391 16099
rect 12633 16065 12667 16099
rect 13645 16065 13679 16099
rect 14841 16065 14875 16099
rect 15669 16065 15703 16099
rect 16129 16065 16163 16099
rect 23397 16065 23431 16099
rect 23857 16065 23891 16099
rect 34161 16065 34195 16099
rect 3801 15997 3835 16031
rect 8401 15997 8435 16031
rect 8677 15997 8711 16031
rect 10517 15997 10551 16031
rect 13185 15997 13219 16031
rect 13461 15997 13495 16031
rect 16865 15997 16899 16031
rect 17049 15997 17083 16031
rect 18613 15997 18647 16031
rect 20085 15997 20119 16031
rect 20269 15997 20303 16031
rect 22109 15997 22143 16031
rect 22293 15997 22327 16031
rect 23949 15997 23983 16031
rect 15485 15929 15519 15963
rect 34253 15929 34287 15963
rect 1777 15861 1811 15895
rect 2605 15861 2639 15895
rect 3249 15861 3283 15895
rect 4537 15861 4571 15895
rect 7021 15861 7055 15895
rect 12173 15861 12207 15895
rect 13829 15861 13863 15895
rect 17233 15861 17267 15895
rect 20453 15861 20487 15895
rect 7205 15657 7239 15691
rect 9321 15657 9355 15691
rect 11069 15657 11103 15691
rect 12633 15657 12667 15691
rect 14565 15657 14599 15691
rect 17141 15657 17175 15691
rect 22845 15657 22879 15691
rect 35081 15657 35115 15691
rect 38117 15657 38151 15691
rect 1593 15589 1627 15623
rect 8493 15589 8527 15623
rect 21465 15589 21499 15623
rect 7941 15521 7975 15555
rect 9965 15521 9999 15555
rect 12173 15521 12207 15555
rect 13277 15521 13311 15555
rect 15301 15521 15335 15555
rect 18337 15521 18371 15555
rect 19533 15521 19567 15555
rect 21097 15521 21131 15555
rect 22201 15521 22235 15555
rect 1777 15453 1811 15487
rect 2421 15453 2455 15487
rect 3249 15453 3283 15487
rect 4537 15453 4571 15487
rect 5365 15453 5399 15487
rect 6193 15453 6227 15487
rect 7389 15453 7423 15487
rect 9229 15453 9263 15487
rect 9873 15453 9907 15487
rect 10517 15453 10551 15487
rect 10701 15453 10735 15487
rect 11989 15453 12023 15487
rect 13093 15453 13127 15487
rect 14473 15453 14507 15487
rect 15117 15453 15151 15487
rect 16497 15453 16531 15487
rect 16681 15453 16715 15487
rect 18153 15453 18187 15487
rect 21281 15453 21315 15487
rect 23029 15453 23063 15487
rect 23673 15453 23707 15487
rect 35265 15453 35299 15487
rect 38301 15453 38335 15487
rect 8033 15385 8067 15419
rect 19625 15385 19659 15419
rect 20545 15385 20579 15419
rect 2513 15317 2547 15351
rect 3065 15317 3099 15351
rect 4629 15317 4663 15351
rect 5181 15317 5215 15351
rect 6285 15317 6319 15351
rect 13737 15317 13771 15351
rect 15761 15317 15795 15351
rect 18797 15317 18831 15351
rect 23489 15317 23523 15351
rect 3157 15113 3191 15147
rect 5089 15113 5123 15147
rect 7205 15113 7239 15147
rect 7849 15113 7883 15147
rect 8585 15113 8619 15147
rect 13369 15113 13403 15147
rect 16221 15113 16255 15147
rect 20177 15113 20211 15147
rect 21281 15113 21315 15147
rect 23121 15113 23155 15147
rect 14105 15045 14139 15079
rect 17302 15045 17336 15079
rect 1869 14977 1903 15011
rect 2697 14977 2731 15011
rect 3341 14977 3375 15011
rect 3985 14977 4019 15011
rect 4629 14977 4663 15011
rect 5273 14977 5307 15011
rect 5733 14977 5767 15011
rect 6745 14977 6779 15011
rect 7389 14977 7423 15011
rect 8033 14977 8067 15011
rect 8493 14977 8527 15011
rect 9229 14977 9263 15011
rect 10517 14977 10551 15011
rect 11161 14977 11195 15011
rect 12817 14977 12851 15011
rect 13277 14977 13311 15011
rect 15669 14977 15703 15011
rect 16129 14977 16163 15011
rect 18613 14977 18647 15011
rect 21189 14977 21223 15011
rect 22017 14977 22051 15011
rect 23305 14977 23339 15011
rect 9413 14909 9447 14943
rect 10701 14909 10735 14943
rect 12173 14909 12207 14943
rect 12326 14909 12360 14943
rect 14013 14909 14047 14943
rect 17234 14909 17268 14943
rect 18429 14909 18463 14943
rect 19533 14909 19567 14943
rect 19717 14909 19751 14943
rect 22201 14909 22235 14943
rect 14565 14841 14599 14875
rect 17785 14841 17819 14875
rect 19073 14841 19107 14875
rect 22385 14841 22419 14875
rect 1961 14773 1995 14807
rect 2513 14773 2547 14807
rect 3801 14773 3835 14807
rect 4445 14773 4479 14807
rect 5825 14773 5859 14807
rect 6561 14773 6595 14807
rect 9597 14773 9631 14807
rect 15485 14773 15519 14807
rect 2605 14569 2639 14603
rect 10333 14569 10367 14603
rect 11069 14569 11103 14603
rect 11713 14569 11747 14603
rect 12265 14569 12299 14603
rect 12909 14569 12943 14603
rect 15025 14569 15059 14603
rect 17693 14569 17727 14603
rect 20821 14569 20855 14603
rect 22661 14569 22695 14603
rect 28457 14569 28491 14603
rect 3985 14433 4019 14467
rect 4169 14433 4203 14467
rect 5549 14433 5583 14467
rect 8585 14433 8619 14467
rect 15577 14433 15611 14467
rect 16957 14433 16991 14467
rect 18429 14433 18463 14467
rect 19625 14433 19659 14467
rect 20085 14433 20119 14467
rect 21465 14433 21499 14467
rect 1593 14365 1627 14399
rect 2513 14365 2547 14399
rect 3433 14365 3467 14399
rect 6837 14365 6871 14399
rect 7297 14365 7331 14399
rect 7941 14365 7975 14399
rect 8125 14365 8159 14399
rect 9873 14365 9907 14399
rect 10517 14365 10551 14399
rect 10977 14365 11011 14399
rect 11621 14365 11655 14399
rect 12449 14365 12483 14399
rect 13093 14365 13127 14399
rect 13553 14365 13587 14399
rect 14473 14365 14507 14399
rect 14933 14365 14967 14399
rect 17601 14365 17635 14399
rect 18245 14365 18279 14399
rect 20729 14365 20763 14399
rect 21649 14365 21683 14399
rect 22569 14365 22603 14399
rect 23213 14365 23247 14399
rect 28365 14365 28399 14399
rect 4629 14297 4663 14331
rect 5273 14297 5307 14331
rect 5365 14297 5399 14331
rect 16314 14297 16348 14331
rect 16405 14297 16439 14331
rect 19717 14297 19751 14331
rect 1777 14229 1811 14263
rect 3249 14229 3283 14263
rect 6653 14229 6687 14263
rect 7389 14229 7423 14263
rect 9689 14229 9723 14263
rect 13645 14229 13679 14263
rect 14289 14229 14323 14263
rect 18889 14229 18923 14263
rect 22109 14229 22143 14263
rect 23305 14229 23339 14263
rect 4997 14025 5031 14059
rect 6837 14025 6871 14059
rect 8125 14025 8159 14059
rect 9137 14025 9171 14059
rect 9781 14025 9815 14059
rect 18889 14025 18923 14059
rect 19809 14025 19843 14059
rect 1869 13957 1903 13991
rect 17049 13957 17083 13991
rect 17601 13957 17635 13991
rect 21465 13957 21499 13991
rect 23765 13957 23799 13991
rect 4077 13889 4111 13923
rect 5181 13889 5215 13923
rect 5825 13889 5859 13923
rect 7021 13889 7055 13923
rect 7665 13889 7699 13923
rect 9045 13889 9079 13923
rect 9689 13889 9723 13923
rect 10517 13889 10551 13923
rect 10977 13889 11011 13923
rect 12265 13889 12299 13923
rect 15669 13889 15703 13923
rect 16313 13889 16347 13923
rect 18245 13889 18279 13923
rect 19993 13889 20027 13923
rect 21005 13889 21039 13923
rect 23121 13889 23155 13923
rect 24409 13889 24443 13923
rect 38025 13889 38059 13923
rect 1593 13821 1627 13855
rect 3893 13821 3927 13855
rect 5917 13821 5951 13855
rect 12725 13821 12759 13855
rect 12909 13821 12943 13855
rect 13369 13821 13403 13855
rect 14013 13821 14047 13855
rect 14197 13821 14231 13855
rect 14657 13821 14691 13855
rect 16957 13821 16991 13855
rect 18429 13821 18463 13855
rect 20821 13821 20855 13855
rect 22017 13821 22051 13855
rect 22201 13821 22235 13855
rect 23305 13821 23339 13855
rect 12081 13753 12115 13787
rect 15485 13753 15519 13787
rect 16129 13753 16163 13787
rect 22385 13753 22419 13787
rect 24225 13753 24259 13787
rect 3341 13685 3375 13719
rect 4537 13685 4571 13719
rect 7481 13685 7515 13719
rect 10333 13685 10367 13719
rect 11069 13685 11103 13719
rect 38209 13685 38243 13719
rect 4353 13481 4387 13515
rect 8033 13481 8067 13515
rect 10701 13481 10735 13515
rect 14381 13481 14415 13515
rect 16037 13481 16071 13515
rect 17693 13481 17727 13515
rect 18613 13481 18647 13515
rect 20637 13481 20671 13515
rect 21833 13481 21867 13515
rect 23581 13481 23615 13515
rect 33425 13481 33459 13515
rect 11253 13413 11287 13447
rect 20085 13413 20119 13447
rect 1593 13345 1627 13379
rect 6745 13345 6779 13379
rect 12081 13345 12115 13379
rect 17049 13345 17083 13379
rect 19533 13345 19567 13379
rect 22477 13345 22511 13379
rect 23121 13345 23155 13379
rect 4537 13277 4571 13311
rect 4997 13277 5031 13311
rect 7389 13277 7423 13311
rect 8217 13277 8251 13311
rect 9505 13277 9539 13311
rect 10149 13277 10183 13311
rect 10609 13277 10643 13311
rect 11437 13277 11471 13311
rect 11897 13277 11931 13311
rect 13737 13277 13771 13311
rect 14565 13277 14599 13311
rect 15209 13277 15243 13311
rect 15669 13277 15703 13311
rect 15853 13277 15887 13311
rect 17233 13277 17267 13311
rect 18245 13277 18279 13311
rect 18429 13277 18463 13311
rect 20821 13277 20855 13311
rect 21741 13277 21775 13311
rect 23765 13277 23799 13311
rect 33333 13277 33367 13311
rect 1869 13209 1903 13243
rect 5273 13209 5307 13243
rect 7481 13209 7515 13243
rect 19625 13209 19659 13243
rect 22569 13209 22603 13243
rect 3341 13141 3375 13175
rect 9321 13141 9355 13175
rect 9965 13141 9999 13175
rect 12541 13141 12575 13175
rect 13553 13141 13587 13175
rect 15025 13141 15059 13175
rect 3433 12937 3467 12971
rect 10977 12937 11011 12971
rect 11805 12937 11839 12971
rect 15025 12937 15059 12971
rect 16221 12937 16255 12971
rect 18153 12937 18187 12971
rect 19441 12937 19475 12971
rect 19901 12937 19935 12971
rect 21281 12937 21315 12971
rect 22017 12937 22051 12971
rect 4169 12869 4203 12903
rect 8125 12869 8159 12903
rect 12633 12869 12667 12903
rect 23213 12869 23247 12903
rect 1685 12801 1719 12835
rect 3893 12801 3927 12835
rect 6561 12801 6595 12835
rect 8033 12801 8067 12835
rect 8861 12801 8895 12835
rect 10517 12801 10551 12835
rect 11161 12801 11195 12835
rect 11989 12801 12023 12835
rect 13921 12801 13955 12835
rect 14565 12801 14599 12835
rect 15761 12801 15795 12835
rect 18061 12801 18095 12835
rect 20085 12801 20119 12835
rect 20729 12801 20763 12835
rect 21465 12801 21499 12835
rect 22201 12801 22235 12835
rect 24409 12801 24443 12835
rect 31401 12801 31435 12835
rect 1961 12733 1995 12767
rect 6745 12733 6779 12767
rect 8677 12733 8711 12767
rect 12541 12733 12575 12767
rect 13185 12733 13219 12767
rect 14381 12733 14415 12767
rect 15577 12733 15611 12767
rect 16865 12733 16899 12767
rect 17049 12733 17083 12767
rect 18797 12733 18831 12767
rect 18981 12733 19015 12767
rect 23121 12733 23155 12767
rect 23765 12733 23799 12767
rect 13737 12665 13771 12699
rect 31493 12665 31527 12699
rect 5641 12597 5675 12631
rect 6929 12597 6963 12631
rect 9321 12597 9355 12631
rect 10333 12597 10367 12631
rect 17233 12597 17267 12631
rect 20545 12597 20579 12631
rect 24225 12597 24259 12631
rect 9873 12393 9907 12427
rect 10793 12393 10827 12427
rect 17693 12393 17727 12427
rect 19625 12393 19659 12427
rect 11805 12325 11839 12359
rect 24961 12325 24995 12359
rect 4537 12257 4571 12291
rect 5457 12257 5491 12291
rect 7849 12257 7883 12291
rect 9229 12257 9263 12291
rect 11437 12257 11471 12291
rect 12633 12257 12667 12291
rect 14473 12257 14507 12291
rect 15117 12257 15151 12291
rect 16313 12257 16347 12291
rect 16589 12257 16623 12291
rect 18337 12257 18371 12291
rect 20453 12257 20487 12291
rect 23397 12257 23431 12291
rect 24041 12257 24075 12291
rect 1685 12189 1719 12223
rect 4353 12189 4387 12223
rect 7665 12189 7699 12223
rect 9413 12189 9447 12223
rect 10977 12189 11011 12223
rect 11621 12189 11655 12223
rect 15301 12189 15335 12223
rect 17877 12189 17911 12223
rect 19809 12189 19843 12223
rect 20637 12189 20671 12223
rect 21557 12189 21591 12223
rect 22385 12189 22419 12223
rect 24593 12189 24627 12223
rect 24777 12189 24811 12223
rect 35449 12189 35483 12223
rect 1961 12121 1995 12155
rect 4997 12121 5031 12155
rect 5733 12121 5767 12155
rect 12725 12121 12759 12155
rect 13277 12121 13311 12155
rect 16405 12121 16439 12155
rect 21649 12121 21683 12155
rect 23489 12121 23523 12155
rect 3433 12053 3467 12087
rect 7205 12053 7239 12087
rect 8309 12053 8343 12087
rect 15761 12053 15795 12087
rect 21097 12053 21131 12087
rect 22201 12053 22235 12087
rect 35541 12053 35575 12087
rect 5273 11849 5307 11883
rect 5917 11849 5951 11883
rect 12725 11849 12759 11883
rect 14289 11849 14323 11883
rect 14933 11849 14967 11883
rect 17049 11849 17083 11883
rect 17601 11849 17635 11883
rect 18337 11849 18371 11883
rect 21097 11849 21131 11883
rect 22109 11849 22143 11883
rect 22753 11849 22787 11883
rect 24685 11849 24719 11883
rect 34253 11849 34287 11883
rect 38117 11849 38151 11883
rect 1869 11781 1903 11815
rect 7205 11781 7239 11815
rect 11161 11781 11195 11815
rect 23673 11781 23707 11815
rect 1777 11713 1811 11747
rect 4629 11713 4663 11747
rect 5825 11713 5859 11747
rect 6561 11713 6595 11747
rect 6745 11713 6779 11747
rect 7665 11713 7699 11747
rect 10517 11713 10551 11747
rect 12081 11713 12115 11747
rect 13185 11713 13219 11747
rect 14473 11713 14507 11747
rect 15117 11713 15151 11747
rect 16957 11713 16991 11747
rect 17785 11713 17819 11747
rect 18245 11713 18279 11747
rect 18889 11713 18923 11747
rect 19993 11713 20027 11747
rect 21281 11713 21315 11747
rect 22017 11713 22051 11747
rect 22661 11713 22695 11747
rect 24869 11713 24903 11747
rect 34437 11713 34471 11747
rect 38301 11713 38335 11747
rect 2329 11645 2363 11679
rect 2605 11645 2639 11679
rect 4077 11645 4111 11679
rect 4813 11645 4847 11679
rect 8309 11645 8343 11679
rect 8585 11645 8619 11679
rect 10701 11645 10735 11679
rect 12265 11645 12299 11679
rect 13369 11645 13403 11679
rect 15577 11645 15611 11679
rect 15761 11645 15795 11679
rect 19073 11645 19107 11679
rect 20177 11645 20211 11679
rect 23581 11645 23615 11679
rect 25329 11645 25363 11679
rect 16221 11577 16255 11611
rect 24133 11577 24167 11611
rect 7757 11509 7791 11543
rect 10057 11509 10091 11543
rect 13829 11509 13863 11543
rect 19533 11509 19567 11543
rect 20637 11509 20671 11543
rect 9505 11305 9539 11339
rect 15853 11305 15887 11339
rect 18429 11305 18463 11339
rect 19533 11305 19567 11339
rect 22661 11305 22695 11339
rect 24593 11305 24627 11339
rect 3433 11237 3467 11271
rect 5917 11237 5951 11271
rect 13737 11237 13771 11271
rect 1961 11169 1995 11203
rect 4169 11169 4203 11203
rect 6837 11169 6871 11203
rect 7113 11169 7147 11203
rect 8585 11169 8619 11203
rect 10149 11169 10183 11203
rect 14933 11169 14967 11203
rect 20177 11169 20211 11203
rect 21281 11169 21315 11203
rect 23305 11169 23339 11203
rect 1685 11101 1719 11135
rect 9689 11101 9723 11135
rect 12541 11101 12575 11135
rect 12633 11101 12667 11135
rect 13093 11101 13127 11135
rect 13277 11101 13311 11135
rect 14841 11101 14875 11135
rect 16037 11101 16071 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 17693 11101 17727 11135
rect 18613 11101 18647 11135
rect 19441 11101 19475 11135
rect 20361 11101 20395 11135
rect 22845 11101 22879 11135
rect 24777 11101 24811 11135
rect 29745 11101 29779 11135
rect 4445 11033 4479 11067
rect 10425 11033 10459 11067
rect 17785 11033 17819 11067
rect 29837 11033 29871 11067
rect 4077 10965 4111 10999
rect 11897 10965 11931 10999
rect 17141 10965 17175 10999
rect 20821 10965 20855 10999
rect 1685 10761 1719 10795
rect 2329 10761 2363 10795
rect 5825 10761 5859 10795
rect 8493 10761 8527 10795
rect 15577 10761 15611 10795
rect 16221 10761 16255 10795
rect 18889 10761 18923 10795
rect 19441 10761 19475 10795
rect 20269 10761 20303 10795
rect 20821 10761 20855 10795
rect 23397 10761 23431 10795
rect 24041 10761 24075 10795
rect 27261 10761 27295 10795
rect 7021 10693 7055 10727
rect 1593 10625 1627 10659
rect 2237 10625 2271 10659
rect 5181 10625 5215 10659
rect 6009 10625 6043 10659
rect 6745 10625 6779 10659
rect 14381 10625 14415 10659
rect 14841 10625 14875 10659
rect 15485 10625 15519 10659
rect 16129 10625 16163 10659
rect 20177 10625 20211 10659
rect 21005 10625 21039 10659
rect 22661 10625 22695 10659
rect 23581 10625 23615 10659
rect 24225 10625 24259 10659
rect 27169 10625 27203 10659
rect 35081 10625 35115 10659
rect 36461 10625 36495 10659
rect 38025 10625 38059 10659
rect 2881 10557 2915 10591
rect 3157 10557 3191 10591
rect 5273 10557 5307 10591
rect 9413 10557 9447 10591
rect 11713 10557 11747 10591
rect 11989 10557 12023 10591
rect 16865 10557 16899 10591
rect 17049 10557 17083 10591
rect 18245 10557 18279 10591
rect 18429 10557 18463 10591
rect 11161 10489 11195 10523
rect 14933 10489 14967 10523
rect 17233 10489 17267 10523
rect 22753 10489 22787 10523
rect 34897 10489 34931 10523
rect 4629 10421 4663 10455
rect 9670 10421 9704 10455
rect 13461 10421 13495 10455
rect 14197 10421 14231 10455
rect 36277 10421 36311 10455
rect 38209 10421 38243 10455
rect 4629 10217 4663 10251
rect 7665 10217 7699 10251
rect 13553 10217 13587 10251
rect 14657 10217 14691 10251
rect 15669 10217 15703 10251
rect 18613 10217 18647 10251
rect 20177 10217 20211 10251
rect 23489 10217 23523 10251
rect 8493 10149 8527 10183
rect 11897 10149 11931 10183
rect 17601 10149 17635 10183
rect 19625 10149 19659 10183
rect 1961 10081 1995 10115
rect 3985 10081 4019 10115
rect 4169 10081 4203 10115
rect 5917 10081 5951 10115
rect 10149 10081 10183 10115
rect 12541 10081 12575 10115
rect 16313 10081 16347 10115
rect 17049 10081 17083 10115
rect 33977 10081 34011 10115
rect 1685 10013 1719 10047
rect 5457 10013 5491 10047
rect 8401 10013 8435 10047
rect 9689 10013 9723 10047
rect 12357 10013 12391 10047
rect 13461 10013 13495 10047
rect 14289 10013 14323 10047
rect 14473 10013 14507 10047
rect 15853 10013 15887 10047
rect 18521 10013 18555 10047
rect 19533 10013 19567 10047
rect 20361 10013 20395 10047
rect 23121 10013 23155 10047
rect 23305 10013 23339 10047
rect 33885 10013 33919 10047
rect 6193 9945 6227 9979
rect 10425 9945 10459 9979
rect 17141 9945 17175 9979
rect 3433 9877 3467 9911
rect 5273 9877 5307 9911
rect 9505 9877 9539 9911
rect 13001 9877 13035 9911
rect 23305 9673 23339 9707
rect 4353 9605 4387 9639
rect 6929 9605 6963 9639
rect 9321 9605 9355 9639
rect 12265 9605 12299 9639
rect 15761 9605 15795 9639
rect 17049 9605 17083 9639
rect 6653 9537 6687 9571
rect 12173 9537 12207 9571
rect 13001 9537 13035 9571
rect 13461 9537 13495 9571
rect 14289 9537 14323 9571
rect 15117 9537 15151 9571
rect 18337 9537 18371 9571
rect 23213 9537 23247 9571
rect 1593 9469 1627 9503
rect 1869 9469 1903 9503
rect 3617 9469 3651 9503
rect 4077 9469 4111 9503
rect 8401 9469 8435 9503
rect 9045 9469 9079 9503
rect 15669 9469 15703 9503
rect 16957 9469 16991 9503
rect 14105 9401 14139 9435
rect 16221 9401 16255 9435
rect 17509 9401 17543 9435
rect 5825 9333 5859 9367
rect 10793 9333 10827 9367
rect 12817 9333 12851 9367
rect 13553 9333 13587 9367
rect 14933 9333 14967 9367
rect 18429 9333 18463 9367
rect 5733 9129 5767 9163
rect 9413 9129 9447 9163
rect 12449 9129 12483 9163
rect 16681 9129 16715 9163
rect 18061 9129 18095 9163
rect 3341 9061 3375 9095
rect 11805 9061 11839 9095
rect 14841 9061 14875 9095
rect 22385 9061 22419 9095
rect 3985 8993 4019 9027
rect 4261 8993 4295 9027
rect 10333 8993 10367 9027
rect 13093 8993 13127 9027
rect 13277 8993 13311 9027
rect 16037 8993 16071 9027
rect 16221 8993 16255 9027
rect 21833 8993 21867 9027
rect 24961 8993 24995 9027
rect 1593 8925 1627 8959
rect 6837 8925 6871 8959
rect 9597 8925 9631 8959
rect 10057 8925 10091 8959
rect 12633 8925 12667 8959
rect 14749 8925 14783 8959
rect 15393 8925 15427 8959
rect 18245 8925 18279 8959
rect 21097 8925 21131 8959
rect 24869 8925 24903 8959
rect 38025 8925 38059 8959
rect 1869 8857 1903 8891
rect 7113 8857 7147 8891
rect 21189 8857 21223 8891
rect 21925 8857 21959 8891
rect 8585 8789 8619 8823
rect 13737 8789 13771 8823
rect 15485 8789 15519 8823
rect 17417 8789 17451 8823
rect 38209 8789 38243 8823
rect 8769 8585 8803 8619
rect 10977 8585 11011 8619
rect 15025 8585 15059 8619
rect 2237 8517 2271 8551
rect 5273 8517 5307 8551
rect 15770 8517 15804 8551
rect 17325 8517 17359 8551
rect 17417 8517 17451 8551
rect 18521 8517 18555 8551
rect 4445 8449 4479 8483
rect 5181 8449 5215 8483
rect 6009 8449 6043 8483
rect 9229 8449 9263 8483
rect 14473 8449 14507 8483
rect 14933 8449 14967 8483
rect 18429 8449 18463 8483
rect 20085 8449 20119 8483
rect 20545 8449 20579 8483
rect 28273 8449 28307 8483
rect 1961 8381 1995 8415
rect 3985 8381 4019 8415
rect 7021 8381 7055 8415
rect 7297 8381 7331 8415
rect 11713 8381 11747 8415
rect 11989 8381 12023 8415
rect 13461 8381 13495 8415
rect 15669 8381 15703 8415
rect 15945 8381 15979 8415
rect 17601 8381 17635 8415
rect 20729 8381 20763 8415
rect 5825 8313 5859 8347
rect 14289 8313 14323 8347
rect 21189 8313 21223 8347
rect 28365 8313 28399 8347
rect 4629 8245 4663 8279
rect 9486 8245 9520 8279
rect 19901 8245 19935 8279
rect 4629 8041 4663 8075
rect 12449 8041 12483 8075
rect 15669 8041 15703 8075
rect 17417 8041 17451 8075
rect 20453 8041 20487 8075
rect 4077 7973 4111 8007
rect 7297 7973 7331 8007
rect 9505 7973 9539 8007
rect 27813 7973 27847 8007
rect 1869 7905 1903 7939
rect 10057 7905 10091 7939
rect 14473 7905 14507 7939
rect 16313 7905 16347 7939
rect 1593 7837 1627 7871
rect 3985 7837 4019 7871
rect 4813 7837 4847 7871
rect 5549 7837 5583 7871
rect 8401 7837 8435 7871
rect 9413 7837 9447 7871
rect 12357 7837 12391 7871
rect 13093 7837 13127 7871
rect 13277 7837 13311 7871
rect 14289 7837 14323 7871
rect 15853 7837 15887 7871
rect 16497 7837 16531 7871
rect 17601 7837 17635 7871
rect 18245 7837 18279 7871
rect 18705 7837 18739 7871
rect 20637 7837 20671 7871
rect 21925 7837 21959 7871
rect 22753 7837 22787 7871
rect 27721 7837 27755 7871
rect 5825 7769 5859 7803
rect 8493 7769 8527 7803
rect 10333 7769 10367 7803
rect 3341 7701 3375 7735
rect 11805 7701 11839 7735
rect 13737 7701 13771 7735
rect 14933 7701 14967 7735
rect 16957 7701 16991 7735
rect 18061 7701 18095 7735
rect 18797 7701 18831 7735
rect 22017 7701 22051 7735
rect 22569 7701 22603 7735
rect 23213 7701 23247 7735
rect 6653 7497 6687 7531
rect 11161 7497 11195 7531
rect 16037 7497 16071 7531
rect 16957 7497 16991 7531
rect 17509 7497 17543 7531
rect 18245 7497 18279 7531
rect 18889 7497 18923 7531
rect 29561 7497 29595 7531
rect 33885 7497 33919 7531
rect 38117 7497 38151 7531
rect 1869 7429 1903 7463
rect 6009 7429 6043 7463
rect 8217 7429 8251 7463
rect 11989 7429 12023 7463
rect 14105 7429 14139 7463
rect 22201 7429 22235 7463
rect 23305 7429 23339 7463
rect 23397 7429 23431 7463
rect 6561 7361 6595 7395
rect 7481 7361 7515 7395
rect 9965 7361 9999 7395
rect 11713 7361 11747 7395
rect 14657 7361 14691 7395
rect 15301 7361 15335 7395
rect 16221 7361 16255 7395
rect 16865 7361 16899 7395
rect 17693 7361 17727 7395
rect 18153 7361 18187 7395
rect 18797 7361 18831 7395
rect 19441 7361 19475 7395
rect 20545 7361 20579 7395
rect 29469 7361 29503 7395
rect 33793 7361 33827 7395
rect 38301 7361 38335 7395
rect 1593 7293 1627 7327
rect 3985 7293 4019 7327
rect 4261 7293 4295 7327
rect 7941 7293 7975 7327
rect 10517 7293 10551 7327
rect 10701 7293 10735 7327
rect 14013 7293 14047 7327
rect 22109 7293 22143 7327
rect 22753 7293 22787 7327
rect 23949 7293 23983 7327
rect 7297 7225 7331 7259
rect 15117 7225 15151 7259
rect 19533 7225 19567 7259
rect 3341 7157 3375 7191
rect 13461 7157 13495 7191
rect 20637 7157 20671 7191
rect 1948 6953 1982 6987
rect 4248 6953 4282 6987
rect 7100 6953 7134 6987
rect 17601 6953 17635 6987
rect 22477 6953 22511 6987
rect 3985 6817 4019 6851
rect 6837 6817 6871 6851
rect 10333 6817 10367 6851
rect 13277 6817 13311 6851
rect 15853 6817 15887 6851
rect 16037 6817 16071 6851
rect 17049 6817 17083 6851
rect 20269 6817 20303 6851
rect 21005 6817 21039 6851
rect 21465 6817 21499 6851
rect 31953 6817 31987 6851
rect 1685 6749 1719 6783
rect 6009 6749 6043 6783
rect 9873 6749 9907 6783
rect 13093 6749 13127 6783
rect 14289 6749 14323 6783
rect 14473 6749 14507 6783
rect 16957 6749 16991 6783
rect 17785 6749 17819 6783
rect 18429 6749 18463 6783
rect 19441 6749 19475 6783
rect 19533 6749 19567 6783
rect 20177 6749 20211 6783
rect 20821 6749 20855 6783
rect 22661 6749 22695 6783
rect 31861 6749 31895 6783
rect 10609 6681 10643 6715
rect 3433 6613 3467 6647
rect 8585 6613 8619 6647
rect 9689 6613 9723 6647
rect 12081 6613 12115 6647
rect 13737 6613 13771 6647
rect 14933 6613 14967 6647
rect 16497 6613 16531 6647
rect 18245 6613 18279 6647
rect 15669 6409 15703 6443
rect 16129 6409 16163 6443
rect 18797 6409 18831 6443
rect 19441 6409 19475 6443
rect 20729 6409 20763 6443
rect 4077 6341 4111 6375
rect 4629 6341 4663 6375
rect 7297 6341 7331 6375
rect 14197 6341 14231 6375
rect 17049 6341 17083 6375
rect 20085 6341 20119 6375
rect 4537 6273 4571 6307
rect 5181 6273 5215 6307
rect 5273 6273 5307 6307
rect 5825 6273 5859 6307
rect 6561 6273 6595 6307
rect 7205 6273 7239 6307
rect 11161 6273 11195 6307
rect 16313 6273 16347 6307
rect 18245 6273 18279 6307
rect 18705 6273 18739 6307
rect 19349 6273 19383 6307
rect 19993 6273 20027 6307
rect 20637 6273 20671 6307
rect 21281 6273 21315 6307
rect 22293 6273 22327 6307
rect 29561 6273 29595 6307
rect 2053 6205 2087 6239
rect 2329 6205 2363 6239
rect 8125 6205 8159 6239
rect 8401 6205 8435 6239
rect 10149 6205 10183 6239
rect 11713 6205 11747 6239
rect 11989 6205 12023 6239
rect 13921 6205 13955 6239
rect 16957 6205 16991 6239
rect 17233 6205 17267 6239
rect 5917 6137 5951 6171
rect 10977 6137 11011 6171
rect 13461 6137 13495 6171
rect 21373 6137 21407 6171
rect 6653 6069 6687 6103
rect 18061 6069 18095 6103
rect 22385 6069 22419 6103
rect 29653 6069 29687 6103
rect 1856 5865 1890 5899
rect 7665 5865 7699 5899
rect 9321 5865 9355 5899
rect 9965 5865 9999 5899
rect 18521 5865 18555 5899
rect 19533 5865 19567 5899
rect 20821 5865 20855 5899
rect 21465 5865 21499 5899
rect 22109 5865 22143 5899
rect 3341 5797 3375 5831
rect 5365 5729 5399 5763
rect 8309 5729 8343 5763
rect 10517 5729 10551 5763
rect 12541 5729 12575 5763
rect 13093 5729 13127 5763
rect 13737 5729 13771 5763
rect 14289 5729 14323 5763
rect 16037 5729 16071 5763
rect 16497 5729 16531 5763
rect 1593 5661 1627 5695
rect 4169 5661 4203 5695
rect 5089 5661 5123 5695
rect 7573 5661 7607 5695
rect 8217 5661 8251 5695
rect 9229 5661 9263 5695
rect 9873 5661 9907 5695
rect 17141 5661 17175 5695
rect 17785 5661 17819 5695
rect 18429 5661 18463 5695
rect 19441 5661 19475 5695
rect 20085 5661 20119 5695
rect 20729 5661 20763 5695
rect 21373 5661 21407 5695
rect 22017 5661 22051 5695
rect 24777 5661 24811 5695
rect 35173 5661 35207 5695
rect 38025 5661 38059 5695
rect 7113 5593 7147 5627
rect 10793 5593 10827 5627
rect 13185 5593 13219 5627
rect 14565 5593 14599 5627
rect 17877 5593 17911 5627
rect 4077 5525 4111 5559
rect 4353 5525 4387 5559
rect 17233 5525 17267 5559
rect 20177 5525 20211 5559
rect 24593 5525 24627 5559
rect 34989 5525 35023 5559
rect 38209 5525 38243 5559
rect 4813 5321 4847 5355
rect 5457 5321 5491 5355
rect 15301 5321 15335 5355
rect 15853 5321 15887 5355
rect 18889 5321 18923 5355
rect 20821 5321 20855 5355
rect 8677 5253 8711 5287
rect 11989 5253 12023 5287
rect 14197 5253 14231 5287
rect 19533 5253 19567 5287
rect 1593 5185 1627 5219
rect 4721 5185 4755 5219
rect 5365 5185 5399 5219
rect 9137 5185 9171 5219
rect 11713 5185 11747 5219
rect 15209 5185 15243 5219
rect 16037 5185 16071 5219
rect 16865 5185 16899 5219
rect 16957 5185 16991 5219
rect 17693 5185 17727 5219
rect 18153 5185 18187 5219
rect 18797 5185 18831 5219
rect 19441 5185 19475 5219
rect 20085 5185 20119 5219
rect 20729 5185 20763 5219
rect 22017 5185 22051 5219
rect 22661 5185 22695 5219
rect 31125 5185 31159 5219
rect 31217 5185 31251 5219
rect 32481 5185 32515 5219
rect 37473 5185 37507 5219
rect 37565 5185 37599 5219
rect 38301 5185 38335 5219
rect 2421 5117 2455 5151
rect 2697 5117 2731 5151
rect 4169 5117 4203 5151
rect 6653 5117 6687 5151
rect 6929 5117 6963 5151
rect 9413 5117 9447 5151
rect 13461 5117 13495 5151
rect 14105 5117 14139 5151
rect 14657 5049 14691 5083
rect 18245 5049 18279 5083
rect 22109 5049 22143 5083
rect 1777 4981 1811 5015
rect 10885 4981 10919 5015
rect 17509 4981 17543 5015
rect 20177 4981 20211 5015
rect 22753 4981 22787 5015
rect 32321 4981 32355 5015
rect 38117 4981 38151 5015
rect 7757 4777 7791 4811
rect 16129 4777 16163 4811
rect 17509 4777 17543 4811
rect 19533 4777 19567 4811
rect 20821 4777 20855 4811
rect 21465 4777 21499 4811
rect 7113 4709 7147 4743
rect 15577 4709 15611 4743
rect 18613 4709 18647 4743
rect 2145 4641 2179 4675
rect 6561 4641 6595 4675
rect 10609 4641 10643 4675
rect 13277 4641 13311 4675
rect 20177 4641 20211 4675
rect 1869 4573 1903 4607
rect 2881 4573 2915 4607
rect 4537 4573 4571 4607
rect 7297 4573 7331 4607
rect 7941 4573 7975 4607
rect 8401 4573 8435 4607
rect 9137 4573 9171 4607
rect 9965 4573 9999 4607
rect 12633 4573 12667 4607
rect 13093 4573 13127 4607
rect 13737 4573 13771 4607
rect 15025 4573 15059 4607
rect 15485 4573 15519 4607
rect 16313 4573 16347 4607
rect 16773 4573 16807 4607
rect 17417 4573 17451 4607
rect 18797 4573 18831 4607
rect 19441 4573 19475 4607
rect 20085 4573 20119 4607
rect 20729 4573 20763 4607
rect 21373 4573 21407 4607
rect 22009 4573 22043 4607
rect 22661 4573 22695 4607
rect 3157 4505 3191 4539
rect 4813 4505 4847 4539
rect 8493 4505 8527 4539
rect 10885 4505 10919 4539
rect 14381 4505 14415 4539
rect 14473 4505 14507 4539
rect 16865 4505 16899 4539
rect 22109 4505 22143 4539
rect 9321 4437 9355 4471
rect 10057 4437 10091 4471
rect 22753 4437 22787 4471
rect 5917 4233 5951 4267
rect 17877 4165 17911 4199
rect 1869 4097 1903 4131
rect 2973 4097 3007 4131
rect 7113 4097 7147 4131
rect 10517 4097 10551 4131
rect 10977 4097 11011 4131
rect 11069 4097 11103 4131
rect 11713 4097 11747 4131
rect 17325 4097 17359 4131
rect 17785 4097 17819 4131
rect 18429 4097 18463 4131
rect 19073 4097 19107 4131
rect 19717 4097 19751 4131
rect 20361 4097 20395 4131
rect 21005 4097 21039 4131
rect 22017 4097 22051 4131
rect 22661 4097 22695 4131
rect 27353 4097 27387 4131
rect 2145 4029 2179 4063
rect 3249 4029 3283 4063
rect 4169 4029 4203 4063
rect 4445 4029 4479 4063
rect 7757 4029 7791 4063
rect 8033 4029 8067 4063
rect 9781 4029 9815 4063
rect 11989 4029 12023 4063
rect 14013 4029 14047 4063
rect 14289 4029 14323 4063
rect 18521 4029 18555 4063
rect 17141 3961 17175 3995
rect 22753 3961 22787 3995
rect 7205 3893 7239 3927
rect 10333 3893 10367 3927
rect 13461 3893 13495 3927
rect 15761 3893 15795 3927
rect 19165 3893 19199 3927
rect 19809 3893 19843 3927
rect 20453 3893 20487 3927
rect 21097 3893 21131 3927
rect 22109 3893 22143 3927
rect 27169 3893 27203 3927
rect 19533 3689 19567 3723
rect 21465 3689 21499 3723
rect 22477 3689 22511 3723
rect 23305 3689 23339 3723
rect 26709 3689 26743 3723
rect 38117 3689 38151 3723
rect 13737 3621 13771 3655
rect 16037 3621 16071 3655
rect 16589 3621 16623 3655
rect 2881 3553 2915 3587
rect 4261 3553 4295 3587
rect 6009 3553 6043 3587
rect 11529 3553 11563 3587
rect 11989 3553 12023 3587
rect 18613 3553 18647 3587
rect 22109 3553 22143 3587
rect 1685 3485 1719 3519
rect 2605 3485 2639 3519
rect 3985 3485 4019 3519
rect 4905 3485 4939 3519
rect 8033 3485 8067 3519
rect 9505 3485 9539 3519
rect 14289 3485 14323 3519
rect 16773 3485 16807 3519
rect 17233 3485 17267 3519
rect 17877 3485 17911 3519
rect 18521 3485 18555 3519
rect 19441 3485 19475 3519
rect 20085 3485 20119 3519
rect 20729 3485 20763 3519
rect 21373 3485 21407 3519
rect 22661 3485 22695 3519
rect 22753 3485 22787 3519
rect 23489 3485 23523 3519
rect 23765 3485 23799 3519
rect 26617 3485 26651 3519
rect 38301 3485 38335 3519
rect 1961 3417 1995 3451
rect 5181 3417 5215 3451
rect 6285 3417 6319 3451
rect 9781 3417 9815 3451
rect 12265 3417 12299 3451
rect 14565 3417 14599 3451
rect 17325 3417 17359 3451
rect 17969 3349 18003 3383
rect 20177 3349 20211 3383
rect 20821 3349 20855 3383
rect 22845 3349 22879 3383
rect 6929 3145 6963 3179
rect 13461 3145 13495 3179
rect 18153 3145 18187 3179
rect 23213 3145 23247 3179
rect 23949 3145 23983 3179
rect 36737 3145 36771 3179
rect 8224 3077 8258 3111
rect 10517 3077 10551 3111
rect 10609 3077 10643 3111
rect 11989 3077 12023 3111
rect 4169 3009 4203 3043
rect 6653 3009 6687 3043
rect 7941 3009 7975 3043
rect 11713 3009 11747 3043
rect 17049 3009 17083 3043
rect 17693 3009 17727 3043
rect 18797 3009 18831 3043
rect 19441 3009 19475 3043
rect 20085 3009 20119 3043
rect 20729 3009 20763 3043
rect 22017 3009 22051 3043
rect 22661 3009 22695 3043
rect 23121 3009 23155 3043
rect 23673 3009 23707 3043
rect 24133 3009 24167 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 1593 2941 1627 2975
rect 1869 2941 1903 2975
rect 5917 2941 5951 2975
rect 9965 2941 9999 2975
rect 11161 2941 11195 2975
rect 14002 2941 14036 2975
rect 3341 2873 3375 2907
rect 15761 2873 15795 2907
rect 16865 2873 16899 2907
rect 22753 2873 22787 2907
rect 4432 2805 4466 2839
rect 14270 2805 14304 2839
rect 17509 2805 17543 2839
rect 18889 2805 18923 2839
rect 19533 2805 19567 2839
rect 20177 2805 20211 2839
rect 20821 2805 20855 2839
rect 22109 2805 22143 2839
rect 38209 2805 38243 2839
rect 3433 2601 3467 2635
rect 11069 2601 11103 2635
rect 17509 2601 17543 2635
rect 22017 2601 22051 2635
rect 27169 2601 27203 2635
rect 29745 2601 29779 2635
rect 32321 2601 32355 2635
rect 34897 2601 34931 2635
rect 16865 2533 16899 2567
rect 24593 2533 24627 2567
rect 35541 2533 35575 2567
rect 36737 2533 36771 2567
rect 4169 2465 4203 2499
rect 6561 2465 6595 2499
rect 6837 2465 6871 2499
rect 9321 2465 9355 2499
rect 11713 2465 11747 2499
rect 14289 2465 14323 2499
rect 22753 2465 22787 2499
rect 1685 2397 1719 2431
rect 17049 2397 17083 2431
rect 17693 2397 17727 2431
rect 18613 2397 18647 2431
rect 19625 2397 19659 2431
rect 19901 2397 19935 2431
rect 21005 2397 21039 2431
rect 22201 2397 22235 2431
rect 22661 2397 22695 2431
rect 23305 2397 23339 2431
rect 24777 2397 24811 2431
rect 27353 2397 27387 2431
rect 27813 2397 27847 2431
rect 29929 2397 29963 2431
rect 31033 2397 31067 2431
rect 32505 2397 32539 2431
rect 35081 2397 35115 2431
rect 35725 2397 35759 2431
rect 36921 2397 36955 2431
rect 37473 2397 37507 2431
rect 1961 2329 1995 2363
rect 4445 2329 4479 2363
rect 8585 2329 8619 2363
rect 9597 2329 9631 2363
rect 11989 2329 12023 2363
rect 14565 2329 14599 2363
rect 5917 2261 5951 2295
rect 13461 2261 13495 2295
rect 16037 2261 16071 2295
rect 18797 2261 18831 2295
rect 19441 2261 19475 2295
rect 20085 2261 20119 2295
rect 20453 2261 20487 2295
rect 20821 2261 20855 2295
rect 23489 2261 23523 2295
rect 27997 2261 28031 2295
rect 31217 2261 31251 2295
rect 37657 2261 37691 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 7098 37272 7104 37324
rect 7156 37312 7162 37324
rect 7193 37315 7251 37321
rect 7193 37312 7205 37315
rect 7156 37284 7205 37312
rect 7156 37272 7162 37284
rect 7193 37281 7205 37284
rect 7239 37281 7251 37315
rect 7193 37275 7251 37281
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37244 1639 37247
rect 1854 37244 1860 37256
rect 1627 37216 1860 37244
rect 1627 37213 1639 37216
rect 1581 37207 1639 37213
rect 1854 37204 1860 37216
rect 1912 37204 1918 37256
rect 1946 37204 1952 37256
rect 2004 37244 2010 37256
rect 2501 37247 2559 37253
rect 2501 37244 2513 37247
rect 2004 37216 2513 37244
rect 2004 37204 2010 37216
rect 2501 37213 2513 37216
rect 2547 37213 2559 37247
rect 3142 37244 3148 37256
rect 3103 37216 3148 37244
rect 2501 37207 2559 37213
rect 3142 37204 3148 37216
rect 3200 37204 3206 37256
rect 3970 37244 3976 37256
rect 3931 37216 3976 37244
rect 3970 37204 3976 37216
rect 4028 37204 4034 37256
rect 5261 37247 5319 37253
rect 5261 37213 5273 37247
rect 5307 37244 5319 37247
rect 6730 37244 6736 37256
rect 5307 37216 6736 37244
rect 5307 37213 5319 37216
rect 5261 37207 5319 37213
rect 6730 37204 6736 37216
rect 6788 37204 6794 37256
rect 7466 37244 7472 37256
rect 7427 37216 7472 37244
rect 7466 37204 7472 37216
rect 7524 37204 7530 37256
rect 8386 37204 8392 37256
rect 8444 37244 8450 37256
rect 9309 37247 9367 37253
rect 9309 37244 9321 37247
rect 8444 37216 9321 37244
rect 8444 37204 8450 37216
rect 9309 37213 9321 37216
rect 9355 37213 9367 37247
rect 9309 37207 9367 37213
rect 10318 37204 10324 37256
rect 10376 37244 10382 37256
rect 10597 37247 10655 37253
rect 10597 37244 10609 37247
rect 10376 37216 10609 37244
rect 10376 37204 10382 37216
rect 10597 37213 10609 37216
rect 10643 37213 10655 37247
rect 10597 37207 10655 37213
rect 11606 37204 11612 37256
rect 11664 37244 11670 37256
rect 11885 37247 11943 37253
rect 11885 37244 11897 37247
rect 11664 37216 11897 37244
rect 11664 37204 11670 37216
rect 11885 37213 11897 37216
rect 11931 37213 11943 37247
rect 11885 37207 11943 37213
rect 12894 37204 12900 37256
rect 12952 37244 12958 37256
rect 13173 37247 13231 37253
rect 13173 37244 13185 37247
rect 12952 37216 13185 37244
rect 12952 37204 12958 37216
rect 13173 37213 13185 37216
rect 13219 37213 13231 37247
rect 14918 37244 14924 37256
rect 14879 37216 14924 37244
rect 13173 37207 13231 37213
rect 14918 37204 14924 37216
rect 14976 37204 14982 37256
rect 16850 37244 16856 37256
rect 16811 37216 16856 37244
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 18138 37244 18144 37256
rect 18099 37216 18144 37244
rect 18138 37204 18144 37216
rect 18196 37204 18202 37256
rect 19426 37244 19432 37256
rect 19387 37216 19432 37244
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 20714 37204 20720 37256
rect 20772 37244 20778 37256
rect 20901 37247 20959 37253
rect 20901 37244 20913 37247
rect 20772 37216 20913 37244
rect 20772 37204 20778 37216
rect 20901 37213 20913 37216
rect 20947 37213 20959 37247
rect 20901 37207 20959 37213
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 22612 37216 22845 37244
rect 22612 37204 22618 37216
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 22833 37207 22891 37213
rect 22922 37204 22928 37256
rect 22980 37244 22986 37256
rect 24581 37247 24639 37253
rect 24581 37244 24593 37247
rect 22980 37216 24593 37244
rect 22980 37204 22986 37216
rect 24581 37213 24593 37216
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 24670 37204 24676 37256
rect 24728 37244 24734 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 24728 37216 25881 37244
rect 24728 37204 24734 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 27062 37204 27068 37256
rect 27120 37244 27126 37256
rect 27341 37247 27399 37253
rect 27341 37244 27353 37247
rect 27120 37216 27353 37244
rect 27120 37204 27126 37216
rect 27341 37213 27353 37216
rect 27387 37213 27399 37247
rect 27341 37207 27399 37213
rect 27798 37204 27804 37256
rect 27856 37244 27862 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 27856 37216 29745 37244
rect 27856 37204 27862 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30653 37247 30711 37253
rect 30653 37244 30665 37247
rect 30432 37216 30665 37244
rect 30432 37204 30438 37216
rect 30653 37213 30665 37216
rect 30699 37213 30711 37247
rect 30653 37207 30711 37213
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 31812 37216 32505 37244
rect 31812 37204 31818 37216
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33560 37216 33793 37244
rect 33560 37204 33566 37216
rect 33781 37213 33793 37216
rect 33827 37213 33839 37247
rect 33781 37207 33839 37213
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34848 37216 35081 37244
rect 34848 37204 34854 37216
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 36722 37204 36728 37256
rect 36780 37244 36786 37256
rect 36909 37247 36967 37253
rect 36909 37244 36921 37247
rect 36780 37216 36921 37244
rect 36780 37204 36786 37216
rect 36909 37213 36921 37216
rect 36955 37213 36967 37247
rect 36909 37207 36967 37213
rect 38013 37247 38071 37253
rect 38013 37213 38025 37247
rect 38059 37213 38071 37247
rect 38013 37207 38071 37213
rect 2774 37176 2780 37188
rect 1780 37148 2780 37176
rect 1780 37117 1808 37148
rect 2774 37136 2780 37148
rect 2832 37136 2838 37188
rect 6546 37176 6552 37188
rect 2976 37148 6552 37176
rect 1765 37111 1823 37117
rect 1765 37077 1777 37111
rect 1811 37077 1823 37111
rect 1765 37071 1823 37077
rect 2317 37111 2375 37117
rect 2317 37077 2329 37111
rect 2363 37108 2375 37111
rect 2866 37108 2872 37120
rect 2363 37080 2872 37108
rect 2363 37077 2375 37080
rect 2317 37071 2375 37077
rect 2866 37068 2872 37080
rect 2924 37068 2930 37120
rect 2976 37117 3004 37148
rect 6546 37136 6552 37148
rect 6604 37136 6610 37188
rect 11974 37176 11980 37188
rect 10428 37148 11980 37176
rect 2961 37111 3019 37117
rect 2961 37077 2973 37111
rect 3007 37077 3019 37111
rect 2961 37071 3019 37077
rect 3878 37068 3884 37120
rect 3936 37108 3942 37120
rect 4157 37111 4215 37117
rect 4157 37108 4169 37111
rect 3936 37080 4169 37108
rect 3936 37068 3942 37080
rect 4157 37077 4169 37080
rect 4203 37077 4215 37111
rect 4157 37071 4215 37077
rect 5166 37068 5172 37120
rect 5224 37108 5230 37120
rect 5445 37111 5503 37117
rect 5445 37108 5457 37111
rect 5224 37080 5457 37108
rect 5224 37068 5230 37080
rect 5445 37077 5457 37080
rect 5491 37077 5503 37111
rect 9122 37108 9128 37120
rect 9083 37080 9128 37108
rect 5445 37071 5503 37077
rect 9122 37068 9128 37080
rect 9180 37068 9186 37120
rect 10428 37117 10456 37148
rect 11974 37136 11980 37148
rect 12032 37136 12038 37188
rect 31846 37136 31852 37188
rect 31904 37176 31910 37188
rect 31904 37148 34928 37176
rect 31904 37136 31910 37148
rect 10413 37111 10471 37117
rect 10413 37077 10425 37111
rect 10459 37077 10471 37111
rect 10413 37071 10471 37077
rect 10778 37068 10784 37120
rect 10836 37108 10842 37120
rect 11701 37111 11759 37117
rect 11701 37108 11713 37111
rect 10836 37080 11713 37108
rect 10836 37068 10842 37080
rect 11701 37077 11713 37080
rect 11747 37077 11759 37111
rect 12986 37108 12992 37120
rect 12947 37080 12992 37108
rect 11701 37071 11759 37077
rect 12986 37068 12992 37080
rect 13044 37068 13050 37120
rect 14826 37068 14832 37120
rect 14884 37108 14890 37120
rect 15105 37111 15163 37117
rect 15105 37108 15117 37111
rect 14884 37080 15117 37108
rect 14884 37068 14890 37080
rect 15105 37077 15117 37080
rect 15151 37077 15163 37111
rect 15105 37071 15163 37077
rect 16574 37068 16580 37120
rect 16632 37108 16638 37120
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 16632 37080 17049 37108
rect 16632 37068 16638 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 17037 37071 17095 37077
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18325 37111 18383 37117
rect 18325 37108 18337 37111
rect 18104 37080 18337 37108
rect 18104 37068 18110 37080
rect 18325 37077 18337 37080
rect 18371 37077 18383 37111
rect 18325 37071 18383 37077
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 19613 37111 19671 37117
rect 19613 37108 19625 37111
rect 19392 37080 19625 37108
rect 19392 37068 19398 37080
rect 19613 37077 19625 37080
rect 19659 37077 19671 37111
rect 20714 37108 20720 37120
rect 20675 37080 20720 37108
rect 19613 37071 19671 37077
rect 20714 37068 20720 37080
rect 20772 37068 20778 37120
rect 21726 37068 21732 37120
rect 21784 37108 21790 37120
rect 22649 37111 22707 37117
rect 22649 37108 22661 37111
rect 21784 37080 22661 37108
rect 21784 37068 21790 37080
rect 22649 37077 22661 37080
rect 22695 37077 22707 37111
rect 22649 37071 22707 37077
rect 23842 37068 23848 37120
rect 23900 37108 23906 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 23900 37080 24777 37108
rect 23900 37068 23906 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25774 37068 25780 37120
rect 25832 37108 25838 37120
rect 26053 37111 26111 37117
rect 26053 37108 26065 37111
rect 25832 37080 26065 37108
rect 25832 37068 25838 37080
rect 26053 37077 26065 37080
rect 26099 37077 26111 37111
rect 27154 37108 27160 37120
rect 27115 37080 27160 37108
rect 26053 37071 26111 37077
rect 27154 37068 27160 37080
rect 27212 37068 27218 37120
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29052 37080 29929 37108
rect 29052 37068 29058 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 30006 37068 30012 37120
rect 30064 37108 30070 37120
rect 30469 37111 30527 37117
rect 30469 37108 30481 37111
rect 30064 37080 30481 37108
rect 30064 37068 30070 37080
rect 30469 37077 30481 37080
rect 30515 37077 30527 37111
rect 32306 37108 32312 37120
rect 32267 37080 32312 37108
rect 30469 37071 30527 37077
rect 32306 37068 32312 37080
rect 32364 37068 32370 37120
rect 33594 37108 33600 37120
rect 33555 37080 33600 37108
rect 33594 37068 33600 37080
rect 33652 37068 33658 37120
rect 34900 37117 34928 37148
rect 35526 37136 35532 37188
rect 35584 37176 35590 37188
rect 38028 37176 38056 37207
rect 35584 37148 38056 37176
rect 35584 37136 35590 37148
rect 34885 37111 34943 37117
rect 34885 37077 34897 37111
rect 34931 37077 34943 37111
rect 34885 37071 34943 37077
rect 35894 37068 35900 37120
rect 35952 37108 35958 37120
rect 36725 37111 36783 37117
rect 36725 37108 36737 37111
rect 35952 37080 36737 37108
rect 35952 37068 35958 37080
rect 36725 37077 36737 37080
rect 36771 37077 36783 37111
rect 38194 37108 38200 37120
rect 38155 37080 38200 37108
rect 36725 37071 36783 37077
rect 38194 37068 38200 37080
rect 38252 37068 38258 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 658 36864 664 36916
rect 716 36904 722 36916
rect 1765 36907 1823 36913
rect 1765 36904 1777 36907
rect 716 36876 1777 36904
rect 716 36864 722 36876
rect 1765 36873 1777 36876
rect 1811 36873 1823 36907
rect 1765 36867 1823 36873
rect 1854 36864 1860 36916
rect 1912 36904 1918 36916
rect 2317 36907 2375 36913
rect 2317 36904 2329 36907
rect 1912 36876 2329 36904
rect 1912 36864 1918 36876
rect 2317 36873 2329 36876
rect 2363 36873 2375 36907
rect 2317 36867 2375 36873
rect 2866 36864 2872 36916
rect 2924 36904 2930 36916
rect 5442 36904 5448 36916
rect 2924 36876 5448 36904
rect 2924 36864 2930 36876
rect 5442 36864 5448 36876
rect 5500 36864 5506 36916
rect 29730 36864 29736 36916
rect 29788 36904 29794 36916
rect 33594 36904 33600 36916
rect 29788 36876 33600 36904
rect 29788 36864 29794 36876
rect 33594 36864 33600 36876
rect 33652 36864 33658 36916
rect 38197 36907 38255 36913
rect 38197 36873 38209 36907
rect 38243 36904 38255 36907
rect 38286 36904 38292 36916
rect 38243 36876 38292 36904
rect 38243 36873 38255 36876
rect 38197 36867 38255 36873
rect 38286 36864 38292 36876
rect 38344 36864 38350 36916
rect 39298 36836 39304 36848
rect 36924 36808 39304 36836
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36737 1639 36771
rect 2498 36768 2504 36780
rect 2459 36740 2504 36768
rect 1581 36731 1639 36737
rect 1596 36700 1624 36731
rect 2498 36728 2504 36740
rect 2556 36728 2562 36780
rect 36924 36777 36952 36808
rect 39298 36796 39304 36808
rect 39356 36796 39362 36848
rect 36909 36771 36967 36777
rect 36909 36737 36921 36771
rect 36955 36737 36967 36771
rect 36909 36731 36967 36737
rect 38013 36771 38071 36777
rect 38013 36737 38025 36771
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 4062 36700 4068 36712
rect 1596 36672 4068 36700
rect 4062 36660 4068 36672
rect 4120 36660 4126 36712
rect 35342 36660 35348 36712
rect 35400 36700 35406 36712
rect 38028 36700 38056 36731
rect 35400 36672 38056 36700
rect 35400 36660 35406 36672
rect 36722 36564 36728 36576
rect 36683 36536 36728 36564
rect 36722 36524 36728 36536
rect 36780 36524 36786 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1762 36156 1768 36168
rect 1723 36128 1768 36156
rect 1762 36116 1768 36128
rect 1820 36116 1826 36168
rect 38010 36116 38016 36168
rect 38068 36156 38074 36168
rect 38289 36159 38347 36165
rect 38289 36156 38301 36159
rect 38068 36128 38301 36156
rect 38068 36116 38074 36128
rect 38289 36125 38301 36128
rect 38335 36125 38347 36159
rect 38289 36119 38347 36125
rect 1581 36023 1639 36029
rect 1581 35989 1593 36023
rect 1627 36020 1639 36023
rect 2682 36020 2688 36032
rect 1627 35992 2688 36020
rect 1627 35989 1639 35992
rect 1581 35983 1639 35989
rect 2682 35980 2688 35992
rect 2740 35980 2746 36032
rect 34514 35980 34520 36032
rect 34572 36020 34578 36032
rect 38105 36023 38163 36029
rect 38105 36020 38117 36023
rect 34572 35992 38117 36020
rect 34572 35980 34578 35992
rect 38105 35989 38117 35992
rect 38151 35989 38163 36023
rect 38105 35983 38163 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 2498 35816 2504 35828
rect 2459 35788 2504 35816
rect 2498 35776 2504 35788
rect 2556 35776 2562 35828
rect 2406 35680 2412 35692
rect 2367 35652 2412 35680
rect 2406 35640 2412 35652
rect 2464 35640 2470 35692
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 4062 35232 4068 35284
rect 4120 35272 4126 35284
rect 5721 35275 5779 35281
rect 5721 35272 5733 35275
rect 4120 35244 5733 35272
rect 4120 35232 4126 35244
rect 5721 35241 5733 35244
rect 5767 35241 5779 35275
rect 5721 35235 5779 35241
rect 14918 35232 14924 35284
rect 14976 35272 14982 35284
rect 15105 35275 15163 35281
rect 15105 35272 15117 35275
rect 14976 35244 15117 35272
rect 14976 35232 14982 35244
rect 15105 35241 15117 35244
rect 15151 35241 15163 35275
rect 15105 35235 15163 35241
rect 16485 35275 16543 35281
rect 16485 35241 16497 35275
rect 16531 35272 16543 35275
rect 16850 35272 16856 35284
rect 16531 35244 16856 35272
rect 16531 35241 16543 35244
rect 16485 35235 16543 35241
rect 16850 35232 16856 35244
rect 16908 35232 16914 35284
rect 17405 35275 17463 35281
rect 17405 35241 17417 35275
rect 17451 35272 17463 35275
rect 18138 35272 18144 35284
rect 17451 35244 18144 35272
rect 17451 35241 17463 35244
rect 17405 35235 17463 35241
rect 18138 35232 18144 35244
rect 18196 35232 18202 35284
rect 21085 35275 21143 35281
rect 21085 35241 21097 35275
rect 21131 35272 21143 35275
rect 22922 35272 22928 35284
rect 21131 35244 22928 35272
rect 21131 35241 21143 35244
rect 21085 35235 21143 35241
rect 22922 35232 22928 35244
rect 22980 35232 22986 35284
rect 23201 35275 23259 35281
rect 23201 35241 23213 35275
rect 23247 35272 23259 35275
rect 24670 35272 24676 35284
rect 23247 35244 24676 35272
rect 23247 35241 23259 35244
rect 23201 35235 23259 35241
rect 24670 35232 24676 35244
rect 24728 35232 24734 35284
rect 5905 35071 5963 35077
rect 5905 35037 5917 35071
rect 5951 35068 5963 35071
rect 7190 35068 7196 35080
rect 5951 35040 7196 35068
rect 5951 35037 5963 35040
rect 5905 35031 5963 35037
rect 7190 35028 7196 35040
rect 7248 35028 7254 35080
rect 12069 35071 12127 35077
rect 12069 35037 12081 35071
rect 12115 35068 12127 35071
rect 12986 35068 12992 35080
rect 12115 35040 12992 35068
rect 12115 35037 12127 35040
rect 12069 35031 12127 35037
rect 12986 35028 12992 35040
rect 13044 35028 13050 35080
rect 15289 35071 15347 35077
rect 15289 35037 15301 35071
rect 15335 35068 15347 35071
rect 15654 35068 15660 35080
rect 15335 35040 15660 35068
rect 15335 35037 15347 35040
rect 15289 35031 15347 35037
rect 15654 35028 15660 35040
rect 15712 35028 15718 35080
rect 16666 35068 16672 35080
rect 16627 35040 16672 35068
rect 16666 35028 16672 35040
rect 16724 35028 16730 35080
rect 17586 35068 17592 35080
rect 17547 35040 17592 35068
rect 17586 35028 17592 35040
rect 17644 35028 17650 35080
rect 19978 35028 19984 35080
rect 20036 35068 20042 35080
rect 21269 35071 21327 35077
rect 21269 35068 21281 35071
rect 20036 35040 21281 35068
rect 20036 35028 20042 35040
rect 21269 35037 21281 35040
rect 21315 35037 21327 35071
rect 21269 35031 21327 35037
rect 22002 35028 22008 35080
rect 22060 35068 22066 35080
rect 23385 35071 23443 35077
rect 23385 35068 23397 35071
rect 22060 35040 23397 35068
rect 22060 35028 22066 35040
rect 23385 35037 23397 35040
rect 23431 35037 23443 35071
rect 23385 35031 23443 35037
rect 30469 35071 30527 35077
rect 30469 35037 30481 35071
rect 30515 35068 30527 35071
rect 31846 35068 31852 35080
rect 30515 35040 31852 35068
rect 30515 35037 30527 35040
rect 30469 35031 30527 35037
rect 31846 35028 31852 35040
rect 31904 35028 31910 35080
rect 35434 35028 35440 35080
rect 35492 35068 35498 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 35492 35040 38025 35068
rect 35492 35028 35498 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 11698 34892 11704 34944
rect 11756 34932 11762 34944
rect 12161 34935 12219 34941
rect 12161 34932 12173 34935
rect 11756 34904 12173 34932
rect 11756 34892 11762 34904
rect 12161 34901 12173 34904
rect 12207 34901 12219 34935
rect 30558 34932 30564 34944
rect 30519 34904 30564 34932
rect 12161 34895 12219 34901
rect 30558 34892 30564 34904
rect 30616 34892 30622 34944
rect 38194 34932 38200 34944
rect 38155 34904 38200 34932
rect 38194 34892 38200 34904
rect 38252 34892 38258 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 6730 34688 6736 34740
rect 6788 34728 6794 34740
rect 7929 34731 7987 34737
rect 7929 34728 7941 34731
rect 6788 34700 7941 34728
rect 6788 34688 6794 34700
rect 7929 34697 7941 34700
rect 7975 34697 7987 34731
rect 7929 34691 7987 34697
rect 18325 34731 18383 34737
rect 18325 34697 18337 34731
rect 18371 34728 18383 34731
rect 19426 34728 19432 34740
rect 18371 34700 19432 34728
rect 18371 34697 18383 34700
rect 18325 34691 18383 34697
rect 19426 34688 19432 34700
rect 19484 34688 19490 34740
rect 27157 34731 27215 34737
rect 27157 34697 27169 34731
rect 27203 34728 27215 34731
rect 27798 34728 27804 34740
rect 27203 34700 27804 34728
rect 27203 34697 27215 34700
rect 27157 34691 27215 34697
rect 27798 34688 27804 34700
rect 27856 34688 27862 34740
rect 1581 34595 1639 34601
rect 1581 34561 1593 34595
rect 1627 34592 1639 34595
rect 4062 34592 4068 34604
rect 1627 34564 4068 34592
rect 1627 34561 1639 34564
rect 1581 34555 1639 34561
rect 4062 34552 4068 34564
rect 4120 34552 4126 34604
rect 8113 34595 8171 34601
rect 8113 34561 8125 34595
rect 8159 34592 8171 34595
rect 9858 34592 9864 34604
rect 8159 34564 9864 34592
rect 8159 34561 8171 34564
rect 8113 34555 8171 34561
rect 9858 34552 9864 34564
rect 9916 34552 9922 34604
rect 11974 34592 11980 34604
rect 11935 34564 11980 34592
rect 11974 34552 11980 34564
rect 12032 34552 12038 34604
rect 18506 34592 18512 34604
rect 18467 34564 18512 34592
rect 18506 34552 18512 34564
rect 18564 34552 18570 34604
rect 19889 34595 19947 34601
rect 19889 34561 19901 34595
rect 19935 34592 19947 34595
rect 20714 34592 20720 34604
rect 19935 34564 20720 34592
rect 19935 34561 19947 34564
rect 19889 34555 19947 34561
rect 20714 34552 20720 34564
rect 20772 34552 20778 34604
rect 27338 34592 27344 34604
rect 27299 34564 27344 34592
rect 27338 34552 27344 34564
rect 27396 34552 27402 34604
rect 33229 34595 33287 34601
rect 33229 34561 33241 34595
rect 33275 34592 33287 34595
rect 34514 34592 34520 34604
rect 33275 34564 34520 34592
rect 33275 34561 33287 34564
rect 33229 34555 33287 34561
rect 34514 34552 34520 34564
rect 34572 34552 34578 34604
rect 12069 34527 12127 34533
rect 12069 34493 12081 34527
rect 12115 34524 12127 34527
rect 12158 34524 12164 34536
rect 12115 34496 12164 34524
rect 12115 34493 12127 34496
rect 12069 34487 12127 34493
rect 12158 34484 12164 34496
rect 12216 34484 12222 34536
rect 19058 34484 19064 34536
rect 19116 34524 19122 34536
rect 19981 34527 20039 34533
rect 19981 34524 19993 34527
rect 19116 34496 19993 34524
rect 19116 34484 19122 34496
rect 19981 34493 19993 34496
rect 20027 34493 20039 34527
rect 33318 34524 33324 34536
rect 33279 34496 33324 34524
rect 19981 34487 20039 34493
rect 33318 34484 33324 34496
rect 33376 34484 33382 34536
rect 1762 34388 1768 34400
rect 1723 34360 1768 34388
rect 1762 34348 1768 34360
rect 1820 34348 1826 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 7190 34184 7196 34196
rect 7151 34156 7196 34184
rect 7190 34144 7196 34156
rect 7248 34144 7254 34196
rect 25961 34187 26019 34193
rect 25961 34153 25973 34187
rect 26007 34184 26019 34187
rect 27338 34184 27344 34196
rect 26007 34156 27344 34184
rect 26007 34153 26019 34156
rect 25961 34147 26019 34153
rect 27338 34144 27344 34156
rect 27396 34144 27402 34196
rect 34885 34187 34943 34193
rect 34885 34153 34897 34187
rect 34931 34184 34943 34187
rect 35342 34184 35348 34196
rect 34931 34156 35348 34184
rect 34931 34153 34943 34156
rect 34885 34147 34943 34153
rect 35342 34144 35348 34156
rect 35400 34144 35406 34196
rect 7098 33980 7104 33992
rect 7059 33952 7104 33980
rect 7098 33940 7104 33952
rect 7156 33940 7162 33992
rect 21726 33980 21732 33992
rect 21687 33952 21732 33980
rect 21726 33940 21732 33952
rect 21784 33940 21790 33992
rect 23198 33940 23204 33992
rect 23256 33980 23262 33992
rect 25869 33983 25927 33989
rect 25869 33980 25881 33983
rect 23256 33952 25881 33980
rect 23256 33940 23262 33952
rect 25869 33949 25881 33952
rect 25915 33949 25927 33983
rect 29730 33980 29736 33992
rect 29691 33952 29736 33980
rect 25869 33943 25927 33949
rect 29730 33940 29736 33952
rect 29788 33940 29794 33992
rect 30098 33940 30104 33992
rect 30156 33980 30162 33992
rect 35069 33983 35127 33989
rect 35069 33980 35081 33983
rect 30156 33952 35081 33980
rect 30156 33940 30162 33952
rect 35069 33949 35081 33952
rect 35115 33949 35127 33983
rect 35069 33943 35127 33949
rect 21818 33844 21824 33856
rect 21779 33816 21824 33844
rect 21818 33804 21824 33816
rect 21876 33804 21882 33856
rect 29822 33844 29828 33856
rect 29783 33816 29828 33844
rect 29822 33804 29828 33816
rect 29880 33804 29886 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 19334 33600 19340 33652
rect 19392 33640 19398 33652
rect 29822 33640 29828 33652
rect 19392 33612 29828 33640
rect 19392 33600 19398 33612
rect 29822 33600 29828 33612
rect 29880 33600 29886 33652
rect 10778 33504 10784 33516
rect 10739 33476 10784 33504
rect 10778 33464 10784 33476
rect 10836 33464 10842 33516
rect 35342 33464 35348 33516
rect 35400 33504 35406 33516
rect 38013 33507 38071 33513
rect 38013 33504 38025 33507
rect 35400 33476 38025 33504
rect 35400 33464 35406 33476
rect 38013 33473 38025 33476
rect 38059 33473 38071 33507
rect 38013 33467 38071 33473
rect 38194 33368 38200 33380
rect 38155 33340 38200 33368
rect 38194 33328 38200 33340
rect 38252 33328 38258 33380
rect 10134 33260 10140 33312
rect 10192 33300 10198 33312
rect 10873 33303 10931 33309
rect 10873 33300 10885 33303
rect 10192 33272 10885 33300
rect 10192 33260 10198 33272
rect 10873 33269 10885 33272
rect 10919 33269 10931 33303
rect 10873 33263 10931 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1762 32892 1768 32904
rect 1723 32864 1768 32892
rect 1762 32852 1768 32864
rect 1820 32852 1826 32904
rect 1581 32759 1639 32765
rect 1581 32725 1593 32759
rect 1627 32756 1639 32759
rect 5534 32756 5540 32768
rect 1627 32728 5540 32756
rect 1627 32725 1639 32728
rect 1581 32719 1639 32725
rect 5534 32716 5540 32728
rect 5592 32716 5598 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 34701 32555 34759 32561
rect 34701 32521 34713 32555
rect 34747 32552 34759 32555
rect 35526 32552 35532 32564
rect 34747 32524 35532 32552
rect 34747 32521 34759 32524
rect 34701 32515 34759 32521
rect 35526 32512 35532 32524
rect 35584 32512 35590 32564
rect 6546 32416 6552 32428
rect 6507 32388 6552 32416
rect 6546 32376 6552 32388
rect 6604 32376 6610 32428
rect 7098 32376 7104 32428
rect 7156 32416 7162 32428
rect 20162 32416 20168 32428
rect 7156 32388 20168 32416
rect 7156 32376 7162 32388
rect 20162 32376 20168 32388
rect 20220 32376 20226 32428
rect 23201 32419 23259 32425
rect 23201 32385 23213 32419
rect 23247 32416 23259 32419
rect 27154 32416 27160 32428
rect 23247 32388 27160 32416
rect 23247 32385 23259 32388
rect 23201 32379 23259 32385
rect 27154 32376 27160 32388
rect 27212 32376 27218 32428
rect 29914 32376 29920 32428
rect 29972 32416 29978 32428
rect 34885 32419 34943 32425
rect 34885 32416 34897 32419
rect 29972 32388 34897 32416
rect 29972 32376 29978 32388
rect 34885 32385 34897 32388
rect 34931 32385 34943 32419
rect 34885 32379 34943 32385
rect 28994 32308 29000 32360
rect 29052 32348 29058 32360
rect 30006 32348 30012 32360
rect 29052 32320 30012 32348
rect 29052 32308 29058 32320
rect 30006 32308 30012 32320
rect 30064 32308 30070 32360
rect 6638 32212 6644 32224
rect 6599 32184 6644 32212
rect 6638 32172 6644 32184
rect 6696 32172 6702 32224
rect 18782 32172 18788 32224
rect 18840 32212 18846 32224
rect 23293 32215 23351 32221
rect 23293 32212 23305 32215
rect 18840 32184 23305 32212
rect 18840 32172 18846 32184
rect 23293 32181 23305 32184
rect 23339 32181 23351 32215
rect 23293 32175 23351 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 9858 32008 9864 32020
rect 9819 31980 9864 32008
rect 9858 31968 9864 31980
rect 9916 31968 9922 32020
rect 32306 32008 32312 32020
rect 29288 31980 32312 32008
rect 18414 31900 18420 31952
rect 18472 31940 18478 31952
rect 26053 31943 26111 31949
rect 26053 31940 26065 31943
rect 18472 31912 26065 31940
rect 18472 31900 18478 31912
rect 26053 31909 26065 31912
rect 26099 31909 26111 31943
rect 26053 31903 26111 31909
rect 28994 31872 29000 31884
rect 25148 31844 29000 31872
rect 5442 31764 5448 31816
rect 5500 31804 5506 31816
rect 8389 31807 8447 31813
rect 8389 31804 8401 31807
rect 5500 31776 8401 31804
rect 5500 31764 5506 31776
rect 8389 31773 8401 31776
rect 8435 31773 8447 31807
rect 8389 31767 8447 31773
rect 8481 31807 8539 31813
rect 8481 31773 8493 31807
rect 8527 31804 8539 31807
rect 8846 31804 8852 31816
rect 8527 31776 8852 31804
rect 8527 31773 8539 31776
rect 8481 31767 8539 31773
rect 8846 31764 8852 31776
rect 8904 31764 8910 31816
rect 9122 31804 9128 31816
rect 9083 31776 9128 31804
rect 9122 31764 9128 31776
rect 9180 31764 9186 31816
rect 9217 31807 9275 31813
rect 9217 31773 9229 31807
rect 9263 31804 9275 31807
rect 9306 31804 9312 31816
rect 9263 31776 9312 31804
rect 9263 31773 9275 31776
rect 9217 31767 9275 31773
rect 9306 31764 9312 31776
rect 9364 31764 9370 31816
rect 9769 31807 9827 31813
rect 9769 31773 9781 31807
rect 9815 31804 9827 31807
rect 10870 31804 10876 31816
rect 9815 31776 10876 31804
rect 9815 31773 9827 31776
rect 9769 31767 9827 31773
rect 10870 31764 10876 31776
rect 10928 31764 10934 31816
rect 25148 31813 25176 31844
rect 28994 31832 29000 31844
rect 29052 31832 29058 31884
rect 25133 31807 25191 31813
rect 25133 31773 25145 31807
rect 25179 31773 25191 31807
rect 25133 31767 25191 31773
rect 25222 31764 25228 31816
rect 25280 31804 25286 31816
rect 25961 31807 26019 31813
rect 25280 31776 25325 31804
rect 25280 31764 25286 31776
rect 25961 31773 25973 31807
rect 26007 31804 26019 31807
rect 29288 31804 29316 31980
rect 32306 31968 32312 31980
rect 32364 31968 32370 32020
rect 36998 31900 37004 31952
rect 37056 31940 37062 31952
rect 38105 31943 38163 31949
rect 38105 31940 38117 31943
rect 37056 31912 38117 31940
rect 37056 31900 37062 31912
rect 38105 31909 38117 31912
rect 38151 31909 38163 31943
rect 38105 31903 38163 31909
rect 29822 31872 29828 31884
rect 29783 31844 29828 31872
rect 29822 31832 29828 31844
rect 29880 31832 29886 31884
rect 26007 31776 29316 31804
rect 29733 31807 29791 31813
rect 26007 31773 26019 31776
rect 25961 31767 26019 31773
rect 29733 31773 29745 31807
rect 29779 31804 29791 31807
rect 35894 31804 35900 31816
rect 29779 31776 35900 31804
rect 29779 31773 29791 31776
rect 29733 31767 29791 31773
rect 35894 31764 35900 31776
rect 35952 31764 35958 31816
rect 38286 31804 38292 31816
rect 38247 31776 38292 31804
rect 38286 31764 38292 31776
rect 38344 31764 38350 31816
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 30745 31331 30803 31337
rect 30745 31297 30757 31331
rect 30791 31328 30803 31331
rect 36722 31328 36728 31340
rect 30791 31300 36728 31328
rect 30791 31297 30803 31300
rect 30745 31291 30803 31297
rect 36722 31288 36728 31300
rect 36780 31288 36786 31340
rect 20438 31084 20444 31136
rect 20496 31124 20502 31136
rect 30837 31127 30895 31133
rect 30837 31124 30849 31127
rect 20496 31096 30849 31124
rect 20496 31084 20502 31096
rect 30837 31093 30849 31096
rect 30883 31093 30895 31127
rect 30837 31087 30895 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 4062 30880 4068 30932
rect 4120 30920 4126 30932
rect 4157 30923 4215 30929
rect 4157 30920 4169 30923
rect 4120 30892 4169 30920
rect 4120 30880 4126 30892
rect 4157 30889 4169 30892
rect 4203 30889 4215 30923
rect 4157 30883 4215 30889
rect 16666 30880 16672 30932
rect 16724 30920 16730 30932
rect 17313 30923 17371 30929
rect 17313 30920 17325 30923
rect 16724 30892 17325 30920
rect 16724 30880 16730 30892
rect 17313 30889 17325 30892
rect 17359 30889 17371 30923
rect 17313 30883 17371 30889
rect 34885 30923 34943 30929
rect 34885 30889 34897 30923
rect 34931 30920 34943 30923
rect 35434 30920 35440 30932
rect 34931 30892 35440 30920
rect 34931 30889 34943 30892
rect 34885 30883 34943 30889
rect 35434 30880 35440 30892
rect 35492 30880 35498 30932
rect 1762 30716 1768 30728
rect 1723 30688 1768 30716
rect 1762 30676 1768 30688
rect 1820 30676 1826 30728
rect 4341 30719 4399 30725
rect 4341 30685 4353 30719
rect 4387 30716 4399 30719
rect 6086 30716 6092 30728
rect 4387 30688 6092 30716
rect 4387 30685 4399 30688
rect 4341 30679 4399 30685
rect 6086 30676 6092 30688
rect 6144 30676 6150 30728
rect 17221 30719 17279 30725
rect 17221 30685 17233 30719
rect 17267 30716 17279 30719
rect 17402 30716 17408 30728
rect 17267 30688 17408 30716
rect 17267 30685 17279 30688
rect 17221 30679 17279 30685
rect 17402 30676 17408 30688
rect 17460 30676 17466 30728
rect 30006 30676 30012 30728
rect 30064 30716 30070 30728
rect 35069 30719 35127 30725
rect 35069 30716 35081 30719
rect 30064 30688 35081 30716
rect 30064 30676 30070 30688
rect 35069 30685 35081 30688
rect 35115 30685 35127 30719
rect 35069 30679 35127 30685
rect 1581 30583 1639 30589
rect 1581 30549 1593 30583
rect 1627 30580 1639 30583
rect 3786 30580 3792 30592
rect 1627 30552 3792 30580
rect 1627 30549 1639 30552
rect 1581 30543 1639 30549
rect 3786 30540 3792 30552
rect 3844 30540 3850 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 15654 30308 15660 30320
rect 15615 30280 15660 30308
rect 15654 30268 15660 30280
rect 15712 30268 15718 30320
rect 15565 30243 15623 30249
rect 15565 30209 15577 30243
rect 15611 30240 15623 30243
rect 16022 30240 16028 30252
rect 15611 30212 16028 30240
rect 15611 30209 15623 30212
rect 15565 30203 15623 30209
rect 16022 30200 16028 30212
rect 16080 30200 16086 30252
rect 38286 30240 38292 30252
rect 38247 30212 38292 30240
rect 38286 30200 38292 30212
rect 38344 30200 38350 30252
rect 34146 29996 34152 30048
rect 34204 30036 34210 30048
rect 38105 30039 38163 30045
rect 38105 30036 38117 30039
rect 34204 30008 38117 30036
rect 34204 29996 34210 30008
rect 38105 30005 38117 30008
rect 38151 30005 38163 30039
rect 38105 29999 38163 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 6086 29832 6092 29844
rect 6047 29804 6092 29832
rect 6086 29792 6092 29804
rect 6144 29792 6150 29844
rect 17221 29835 17279 29841
rect 17221 29801 17233 29835
rect 17267 29832 17279 29835
rect 17586 29832 17592 29844
rect 17267 29804 17592 29832
rect 17267 29801 17279 29804
rect 17221 29795 17279 29801
rect 17586 29792 17592 29804
rect 17644 29792 17650 29844
rect 19521 29835 19579 29841
rect 19521 29801 19533 29835
rect 19567 29832 19579 29835
rect 19978 29832 19984 29844
rect 19567 29804 19984 29832
rect 19567 29801 19579 29804
rect 19521 29795 19579 29801
rect 19978 29792 19984 29804
rect 20036 29792 20042 29844
rect 22002 29832 22008 29844
rect 21963 29804 22008 29832
rect 22002 29792 22008 29804
rect 22060 29792 22066 29844
rect 34885 29835 34943 29841
rect 34885 29801 34897 29835
rect 34931 29832 34943 29835
rect 35342 29832 35348 29844
rect 34931 29804 35348 29832
rect 34931 29801 34943 29804
rect 34885 29795 34943 29801
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29597 1639 29631
rect 1581 29591 1639 29597
rect 1596 29560 1624 29591
rect 2682 29588 2688 29640
rect 2740 29628 2746 29640
rect 3973 29631 4031 29637
rect 3973 29628 3985 29631
rect 2740 29600 3985 29628
rect 2740 29588 2746 29600
rect 3973 29597 3985 29600
rect 4019 29597 4031 29631
rect 3973 29591 4031 29597
rect 5997 29631 6055 29637
rect 5997 29597 6009 29631
rect 6043 29628 6055 29631
rect 7650 29628 7656 29640
rect 6043 29600 7656 29628
rect 6043 29597 6055 29600
rect 5997 29591 6055 29597
rect 7650 29588 7656 29600
rect 7708 29588 7714 29640
rect 17129 29631 17187 29637
rect 17129 29597 17141 29631
rect 17175 29628 17187 29631
rect 17586 29628 17592 29640
rect 17175 29600 17592 29628
rect 17175 29597 17187 29600
rect 17129 29591 17187 29597
rect 17586 29588 17592 29600
rect 17644 29588 17650 29640
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 2774 29560 2780 29572
rect 1596 29532 2780 29560
rect 2774 29520 2780 29532
rect 2832 29520 2838 29572
rect 16758 29520 16764 29572
rect 16816 29560 16822 29572
rect 19444 29560 19472 29591
rect 20622 29588 20628 29640
rect 20680 29628 20686 29640
rect 21913 29631 21971 29637
rect 21913 29628 21925 29631
rect 20680 29600 21925 29628
rect 20680 29588 20686 29600
rect 21913 29597 21925 29600
rect 21959 29597 21971 29631
rect 21913 29591 21971 29597
rect 34698 29588 34704 29640
rect 34756 29628 34762 29640
rect 35069 29631 35127 29637
rect 35069 29628 35081 29631
rect 34756 29600 35081 29628
rect 34756 29588 34762 29600
rect 35069 29597 35081 29600
rect 35115 29597 35127 29631
rect 35069 29591 35127 29597
rect 16816 29532 19472 29560
rect 16816 29520 16822 29532
rect 1762 29492 1768 29504
rect 1723 29464 1768 29492
rect 1762 29452 1768 29464
rect 1820 29452 1826 29504
rect 4062 29492 4068 29504
rect 4023 29464 4068 29492
rect 4062 29452 4068 29464
rect 4120 29452 4126 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 18049 29291 18107 29297
rect 18049 29257 18061 29291
rect 18095 29288 18107 29291
rect 18506 29288 18512 29300
rect 18095 29260 18512 29288
rect 18095 29257 18107 29260
rect 18049 29251 18107 29257
rect 18506 29248 18512 29260
rect 18564 29248 18570 29300
rect 29181 29291 29239 29297
rect 29181 29257 29193 29291
rect 29227 29288 29239 29291
rect 30098 29288 30104 29300
rect 29227 29260 30104 29288
rect 29227 29257 29239 29260
rect 29181 29251 29239 29257
rect 30098 29248 30104 29260
rect 30156 29248 30162 29300
rect 17954 29152 17960 29164
rect 17915 29124 17960 29152
rect 17954 29112 17960 29124
rect 18012 29112 18018 29164
rect 29086 29152 29092 29164
rect 29047 29124 29092 29152
rect 29086 29112 29092 29124
rect 29144 29112 29150 29164
rect 38010 29152 38016 29164
rect 37971 29124 38016 29152
rect 38010 29112 38016 29124
rect 38068 29112 38074 29164
rect 2774 28976 2780 29028
rect 2832 29016 2838 29028
rect 38194 29016 38200 29028
rect 2832 28988 4108 29016
rect 38155 28988 38200 29016
rect 2832 28976 2838 28988
rect 4080 28960 4108 28988
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 4062 28908 4068 28960
rect 4120 28908 4126 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 29825 28747 29883 28753
rect 29825 28713 29837 28747
rect 29871 28744 29883 28747
rect 29914 28744 29920 28756
rect 29871 28716 29920 28744
rect 29871 28713 29883 28716
rect 29825 28707 29883 28713
rect 29914 28704 29920 28716
rect 29972 28704 29978 28756
rect 5534 28500 5540 28552
rect 5592 28540 5598 28552
rect 6917 28543 6975 28549
rect 6917 28540 6929 28543
rect 5592 28512 6929 28540
rect 5592 28500 5598 28512
rect 6917 28509 6929 28512
rect 6963 28509 6975 28543
rect 29730 28540 29736 28552
rect 29691 28512 29736 28540
rect 6917 28503 6975 28509
rect 29730 28500 29736 28512
rect 29788 28500 29794 28552
rect 7006 28404 7012 28416
rect 6967 28376 7012 28404
rect 7006 28364 7012 28376
rect 7064 28364 7070 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 1762 28064 1768 28076
rect 1723 28036 1768 28064
rect 1762 28024 1768 28036
rect 1820 28024 1826 28076
rect 32309 28067 32367 28073
rect 32309 28033 32321 28067
rect 32355 28064 32367 28067
rect 36998 28064 37004 28076
rect 32355 28036 37004 28064
rect 32355 28033 32367 28036
rect 32309 28027 32367 28033
rect 36998 28024 37004 28036
rect 37056 28024 37062 28076
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 3878 27860 3884 27872
rect 1627 27832 3884 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 3878 27820 3884 27832
rect 3936 27820 3942 27872
rect 32398 27860 32404 27872
rect 32359 27832 32404 27860
rect 32398 27820 32404 27832
rect 32456 27820 32462 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 3786 27412 3792 27464
rect 3844 27452 3850 27464
rect 7469 27455 7527 27461
rect 7469 27452 7481 27455
rect 3844 27424 7481 27452
rect 3844 27412 3850 27424
rect 7469 27421 7481 27424
rect 7515 27421 7527 27455
rect 34146 27452 34152 27464
rect 34107 27424 34152 27452
rect 7469 27415 7527 27421
rect 34146 27412 34152 27424
rect 34204 27412 34210 27464
rect 7561 27319 7619 27325
rect 7561 27285 7573 27319
rect 7607 27316 7619 27319
rect 8570 27316 8576 27328
rect 7607 27288 8576 27316
rect 7607 27285 7619 27288
rect 7561 27279 7619 27285
rect 8570 27276 8576 27288
rect 8628 27276 8634 27328
rect 20714 27276 20720 27328
rect 20772 27316 20778 27328
rect 34241 27319 34299 27325
rect 34241 27316 34253 27319
rect 20772 27288 34253 27316
rect 20772 27276 20778 27288
rect 34241 27285 34253 27288
rect 34287 27285 34299 27319
rect 34241 27279 34299 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 34790 26936 34796 26988
rect 34848 26976 34854 26988
rect 38013 26979 38071 26985
rect 38013 26976 38025 26979
rect 34848 26948 38025 26976
rect 34848 26936 34854 26948
rect 38013 26945 38025 26948
rect 38059 26945 38071 26979
rect 38013 26939 38071 26945
rect 38194 26772 38200 26784
rect 38155 26744 38200 26772
rect 38194 26732 38200 26744
rect 38252 26732 38258 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 29825 26571 29883 26577
rect 29825 26537 29837 26571
rect 29871 26568 29883 26571
rect 30006 26568 30012 26580
rect 29871 26540 30012 26568
rect 29871 26537 29883 26540
rect 29825 26531 29883 26537
rect 30006 26528 30012 26540
rect 30064 26528 30070 26580
rect 1581 26503 1639 26509
rect 1581 26469 1593 26503
rect 1627 26500 1639 26503
rect 5074 26500 5080 26512
rect 1627 26472 5080 26500
rect 1627 26469 1639 26472
rect 1581 26463 1639 26469
rect 5074 26460 5080 26472
rect 5132 26460 5138 26512
rect 1762 26364 1768 26376
rect 1723 26336 1768 26364
rect 1762 26324 1768 26336
rect 1820 26324 1826 26376
rect 29638 26324 29644 26376
rect 29696 26364 29702 26376
rect 29733 26367 29791 26373
rect 29733 26364 29745 26367
rect 29696 26336 29745 26364
rect 29696 26324 29702 26336
rect 29733 26333 29745 26336
rect 29779 26333 29791 26367
rect 29733 26327 29791 26333
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 4062 26024 4068 26036
rect 4023 25996 4068 26024
rect 4062 25984 4068 25996
rect 4120 25984 4126 26036
rect 4249 25891 4307 25897
rect 4249 25857 4261 25891
rect 4295 25888 4307 25891
rect 4614 25888 4620 25900
rect 4295 25860 4620 25888
rect 4295 25857 4307 25860
rect 4249 25851 4307 25857
rect 4614 25848 4620 25860
rect 4672 25848 4678 25900
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 28813 25483 28871 25489
rect 28813 25449 28825 25483
rect 28859 25480 28871 25483
rect 34698 25480 34704 25492
rect 28859 25452 34704 25480
rect 28859 25449 28871 25452
rect 28813 25443 28871 25449
rect 34698 25440 34704 25452
rect 34756 25440 34762 25492
rect 28718 25276 28724 25288
rect 28679 25248 28724 25276
rect 28718 25236 28724 25248
rect 28776 25236 28782 25288
rect 38286 25276 38292 25288
rect 38247 25248 38292 25276
rect 38286 25236 38292 25248
rect 38344 25236 38350 25288
rect 34606 25100 34612 25152
rect 34664 25140 34670 25152
rect 38105 25143 38163 25149
rect 38105 25140 38117 25143
rect 34664 25112 38117 25140
rect 34664 25100 34670 25112
rect 38105 25109 38117 25112
rect 38151 25109 38163 25143
rect 38105 25103 38163 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24800 1639 24803
rect 5442 24800 5448 24812
rect 1627 24772 5448 24800
rect 1627 24769 1639 24772
rect 1581 24763 1639 24769
rect 5442 24760 5448 24772
rect 5500 24760 5506 24812
rect 19058 24800 19064 24812
rect 19019 24772 19064 24800
rect 19058 24760 19064 24772
rect 19116 24760 19122 24812
rect 32030 24760 32036 24812
rect 32088 24800 32094 24812
rect 34977 24803 35035 24809
rect 34977 24800 34989 24803
rect 32088 24772 34989 24800
rect 32088 24760 32094 24772
rect 34977 24769 34989 24772
rect 35023 24769 35035 24803
rect 34977 24763 35035 24769
rect 17126 24732 17132 24744
rect 17087 24704 17132 24732
rect 17126 24692 17132 24704
rect 17184 24692 17190 24744
rect 18138 24692 18144 24744
rect 18196 24732 18202 24744
rect 19245 24735 19303 24741
rect 19245 24732 19257 24735
rect 18196 24704 19257 24732
rect 18196 24692 18202 24704
rect 19245 24701 19257 24704
rect 19291 24701 19303 24735
rect 19245 24695 19303 24701
rect 19978 24692 19984 24744
rect 20036 24732 20042 24744
rect 20165 24735 20223 24741
rect 20165 24732 20177 24735
rect 20036 24704 20177 24732
rect 20036 24692 20042 24704
rect 20165 24701 20177 24704
rect 20211 24701 20223 24735
rect 20165 24695 20223 24701
rect 34793 24667 34851 24673
rect 34793 24633 34805 24667
rect 34839 24664 34851 24667
rect 38010 24664 38016 24676
rect 34839 24636 38016 24664
rect 34839 24633 34851 24636
rect 34793 24627 34851 24633
rect 38010 24624 38016 24636
rect 38068 24624 38074 24676
rect 1762 24596 1768 24608
rect 1723 24568 1768 24596
rect 1762 24556 1768 24568
rect 1820 24556 1826 24608
rect 19426 24596 19432 24608
rect 19387 24568 19432 24596
rect 19426 24556 19432 24568
rect 19484 24556 19490 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 18138 24392 18144 24404
rect 18099 24364 18144 24392
rect 18138 24352 18144 24364
rect 18196 24352 18202 24404
rect 19978 24256 19984 24268
rect 19939 24228 19984 24256
rect 19978 24216 19984 24228
rect 20036 24216 20042 24268
rect 20622 24256 20628 24268
rect 20583 24228 20628 24256
rect 20622 24216 20628 24228
rect 20680 24216 20686 24268
rect 16114 24148 16120 24200
rect 16172 24188 16178 24200
rect 16853 24191 16911 24197
rect 16853 24188 16865 24191
rect 16172 24160 16865 24188
rect 16172 24148 16178 24160
rect 16853 24157 16865 24160
rect 16899 24157 16911 24191
rect 16853 24151 16911 24157
rect 16942 24148 16948 24200
rect 17000 24188 17006 24200
rect 17313 24191 17371 24197
rect 17313 24188 17325 24191
rect 17000 24160 17325 24188
rect 17000 24148 17006 24160
rect 17313 24157 17325 24160
rect 17359 24157 17371 24191
rect 18046 24188 18052 24200
rect 18007 24160 18052 24188
rect 17313 24151 17371 24157
rect 18046 24148 18052 24160
rect 18104 24148 18110 24200
rect 18322 24148 18328 24200
rect 18380 24188 18386 24200
rect 18877 24191 18935 24197
rect 18877 24188 18889 24191
rect 18380 24160 18889 24188
rect 18380 24148 18386 24160
rect 18877 24157 18889 24160
rect 18923 24157 18935 24191
rect 18877 24151 18935 24157
rect 20073 24123 20131 24129
rect 20073 24089 20085 24123
rect 20119 24089 20131 24123
rect 20073 24083 20131 24089
rect 16669 24055 16727 24061
rect 16669 24021 16681 24055
rect 16715 24052 16727 24055
rect 17218 24052 17224 24064
rect 16715 24024 17224 24052
rect 16715 24021 16727 24024
rect 16669 24015 16727 24021
rect 17218 24012 17224 24024
rect 17276 24012 17282 24064
rect 17405 24055 17463 24061
rect 17405 24021 17417 24055
rect 17451 24052 17463 24055
rect 17494 24052 17500 24064
rect 17451 24024 17500 24052
rect 17451 24021 17463 24024
rect 17405 24015 17463 24021
rect 17494 24012 17500 24024
rect 17552 24012 17558 24064
rect 18693 24055 18751 24061
rect 18693 24021 18705 24055
rect 18739 24052 18751 24055
rect 20088 24052 20116 24083
rect 18739 24024 20116 24052
rect 18739 24021 18751 24024
rect 18693 24015 18751 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 16114 23848 16120 23860
rect 16075 23820 16120 23848
rect 16114 23808 16120 23820
rect 16172 23808 16178 23860
rect 18322 23848 18328 23860
rect 18283 23820 18328 23848
rect 18322 23808 18328 23820
rect 18380 23808 18386 23860
rect 34790 23848 34796 23860
rect 34751 23820 34796 23848
rect 34790 23808 34796 23820
rect 34848 23808 34854 23860
rect 17126 23780 17132 23792
rect 17087 23752 17132 23780
rect 17126 23740 17132 23752
rect 17184 23740 17190 23792
rect 17218 23740 17224 23792
rect 17276 23780 17282 23792
rect 19061 23783 19119 23789
rect 17276 23752 17321 23780
rect 17276 23740 17282 23752
rect 19061 23749 19073 23783
rect 19107 23780 19119 23783
rect 19797 23783 19855 23789
rect 19797 23780 19809 23783
rect 19107 23752 19809 23780
rect 19107 23749 19119 23752
rect 19061 23743 19119 23749
rect 19797 23749 19809 23752
rect 19843 23749 19855 23783
rect 19797 23743 19855 23749
rect 20349 23783 20407 23789
rect 20349 23749 20361 23783
rect 20395 23780 20407 23783
rect 20622 23780 20628 23792
rect 20395 23752 20628 23780
rect 20395 23749 20407 23752
rect 20349 23743 20407 23749
rect 20622 23740 20628 23752
rect 20680 23740 20686 23792
rect 3878 23672 3884 23724
rect 3936 23712 3942 23724
rect 7745 23715 7803 23721
rect 7745 23712 7757 23715
rect 3936 23684 7757 23712
rect 3936 23672 3942 23684
rect 7745 23681 7757 23684
rect 7791 23681 7803 23715
rect 13170 23712 13176 23724
rect 13131 23684 13176 23712
rect 7745 23675 7803 23681
rect 13170 23672 13176 23684
rect 13228 23672 13234 23724
rect 15470 23712 15476 23724
rect 15431 23684 15476 23712
rect 15470 23672 15476 23684
rect 15528 23672 15534 23724
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23712 16359 23715
rect 16942 23712 16948 23724
rect 16347 23684 16948 23712
rect 16347 23681 16359 23684
rect 16301 23675 16359 23681
rect 9490 23604 9496 23656
rect 9548 23644 9554 23656
rect 16316 23644 16344 23675
rect 16942 23672 16948 23684
rect 17000 23672 17006 23724
rect 18506 23712 18512 23724
rect 18467 23684 18512 23712
rect 18506 23672 18512 23684
rect 18564 23712 18570 23724
rect 18969 23715 19027 23721
rect 18969 23712 18981 23715
rect 18564 23684 18981 23712
rect 18564 23672 18570 23684
rect 18969 23681 18981 23684
rect 19015 23681 19027 23715
rect 18969 23675 19027 23681
rect 31754 23672 31760 23724
rect 31812 23712 31818 23724
rect 34977 23715 35035 23721
rect 34977 23712 34989 23715
rect 31812 23684 34989 23712
rect 31812 23672 31818 23684
rect 34977 23681 34989 23684
rect 35023 23681 35035 23715
rect 38286 23712 38292 23724
rect 38247 23684 38292 23712
rect 34977 23675 35035 23681
rect 38286 23672 38292 23684
rect 38344 23672 38350 23724
rect 17402 23644 17408 23656
rect 9548 23616 16344 23644
rect 17363 23616 17408 23644
rect 9548 23604 9554 23616
rect 17402 23604 17408 23616
rect 17460 23604 17466 23656
rect 19426 23604 19432 23656
rect 19484 23644 19490 23656
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 19484 23616 19717 23644
rect 19484 23604 19490 23616
rect 19705 23613 19717 23616
rect 19751 23613 19763 23647
rect 19705 23607 19763 23613
rect 7837 23511 7895 23517
rect 7837 23477 7849 23511
rect 7883 23508 7895 23511
rect 9582 23508 9588 23520
rect 7883 23480 9588 23508
rect 7883 23477 7895 23480
rect 7837 23471 7895 23477
rect 9582 23468 9588 23480
rect 9640 23468 9646 23520
rect 12894 23468 12900 23520
rect 12952 23508 12958 23520
rect 12989 23511 13047 23517
rect 12989 23508 13001 23511
rect 12952 23480 13001 23508
rect 12952 23468 12958 23480
rect 12989 23477 13001 23480
rect 13035 23477 13047 23511
rect 12989 23471 13047 23477
rect 15194 23468 15200 23520
rect 15252 23508 15258 23520
rect 15289 23511 15347 23517
rect 15289 23508 15301 23511
rect 15252 23480 15301 23508
rect 15252 23468 15258 23480
rect 15289 23477 15301 23480
rect 15335 23477 15347 23511
rect 15289 23471 15347 23477
rect 34514 23468 34520 23520
rect 34572 23508 34578 23520
rect 38105 23511 38163 23517
rect 38105 23508 38117 23511
rect 34572 23480 38117 23508
rect 34572 23468 34578 23480
rect 38105 23477 38117 23480
rect 38151 23477 38163 23511
rect 38105 23471 38163 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 18046 23304 18052 23316
rect 16868 23276 18052 23304
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 16868 23168 16896 23276
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 19426 23264 19432 23316
rect 19484 23304 19490 23316
rect 19797 23307 19855 23313
rect 19797 23304 19809 23307
rect 19484 23276 19809 23304
rect 19484 23264 19490 23276
rect 19797 23273 19809 23276
rect 19843 23273 19855 23307
rect 19797 23267 19855 23273
rect 17402 23196 17408 23248
rect 17460 23236 17466 23248
rect 17957 23239 18015 23245
rect 17957 23236 17969 23239
rect 17460 23208 17969 23236
rect 17460 23196 17466 23208
rect 17957 23205 17969 23208
rect 18003 23205 18015 23239
rect 17957 23199 18015 23205
rect 18693 23239 18751 23245
rect 18693 23205 18705 23239
rect 18739 23236 18751 23239
rect 21082 23236 21088 23248
rect 18739 23208 19656 23236
rect 18739 23205 18751 23208
rect 18693 23199 18751 23205
rect 19628 23177 19656 23208
rect 19996 23208 21088 23236
rect 19613 23171 19671 23177
rect 9272 23140 16896 23168
rect 9272 23128 9278 23140
rect 11977 23103 12035 23109
rect 11977 23069 11989 23103
rect 12023 23069 12035 23103
rect 12894 23100 12900 23112
rect 12855 23072 12900 23100
rect 11977 23063 12035 23069
rect 11992 23032 12020 23063
rect 12894 23060 12900 23072
rect 12952 23060 12958 23112
rect 13354 23100 13360 23112
rect 13315 23072 13360 23100
rect 13354 23060 13360 23072
rect 13412 23060 13418 23112
rect 14550 23100 14556 23112
rect 14511 23072 14556 23100
rect 14550 23060 14556 23072
rect 14608 23060 14614 23112
rect 15194 23100 15200 23112
rect 15155 23072 15200 23100
rect 15194 23060 15200 23072
rect 15252 23060 15258 23112
rect 15838 23100 15844 23112
rect 15799 23072 15844 23100
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 16868 23109 16896 23140
rect 17236 23140 19564 23168
rect 16853 23103 16911 23109
rect 16853 23069 16865 23103
rect 16899 23069 16911 23103
rect 16853 23063 16911 23069
rect 13170 23032 13176 23044
rect 11992 23004 13176 23032
rect 13170 22992 13176 23004
rect 13228 23032 13234 23044
rect 13998 23032 14004 23044
rect 13228 23004 14004 23032
rect 13228 22992 13234 23004
rect 13998 22992 14004 23004
rect 14056 22992 14062 23044
rect 17236 23032 17264 23140
rect 18877 23103 18935 23109
rect 18877 23069 18889 23103
rect 18923 23069 18935 23103
rect 18877 23063 18935 23069
rect 19429 23103 19487 23109
rect 19429 23069 19441 23103
rect 19475 23069 19487 23103
rect 19536 23100 19564 23140
rect 19613 23137 19625 23171
rect 19659 23137 19671 23171
rect 19613 23131 19671 23137
rect 19996 23100 20024 23208
rect 21082 23196 21088 23208
rect 21140 23196 21146 23248
rect 20714 23168 20720 23180
rect 20675 23140 20720 23168
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 20898 23100 20904 23112
rect 19536 23072 20024 23100
rect 20859 23072 20904 23100
rect 19429 23063 19487 23069
rect 17405 23035 17463 23041
rect 17405 23032 17417 23035
rect 17236 23004 17417 23032
rect 17405 23001 17417 23004
rect 17451 23001 17463 23035
rect 17405 22995 17463 23001
rect 17494 22992 17500 23044
rect 17552 23032 17558 23044
rect 17552 23004 17597 23032
rect 17552 22992 17558 23004
rect 12066 22964 12072 22976
rect 12027 22936 12072 22964
rect 12066 22924 12072 22936
rect 12124 22924 12130 22976
rect 12710 22964 12716 22976
rect 12671 22936 12716 22964
rect 12710 22924 12716 22936
rect 12768 22924 12774 22976
rect 13446 22964 13452 22976
rect 13407 22936 13452 22964
rect 13446 22924 13452 22936
rect 13504 22924 13510 22976
rect 14366 22964 14372 22976
rect 14327 22936 14372 22964
rect 14366 22924 14372 22936
rect 14424 22924 14430 22976
rect 15010 22964 15016 22976
rect 14971 22936 15016 22964
rect 15010 22924 15016 22936
rect 15068 22924 15074 22976
rect 15654 22964 15660 22976
rect 15615 22936 15660 22964
rect 15654 22924 15660 22936
rect 15712 22924 15718 22976
rect 16669 22967 16727 22973
rect 16669 22933 16681 22967
rect 16715 22964 16727 22967
rect 18892 22964 18920 23063
rect 19444 23032 19472 23063
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 21174 23032 21180 23044
rect 19444 23004 21180 23032
rect 21174 22992 21180 23004
rect 21232 22992 21238 23044
rect 16715 22936 18920 22964
rect 16715 22933 16727 22936
rect 16669 22927 16727 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 5442 22760 5448 22772
rect 5403 22732 5448 22760
rect 5442 22720 5448 22732
rect 5500 22720 5506 22772
rect 14550 22760 14556 22772
rect 14108 22732 14556 22760
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 5629 22627 5687 22633
rect 5629 22593 5641 22627
rect 5675 22624 5687 22627
rect 8202 22624 8208 22636
rect 5675 22596 8208 22624
rect 5675 22593 5687 22596
rect 5629 22587 5687 22593
rect 8202 22584 8208 22596
rect 8260 22584 8266 22636
rect 8570 22584 8576 22636
rect 8628 22624 8634 22636
rect 11885 22627 11943 22633
rect 11885 22624 11897 22627
rect 8628 22596 11897 22624
rect 8628 22584 8634 22596
rect 11885 22593 11897 22596
rect 11931 22593 11943 22627
rect 12066 22624 12072 22636
rect 12027 22596 12072 22624
rect 11885 22587 11943 22593
rect 12066 22584 12072 22596
rect 12124 22584 12130 22636
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22624 13599 22627
rect 14108 22624 14136 22732
rect 14550 22720 14556 22732
rect 14608 22720 14614 22772
rect 15010 22720 15016 22772
rect 15068 22760 15074 22772
rect 19889 22763 19947 22769
rect 15068 22732 17080 22760
rect 15068 22720 15074 22732
rect 17052 22701 17080 22732
rect 19889 22729 19901 22763
rect 19935 22760 19947 22763
rect 20898 22760 20904 22772
rect 19935 22732 20904 22760
rect 19935 22729 19947 22732
rect 19889 22723 19947 22729
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 21082 22760 21088 22772
rect 21043 22732 21088 22760
rect 21082 22720 21088 22732
rect 21140 22720 21146 22772
rect 21174 22720 21180 22772
rect 21232 22760 21238 22772
rect 21542 22760 21548 22772
rect 21232 22732 21548 22760
rect 21232 22720 21238 22732
rect 21542 22720 21548 22732
rect 21600 22760 21606 22772
rect 29822 22760 29828 22772
rect 21600 22732 29828 22760
rect 21600 22720 21606 22732
rect 29822 22720 29828 22732
rect 29880 22720 29886 22772
rect 14277 22695 14335 22701
rect 14277 22661 14289 22695
rect 14323 22692 14335 22695
rect 15657 22695 15715 22701
rect 15657 22692 15669 22695
rect 14323 22664 15669 22692
rect 14323 22661 14335 22664
rect 14277 22655 14335 22661
rect 15657 22661 15669 22664
rect 15703 22661 15715 22695
rect 15657 22655 15715 22661
rect 17037 22695 17095 22701
rect 17037 22661 17049 22695
rect 17083 22661 17095 22695
rect 17586 22692 17592 22704
rect 17547 22664 17592 22692
rect 17037 22655 17095 22661
rect 17586 22652 17592 22664
rect 17644 22652 17650 22704
rect 13587 22596 14136 22624
rect 14185 22627 14243 22633
rect 13587 22593 13599 22596
rect 13541 22587 13599 22593
rect 14185 22593 14197 22627
rect 14231 22593 14243 22627
rect 14185 22587 14243 22593
rect 13722 22448 13728 22500
rect 13780 22488 13786 22500
rect 14200 22488 14228 22587
rect 14366 22584 14372 22636
rect 14424 22624 14430 22636
rect 15013 22627 15071 22633
rect 15013 22624 15025 22627
rect 14424 22596 15025 22624
rect 14424 22584 14430 22596
rect 15013 22593 15025 22596
rect 15059 22593 15071 22627
rect 18690 22624 18696 22636
rect 18651 22596 18696 22624
rect 15013 22587 15071 22593
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 19794 22624 19800 22636
rect 19755 22596 19800 22624
rect 19794 22584 19800 22596
rect 19852 22584 19858 22636
rect 20438 22624 20444 22636
rect 20399 22596 20444 22624
rect 20438 22584 20444 22596
rect 20496 22584 20502 22636
rect 15565 22559 15623 22565
rect 15565 22525 15577 22559
rect 15611 22556 15623 22559
rect 15746 22556 15752 22568
rect 15611 22528 15752 22556
rect 15611 22525 15623 22528
rect 15565 22519 15623 22525
rect 15746 22516 15752 22528
rect 15804 22516 15810 22568
rect 16945 22559 17003 22565
rect 16945 22525 16957 22559
rect 16991 22556 17003 22559
rect 18138 22556 18144 22568
rect 16991 22528 18144 22556
rect 16991 22525 17003 22528
rect 16945 22519 17003 22525
rect 18138 22516 18144 22528
rect 18196 22516 18202 22568
rect 18230 22516 18236 22568
rect 18288 22556 18294 22568
rect 19153 22559 19211 22565
rect 19153 22556 19165 22559
rect 18288 22528 19165 22556
rect 18288 22516 18294 22528
rect 19153 22525 19165 22528
rect 19199 22525 19211 22559
rect 20622 22556 20628 22568
rect 20583 22528 20628 22556
rect 19153 22519 19211 22525
rect 20622 22516 20628 22528
rect 20680 22516 20686 22568
rect 15470 22488 15476 22500
rect 13780 22460 15476 22488
rect 13780 22448 13786 22460
rect 15470 22448 15476 22460
rect 15528 22448 15534 22500
rect 16117 22491 16175 22497
rect 16117 22457 16129 22491
rect 16163 22488 16175 22491
rect 17586 22488 17592 22500
rect 16163 22460 17592 22488
rect 16163 22457 16175 22460
rect 16117 22451 16175 22457
rect 17586 22448 17592 22460
rect 17644 22448 17650 22500
rect 1581 22423 1639 22429
rect 1581 22389 1593 22423
rect 1627 22420 1639 22423
rect 5534 22420 5540 22432
rect 1627 22392 5540 22420
rect 1627 22389 1639 22392
rect 1581 22383 1639 22389
rect 5534 22380 5540 22392
rect 5592 22380 5598 22432
rect 12529 22423 12587 22429
rect 12529 22389 12541 22423
rect 12575 22420 12587 22423
rect 13262 22420 13268 22432
rect 12575 22392 13268 22420
rect 12575 22389 12587 22392
rect 12529 22383 12587 22389
rect 13262 22380 13268 22392
rect 13320 22380 13326 22432
rect 13633 22423 13691 22429
rect 13633 22389 13645 22423
rect 13679 22420 13691 22423
rect 14458 22420 14464 22432
rect 13679 22392 14464 22420
rect 13679 22389 13691 22392
rect 13633 22383 13691 22389
rect 14458 22380 14464 22392
rect 14516 22380 14522 22432
rect 14829 22423 14887 22429
rect 14829 22389 14841 22423
rect 14875 22420 14887 22423
rect 16206 22420 16212 22432
rect 14875 22392 16212 22420
rect 14875 22389 14887 22392
rect 14829 22383 14887 22389
rect 16206 22380 16212 22392
rect 16264 22380 16270 22432
rect 18506 22420 18512 22432
rect 18467 22392 18512 22420
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 13262 22216 13268 22228
rect 13223 22188 13268 22216
rect 13262 22176 13268 22188
rect 13320 22176 13326 22228
rect 18138 22176 18144 22228
rect 18196 22216 18202 22228
rect 18598 22216 18604 22228
rect 18196 22188 18604 22216
rect 18196 22176 18202 22188
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 20533 22219 20591 22225
rect 20533 22185 20545 22219
rect 20579 22216 20591 22219
rect 20622 22216 20628 22228
rect 20579 22188 20628 22216
rect 20579 22185 20591 22188
rect 20533 22179 20591 22185
rect 20622 22176 20628 22188
rect 20680 22176 20686 22228
rect 4433 22083 4491 22089
rect 4433 22049 4445 22083
rect 4479 22080 4491 22083
rect 4614 22080 4620 22092
rect 4479 22052 4620 22080
rect 4479 22049 4491 22052
rect 4433 22043 4491 22049
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 8202 22040 8208 22092
rect 8260 22080 8266 22092
rect 12345 22083 12403 22089
rect 12345 22080 12357 22083
rect 8260 22052 12357 22080
rect 8260 22040 8266 22052
rect 12345 22049 12357 22052
rect 12391 22049 12403 22083
rect 12345 22043 12403 22049
rect 12710 22040 12716 22092
rect 12768 22080 12774 22092
rect 13081 22083 13139 22089
rect 13081 22080 13093 22083
rect 12768 22052 13093 22080
rect 12768 22040 12774 22052
rect 13081 22049 13093 22052
rect 13127 22049 13139 22083
rect 13280 22080 13308 22176
rect 13814 22108 13820 22160
rect 13872 22148 13878 22160
rect 19794 22148 19800 22160
rect 13872 22120 19800 22148
rect 13872 22108 13878 22120
rect 19794 22108 19800 22120
rect 19852 22148 19858 22160
rect 19852 22120 21404 22148
rect 19852 22108 19858 22120
rect 14369 22083 14427 22089
rect 14369 22080 14381 22083
rect 13280 22052 14381 22080
rect 13081 22043 13139 22049
rect 14369 22049 14381 22052
rect 14415 22049 14427 22083
rect 14369 22043 14427 22049
rect 15013 22083 15071 22089
rect 15013 22049 15025 22083
rect 15059 22080 15071 22083
rect 16577 22083 16635 22089
rect 16577 22080 16589 22083
rect 15059 22052 16589 22080
rect 15059 22049 15071 22052
rect 15013 22043 15071 22049
rect 16577 22049 16589 22052
rect 16623 22080 16635 22083
rect 16758 22080 16764 22092
rect 16623 22052 16764 22080
rect 16623 22049 16635 22052
rect 16577 22043 16635 22049
rect 16758 22040 16764 22052
rect 16816 22040 16822 22092
rect 18230 22080 18236 22092
rect 18191 22052 18236 22080
rect 18230 22040 18236 22052
rect 18288 22040 18294 22092
rect 18417 22083 18475 22089
rect 18417 22049 18429 22083
rect 18463 22080 18475 22083
rect 18506 22080 18512 22092
rect 18463 22052 18512 22080
rect 18463 22049 18475 22052
rect 18417 22043 18475 22049
rect 18506 22040 18512 22052
rect 18564 22040 18570 22092
rect 4341 22015 4399 22021
rect 4341 21981 4353 22015
rect 4387 22012 4399 22015
rect 4798 22012 4804 22024
rect 4387 21984 4804 22012
rect 4387 21981 4399 21984
rect 4341 21975 4399 21981
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 7834 21972 7840 22024
rect 7892 22012 7898 22024
rect 10045 22015 10103 22021
rect 10045 22012 10057 22015
rect 7892 21984 10057 22012
rect 7892 21972 7898 21984
rect 10045 21981 10057 21984
rect 10091 21981 10103 22015
rect 11146 22012 11152 22024
rect 11107 21984 11152 22012
rect 10045 21975 10103 21981
rect 11146 21972 11152 21984
rect 11204 21972 11210 22024
rect 11514 21972 11520 22024
rect 11572 22012 11578 22024
rect 11793 22015 11851 22021
rect 11793 22012 11805 22015
rect 11572 21984 11805 22012
rect 11572 21972 11578 21984
rect 11793 21981 11805 21984
rect 11839 21981 11851 22015
rect 12250 22012 12256 22024
rect 12211 21984 12256 22012
rect 11793 21975 11851 21981
rect 12250 21972 12256 21984
rect 12308 21972 12314 22024
rect 12897 22015 12955 22021
rect 12897 21981 12909 22015
rect 12943 21981 12955 22015
rect 12897 21975 12955 21981
rect 11238 21904 11244 21956
rect 11296 21944 11302 21956
rect 12912 21944 12940 21975
rect 17678 21972 17684 22024
rect 17736 22012 17742 22024
rect 21376 22021 21404 22120
rect 28353 22083 28411 22089
rect 28353 22049 28365 22083
rect 28399 22080 28411 22083
rect 31754 22080 31760 22092
rect 28399 22052 31760 22080
rect 28399 22049 28411 22052
rect 28353 22043 28411 22049
rect 31754 22040 31760 22052
rect 31812 22040 31818 22092
rect 17773 22015 17831 22021
rect 17773 22012 17785 22015
rect 17736 21984 17785 22012
rect 17736 21972 17742 21984
rect 17773 21981 17785 21984
rect 17819 22012 17831 22015
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 17819 21984 19441 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 20717 22015 20775 22021
rect 20717 21981 20729 22015
rect 20763 21981 20775 22015
rect 20717 21975 20775 21981
rect 21361 22015 21419 22021
rect 21361 21981 21373 22015
rect 21407 21981 21419 22015
rect 21361 21975 21419 21981
rect 11296 21916 12940 21944
rect 11296 21904 11302 21916
rect 10137 21879 10195 21885
rect 10137 21845 10149 21879
rect 10183 21876 10195 21879
rect 10318 21876 10324 21888
rect 10183 21848 10324 21876
rect 10183 21845 10195 21848
rect 10137 21839 10195 21845
rect 10318 21836 10324 21848
rect 10376 21836 10382 21888
rect 10962 21876 10968 21888
rect 10923 21848 10968 21876
rect 10962 21836 10968 21848
rect 11020 21836 11026 21888
rect 11606 21876 11612 21888
rect 11567 21848 11612 21876
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 12912 21876 12940 21916
rect 14458 21904 14464 21956
rect 14516 21944 14522 21956
rect 16114 21944 16120 21956
rect 14516 21916 14561 21944
rect 16075 21916 16120 21944
rect 14516 21904 14522 21916
rect 16114 21904 16120 21916
rect 16172 21904 16178 21956
rect 16206 21904 16212 21956
rect 16264 21944 16270 21956
rect 18782 21944 18788 21956
rect 16264 21916 16309 21944
rect 16408 21916 18788 21944
rect 16264 21904 16270 21916
rect 16408 21876 16436 21916
rect 18782 21904 18788 21916
rect 18840 21904 18846 21956
rect 12912 21848 16436 21876
rect 17589 21879 17647 21885
rect 17589 21845 17601 21879
rect 17635 21876 17647 21879
rect 18690 21876 18696 21888
rect 17635 21848 18696 21876
rect 17635 21845 17647 21848
rect 17589 21839 17647 21845
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 19521 21879 19579 21885
rect 19521 21876 19533 21879
rect 19484 21848 19533 21876
rect 19484 21836 19490 21848
rect 19521 21845 19533 21848
rect 19567 21845 19579 21879
rect 20732 21876 20760 21975
rect 24854 21972 24860 22024
rect 24912 22012 24918 22024
rect 28261 22015 28319 22021
rect 28261 22012 28273 22015
rect 24912 21984 28273 22012
rect 24912 21972 24918 21984
rect 28261 21981 28273 21984
rect 28307 21981 28319 22015
rect 38286 22012 38292 22024
rect 38247 21984 38292 22012
rect 28261 21975 28319 21981
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 21177 21879 21235 21885
rect 21177 21876 21189 21879
rect 20732 21848 21189 21876
rect 19521 21839 19579 21845
rect 21177 21845 21189 21848
rect 21223 21845 21235 21879
rect 38102 21876 38108 21888
rect 38063 21848 38108 21876
rect 21177 21839 21235 21845
rect 38102 21836 38108 21848
rect 38160 21836 38166 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 10321 21675 10379 21681
rect 10321 21641 10333 21675
rect 10367 21672 10379 21675
rect 11146 21672 11152 21684
rect 10367 21644 11152 21672
rect 10367 21641 10379 21644
rect 10321 21635 10379 21641
rect 11146 21632 11152 21644
rect 11204 21632 11210 21684
rect 13354 21632 13360 21684
rect 13412 21632 13418 21684
rect 14921 21675 14979 21681
rect 14921 21641 14933 21675
rect 14967 21672 14979 21675
rect 15838 21672 15844 21684
rect 14967 21644 15844 21672
rect 14967 21641 14979 21644
rect 14921 21635 14979 21641
rect 15838 21632 15844 21644
rect 15896 21632 15902 21684
rect 18598 21632 18604 21684
rect 18656 21672 18662 21684
rect 20165 21675 20223 21681
rect 20165 21672 20177 21675
rect 18656 21644 20177 21672
rect 18656 21632 18662 21644
rect 20165 21641 20177 21644
rect 20211 21641 20223 21675
rect 20165 21635 20223 21641
rect 13372 21604 13400 21632
rect 17678 21604 17684 21616
rect 13372 21576 17684 21604
rect 1581 21539 1639 21545
rect 1581 21505 1593 21539
rect 1627 21536 1639 21539
rect 4890 21536 4896 21548
rect 1627 21508 4896 21536
rect 1627 21505 1639 21508
rect 1581 21499 1639 21505
rect 4890 21496 4896 21508
rect 4948 21496 4954 21548
rect 5074 21536 5080 21548
rect 5035 21508 5080 21536
rect 5074 21496 5080 21508
rect 5132 21496 5138 21548
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21536 8171 21539
rect 9030 21536 9036 21548
rect 8159 21508 9036 21536
rect 8159 21505 8171 21508
rect 8113 21499 8171 21505
rect 9030 21496 9036 21508
rect 9088 21496 9094 21548
rect 9677 21539 9735 21545
rect 9677 21505 9689 21539
rect 9723 21536 9735 21539
rect 10042 21536 10048 21548
rect 9723 21508 10048 21536
rect 9723 21505 9735 21508
rect 9677 21499 9735 21505
rect 10042 21496 10048 21508
rect 10100 21496 10106 21548
rect 10502 21536 10508 21548
rect 10463 21508 10508 21536
rect 10502 21496 10508 21508
rect 10560 21536 10566 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 10560 21508 10977 21536
rect 10560 21496 10566 21508
rect 10965 21505 10977 21508
rect 11011 21505 11023 21539
rect 11698 21536 11704 21548
rect 11659 21508 11704 21536
rect 10965 21499 11023 21505
rect 11698 21496 11704 21508
rect 11756 21496 11762 21548
rect 12158 21496 12164 21548
rect 12216 21536 12222 21548
rect 13173 21539 13231 21545
rect 13173 21536 13185 21539
rect 12216 21508 13185 21536
rect 12216 21496 12222 21508
rect 13173 21505 13185 21508
rect 13219 21505 13231 21539
rect 13173 21499 13231 21505
rect 13357 21539 13415 21545
rect 13357 21505 13369 21539
rect 13403 21536 13415 21539
rect 13446 21536 13452 21548
rect 13403 21508 13452 21536
rect 13403 21505 13415 21508
rect 13357 21499 13415 21505
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 15120 21545 15148 21576
rect 17678 21564 17684 21576
rect 17736 21564 17742 21616
rect 20625 21607 20683 21613
rect 20625 21604 20637 21607
rect 18432 21576 20637 21604
rect 15105 21539 15163 21545
rect 15105 21505 15117 21539
rect 15151 21505 15163 21539
rect 15105 21499 15163 21505
rect 15654 21496 15660 21548
rect 15712 21536 15718 21548
rect 15749 21539 15807 21545
rect 15749 21536 15761 21539
rect 15712 21508 15761 21536
rect 15712 21496 15718 21508
rect 15749 21505 15761 21508
rect 15795 21505 15807 21539
rect 17310 21536 17316 21548
rect 17271 21508 17316 21536
rect 15749 21499 15807 21505
rect 17310 21496 17316 21508
rect 17368 21496 17374 21548
rect 18432 21545 18460 21576
rect 20625 21573 20637 21576
rect 20671 21573 20683 21607
rect 20625 21567 20683 21573
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21505 17831 21539
rect 17773 21499 17831 21505
rect 18417 21539 18475 21545
rect 18417 21505 18429 21539
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 8754 21468 8760 21480
rect 8715 21440 8760 21468
rect 8754 21428 8760 21440
rect 8812 21428 8818 21480
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21468 11115 21471
rect 11885 21471 11943 21477
rect 11885 21468 11897 21471
rect 11103 21440 11897 21468
rect 11103 21437 11115 21440
rect 11057 21431 11115 21437
rect 11885 21437 11897 21440
rect 11931 21437 11943 21471
rect 11885 21431 11943 21437
rect 14277 21471 14335 21477
rect 14277 21437 14289 21471
rect 14323 21468 14335 21471
rect 15470 21468 15476 21480
rect 14323 21440 15476 21468
rect 14323 21437 14335 21440
rect 14277 21431 14335 21437
rect 15470 21428 15476 21440
rect 15528 21428 15534 21480
rect 15562 21428 15568 21480
rect 15620 21468 15626 21480
rect 15620 21440 15665 21468
rect 15620 21428 15626 21440
rect 16942 21428 16948 21480
rect 17000 21468 17006 21480
rect 17788 21468 17816 21499
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19705 21539 19763 21545
rect 19705 21536 19717 21539
rect 19484 21508 19717 21536
rect 19484 21496 19490 21508
rect 19705 21505 19717 21508
rect 19751 21505 19763 21539
rect 19705 21499 19763 21505
rect 31389 21539 31447 21545
rect 31389 21505 31401 21539
rect 31435 21536 31447 21539
rect 34514 21536 34520 21548
rect 31435 21508 34520 21536
rect 31435 21505 31447 21508
rect 31389 21499 31447 21505
rect 34514 21496 34520 21508
rect 34572 21496 34578 21548
rect 34606 21496 34612 21548
rect 34664 21536 34670 21548
rect 34664 21508 34709 21536
rect 34664 21496 34670 21508
rect 17000 21440 17816 21468
rect 18601 21471 18659 21477
rect 17000 21428 17006 21440
rect 18601 21437 18613 21471
rect 18647 21468 18659 21471
rect 18690 21468 18696 21480
rect 18647 21440 18696 21468
rect 18647 21437 18659 21440
rect 18601 21431 18659 21437
rect 18690 21428 18696 21440
rect 18748 21428 18754 21480
rect 19521 21471 19579 21477
rect 19521 21437 19533 21471
rect 19567 21468 19579 21471
rect 19978 21468 19984 21480
rect 19567 21440 19984 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 19978 21428 19984 21440
rect 20036 21468 20042 21480
rect 20438 21468 20444 21480
rect 20036 21440 20444 21468
rect 20036 21428 20042 21440
rect 20438 21428 20444 21440
rect 20496 21428 20502 21480
rect 22554 21468 22560 21480
rect 22515 21440 22560 21468
rect 22554 21428 22560 21440
rect 22612 21428 22618 21480
rect 5169 21403 5227 21409
rect 5169 21369 5181 21403
rect 5215 21400 5227 21403
rect 6270 21400 6276 21412
rect 5215 21372 6276 21400
rect 5215 21369 5227 21372
rect 5169 21363 5227 21369
rect 6270 21360 6276 21372
rect 6328 21360 6334 21412
rect 8018 21360 8024 21412
rect 8076 21400 8082 21412
rect 13722 21400 13728 21412
rect 8076 21372 13728 21400
rect 8076 21360 8082 21372
rect 13722 21360 13728 21372
rect 13780 21360 13786 21412
rect 13817 21403 13875 21409
rect 13817 21369 13829 21403
rect 13863 21400 13875 21403
rect 15746 21400 15752 21412
rect 13863 21372 15752 21400
rect 13863 21369 13875 21372
rect 13817 21363 13875 21369
rect 15746 21360 15752 21372
rect 15804 21400 15810 21412
rect 15933 21403 15991 21409
rect 15933 21400 15945 21403
rect 15804 21372 15945 21400
rect 15804 21360 15810 21372
rect 15933 21369 15945 21372
rect 15979 21369 15991 21403
rect 15933 21363 15991 21369
rect 17034 21360 17040 21412
rect 17092 21400 17098 21412
rect 18785 21403 18843 21409
rect 18785 21400 18797 21403
rect 17092 21372 18797 21400
rect 17092 21360 17098 21372
rect 18785 21369 18797 21372
rect 18831 21400 18843 21403
rect 19794 21400 19800 21412
rect 18831 21372 19800 21400
rect 18831 21369 18843 21372
rect 18785 21363 18843 21369
rect 19794 21360 19800 21372
rect 19852 21360 19858 21412
rect 1762 21332 1768 21344
rect 1723 21304 1768 21332
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 5534 21292 5540 21344
rect 5592 21332 5598 21344
rect 8205 21335 8263 21341
rect 8205 21332 8217 21335
rect 5592 21304 8217 21332
rect 5592 21292 5598 21304
rect 8205 21301 8217 21304
rect 8251 21301 8263 21335
rect 9766 21332 9772 21344
rect 9727 21304 9772 21332
rect 8205 21295 8263 21301
rect 9766 21292 9772 21304
rect 9824 21292 9830 21344
rect 12066 21332 12072 21344
rect 12027 21304 12072 21332
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 17126 21332 17132 21344
rect 17087 21304 17132 21332
rect 17126 21292 17132 21304
rect 17184 21292 17190 21344
rect 17862 21332 17868 21344
rect 17823 21304 17868 21332
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 31481 21335 31539 21341
rect 31481 21332 31493 21335
rect 20956 21304 31493 21332
rect 20956 21292 20962 21304
rect 31481 21301 31493 21304
rect 31527 21301 31539 21335
rect 34698 21332 34704 21344
rect 34659 21304 34704 21332
rect 31481 21295 31539 21301
rect 34698 21292 34704 21304
rect 34756 21292 34762 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 6362 21088 6368 21140
rect 6420 21128 6426 21140
rect 6420 21100 8708 21128
rect 6420 21088 6426 21100
rect 7745 21063 7803 21069
rect 7745 21029 7757 21063
rect 7791 21029 7803 21063
rect 7745 21023 7803 21029
rect 7760 20992 7788 21023
rect 7760 20964 8616 20992
rect 8588 20933 8616 20964
rect 7929 20927 7987 20933
rect 7929 20893 7941 20927
rect 7975 20893 7987 20927
rect 7929 20887 7987 20893
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20893 8631 20927
rect 8680 20924 8708 21100
rect 9030 21088 9036 21140
rect 9088 21128 9094 21140
rect 9953 21131 10011 21137
rect 9953 21128 9965 21131
rect 9088 21100 9965 21128
rect 9088 21088 9094 21100
rect 9953 21097 9965 21100
rect 9999 21097 10011 21131
rect 9953 21091 10011 21097
rect 12250 21088 12256 21140
rect 12308 21128 12314 21140
rect 15194 21128 15200 21140
rect 12308 21100 15200 21128
rect 12308 21088 12314 21100
rect 15194 21088 15200 21100
rect 15252 21088 15258 21140
rect 16114 21128 16120 21140
rect 16075 21100 16120 21128
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 18690 21128 18696 21140
rect 18651 21100 18696 21128
rect 18690 21088 18696 21100
rect 18748 21088 18754 21140
rect 19794 21128 19800 21140
rect 19755 21100 19800 21128
rect 19794 21088 19800 21100
rect 19852 21088 19858 21140
rect 28905 21131 28963 21137
rect 28905 21097 28917 21131
rect 28951 21128 28963 21131
rect 32030 21128 32036 21140
rect 28951 21100 32036 21128
rect 28951 21097 28963 21100
rect 28905 21091 28963 21097
rect 32030 21088 32036 21100
rect 32088 21088 32094 21140
rect 11609 21063 11667 21069
rect 11609 21060 11621 21063
rect 9600 21032 11621 21060
rect 9600 21001 9628 21032
rect 11609 21029 11621 21032
rect 11655 21060 11667 21063
rect 12066 21060 12072 21072
rect 11655 21032 12072 21060
rect 11655 21029 11667 21032
rect 11609 21023 11667 21029
rect 12066 21020 12072 21032
rect 12124 21020 12130 21072
rect 17862 21020 17868 21072
rect 17920 21060 17926 21072
rect 17920 21032 19656 21060
rect 17920 21020 17926 21032
rect 9585 20995 9643 21001
rect 9585 20961 9597 20995
rect 9631 20961 9643 20995
rect 9766 20992 9772 21004
rect 9727 20964 9772 20992
rect 9585 20955 9643 20961
rect 9766 20952 9772 20964
rect 9824 20952 9830 21004
rect 10962 20952 10968 21004
rect 11020 20992 11026 21004
rect 11425 20995 11483 21001
rect 11425 20992 11437 20995
rect 11020 20964 11437 20992
rect 11020 20952 11026 20964
rect 11425 20961 11437 20964
rect 11471 20961 11483 20995
rect 11425 20955 11483 20961
rect 12989 20995 13047 21001
rect 12989 20961 13001 20995
rect 13035 20992 13047 20995
rect 14829 20995 14887 21001
rect 14829 20992 14841 20995
rect 13035 20964 14841 20992
rect 13035 20961 13047 20964
rect 12989 20955 13047 20961
rect 14829 20961 14841 20964
rect 14875 20961 14887 20995
rect 14829 20955 14887 20961
rect 16945 20995 17003 21001
rect 16945 20961 16957 20995
rect 16991 20992 17003 20995
rect 17681 20995 17739 21001
rect 17681 20992 17693 20995
rect 16991 20964 17693 20992
rect 16991 20961 17003 20964
rect 16945 20955 17003 20961
rect 17681 20961 17693 20964
rect 17727 20961 17739 20995
rect 17681 20955 17739 20961
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 19628 21001 19656 21032
rect 19429 20995 19487 21001
rect 19429 20992 19441 20995
rect 19392 20964 19441 20992
rect 19392 20952 19398 20964
rect 19429 20961 19441 20964
rect 19475 20961 19487 20995
rect 19429 20955 19487 20961
rect 19613 20995 19671 21001
rect 19613 20961 19625 20995
rect 19659 20961 19671 20995
rect 22554 20992 22560 21004
rect 22515 20964 22560 20992
rect 19613 20955 19671 20961
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 23198 20992 23204 21004
rect 23159 20964 23204 20992
rect 23198 20952 23204 20964
rect 23256 20952 23262 21004
rect 11238 20924 11244 20936
rect 8680 20896 10180 20924
rect 11199 20896 11244 20924
rect 8573 20887 8631 20893
rect 7944 20856 7972 20887
rect 10042 20856 10048 20868
rect 7944 20828 10048 20856
rect 10042 20816 10048 20828
rect 10100 20816 10106 20868
rect 10152 20856 10180 20896
rect 11238 20884 11244 20896
rect 11296 20884 11302 20936
rect 12897 20927 12955 20933
rect 12897 20924 12909 20927
rect 12406 20896 12909 20924
rect 12406 20856 12434 20896
rect 12897 20893 12909 20896
rect 12943 20893 12955 20927
rect 12897 20887 12955 20893
rect 13725 20927 13783 20933
rect 13725 20893 13737 20927
rect 13771 20924 13783 20927
rect 14458 20924 14464 20936
rect 13771 20896 14464 20924
rect 13771 20893 13783 20896
rect 13725 20887 13783 20893
rect 10152 20828 12434 20856
rect 12912 20856 12940 20887
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 14645 20927 14703 20933
rect 14645 20893 14657 20927
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 13814 20856 13820 20868
rect 12912 20828 13820 20856
rect 13814 20816 13820 20828
rect 13872 20816 13878 20868
rect 14660 20856 14688 20887
rect 15562 20884 15568 20936
rect 15620 20924 15626 20936
rect 15749 20927 15807 20933
rect 15749 20924 15761 20927
rect 15620 20896 15761 20924
rect 15620 20884 15626 20896
rect 15749 20893 15761 20896
rect 15795 20893 15807 20927
rect 15930 20924 15936 20936
rect 15891 20896 15936 20924
rect 15749 20887 15807 20893
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 16850 20924 16856 20936
rect 16811 20896 16856 20924
rect 16850 20884 16856 20896
rect 16908 20884 16914 20936
rect 17497 20927 17555 20933
rect 17497 20893 17509 20927
rect 17543 20924 17555 20927
rect 18230 20924 18236 20936
rect 17543 20896 18236 20924
rect 17543 20893 17555 20896
rect 17497 20887 17555 20893
rect 18230 20884 18236 20896
rect 18288 20924 18294 20936
rect 18414 20924 18420 20936
rect 18288 20896 18420 20924
rect 18288 20884 18294 20896
rect 18414 20884 18420 20896
rect 18472 20884 18478 20936
rect 18874 20924 18880 20936
rect 18835 20896 18880 20924
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 20533 20927 20591 20933
rect 20533 20893 20545 20927
rect 20579 20893 20591 20927
rect 20533 20887 20591 20893
rect 22005 20927 22063 20933
rect 22005 20893 22017 20927
rect 22051 20924 22063 20927
rect 22370 20924 22376 20936
rect 22051 20896 22376 20924
rect 22051 20893 22063 20896
rect 22005 20887 22063 20893
rect 18046 20856 18052 20868
rect 14660 20828 18052 20856
rect 18046 20816 18052 20828
rect 18104 20856 18110 20868
rect 18141 20859 18199 20865
rect 18141 20856 18153 20859
rect 18104 20828 18153 20856
rect 18104 20816 18110 20828
rect 18141 20825 18153 20828
rect 18187 20825 18199 20859
rect 18141 20819 18199 20825
rect 19334 20816 19340 20868
rect 19392 20856 19398 20868
rect 20548 20856 20576 20887
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 28810 20924 28816 20936
rect 28771 20896 28816 20924
rect 28810 20884 28816 20896
rect 28868 20884 28874 20936
rect 22649 20859 22707 20865
rect 22649 20856 22661 20859
rect 19392 20828 20576 20856
rect 22066 20828 22661 20856
rect 19392 20816 19398 20828
rect 8389 20791 8447 20797
rect 8389 20757 8401 20791
rect 8435 20788 8447 20791
rect 8938 20788 8944 20800
rect 8435 20760 8944 20788
rect 8435 20757 8447 20760
rect 8389 20751 8447 20757
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 13541 20791 13599 20797
rect 13541 20757 13553 20791
rect 13587 20788 13599 20791
rect 15102 20788 15108 20800
rect 13587 20760 15108 20788
rect 13587 20757 13599 20760
rect 13541 20751 13599 20757
rect 15102 20748 15108 20760
rect 15160 20748 15166 20800
rect 20622 20788 20628 20800
rect 20583 20760 20628 20788
rect 20622 20748 20628 20760
rect 20680 20748 20686 20800
rect 21821 20791 21879 20797
rect 21821 20757 21833 20791
rect 21867 20788 21879 20791
rect 22066 20788 22094 20828
rect 22649 20825 22661 20828
rect 22695 20825 22707 20859
rect 22649 20819 22707 20825
rect 21867 20760 22094 20788
rect 21867 20757 21879 20760
rect 21821 20751 21879 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 4890 20544 4896 20596
rect 4948 20584 4954 20596
rect 5261 20587 5319 20593
rect 5261 20584 5273 20587
rect 4948 20556 5273 20584
rect 4948 20544 4954 20556
rect 5261 20553 5273 20556
rect 5307 20553 5319 20587
rect 5261 20547 5319 20553
rect 5810 20544 5816 20596
rect 5868 20584 5874 20596
rect 14461 20587 14519 20593
rect 5868 20556 12434 20584
rect 5868 20544 5874 20556
rect 9582 20476 9588 20528
rect 9640 20516 9646 20528
rect 12406 20516 12434 20556
rect 14461 20553 14473 20587
rect 14507 20584 14519 20587
rect 15930 20584 15936 20596
rect 14507 20556 15936 20584
rect 14507 20553 14519 20556
rect 14461 20547 14519 20553
rect 15930 20544 15936 20556
rect 15988 20544 15994 20596
rect 18046 20584 18052 20596
rect 18007 20556 18052 20584
rect 18046 20544 18052 20556
rect 18104 20544 18110 20596
rect 18785 20587 18843 20593
rect 18785 20553 18797 20587
rect 18831 20584 18843 20587
rect 18874 20584 18880 20596
rect 18831 20556 18880 20584
rect 18831 20553 18843 20556
rect 18785 20547 18843 20553
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 21818 20584 21824 20596
rect 19536 20556 21824 20584
rect 9640 20488 12020 20516
rect 12406 20488 15056 20516
rect 9640 20476 9646 20488
rect 5445 20451 5503 20457
rect 5445 20417 5457 20451
rect 5491 20448 5503 20451
rect 5534 20448 5540 20460
rect 5491 20420 5540 20448
rect 5491 20417 5503 20420
rect 5445 20411 5503 20417
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 8754 20448 8760 20460
rect 8715 20420 8760 20448
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 8938 20448 8944 20460
rect 8899 20420 8944 20448
rect 8938 20408 8944 20420
rect 8996 20408 9002 20460
rect 10134 20448 10140 20460
rect 10095 20420 10140 20448
rect 10134 20408 10140 20420
rect 10192 20408 10198 20460
rect 10318 20448 10324 20460
rect 10279 20420 10324 20448
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 11606 20408 11612 20460
rect 11664 20448 11670 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11664 20420 11897 20448
rect 11664 20408 11670 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 11992 20448 12020 20488
rect 15028 20460 15056 20488
rect 16942 20476 16948 20528
rect 17000 20516 17006 20528
rect 17000 20488 19012 20516
rect 17000 20476 17006 20488
rect 12345 20451 12403 20457
rect 12345 20448 12357 20451
rect 11992 20420 12357 20448
rect 11885 20411 11943 20417
rect 12345 20417 12357 20420
rect 12391 20417 12403 20451
rect 13906 20448 13912 20460
rect 13867 20420 13912 20448
rect 12345 20411 12403 20417
rect 13906 20408 13912 20420
rect 13964 20408 13970 20460
rect 13998 20408 14004 20460
rect 14056 20448 14062 20460
rect 14366 20448 14372 20460
rect 14056 20420 14372 20448
rect 14056 20408 14062 20420
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 15010 20448 15016 20460
rect 14923 20420 15016 20448
rect 15010 20408 15016 20420
rect 15068 20408 15074 20460
rect 15102 20408 15108 20460
rect 15160 20448 15166 20460
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15160 20420 15853 20448
rect 15160 20408 15166 20420
rect 15841 20417 15853 20420
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 18984 20457 19012 20488
rect 19536 20457 19564 20556
rect 21818 20544 21824 20556
rect 21876 20544 21882 20596
rect 22370 20544 22376 20596
rect 22428 20584 22434 20596
rect 23569 20587 23627 20593
rect 23569 20584 23581 20587
rect 22428 20556 23581 20584
rect 22428 20544 22434 20556
rect 23569 20553 23581 20556
rect 23615 20553 23627 20587
rect 23569 20547 23627 20553
rect 20806 20516 20812 20528
rect 20767 20488 20812 20516
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 24213 20519 24271 20525
rect 24213 20516 24225 20519
rect 22480 20488 24225 20516
rect 22480 20457 22508 20488
rect 24213 20485 24225 20488
rect 24259 20485 24271 20519
rect 24213 20479 24271 20485
rect 17589 20451 17647 20457
rect 17589 20448 17601 20451
rect 17184 20420 17601 20448
rect 17184 20408 17190 20420
rect 17589 20417 17601 20420
rect 17635 20417 17647 20451
rect 17589 20411 17647 20417
rect 18969 20451 19027 20457
rect 18969 20417 18981 20451
rect 19015 20417 19027 20451
rect 18969 20411 19027 20417
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 22465 20451 22523 20457
rect 22465 20417 22477 20451
rect 22511 20417 22523 20451
rect 23753 20451 23811 20457
rect 23753 20448 23765 20451
rect 22465 20411 22523 20417
rect 22572 20420 23765 20448
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 9858 20380 9864 20392
rect 8159 20352 9864 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 12529 20383 12587 20389
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 15657 20383 15715 20389
rect 15657 20349 15669 20383
rect 15703 20380 15715 20383
rect 17034 20380 17040 20392
rect 15703 20352 17040 20380
rect 15703 20349 15715 20352
rect 15657 20343 15715 20349
rect 9030 20272 9036 20324
rect 9088 20312 9094 20324
rect 9125 20315 9183 20321
rect 9125 20312 9137 20315
rect 9088 20284 9137 20312
rect 9088 20272 9094 20284
rect 9125 20281 9137 20284
rect 9171 20281 9183 20315
rect 9125 20275 9183 20281
rect 11701 20315 11759 20321
rect 11701 20281 11713 20315
rect 11747 20312 11759 20315
rect 12544 20312 12572 20343
rect 17034 20340 17040 20352
rect 17092 20340 17098 20392
rect 17405 20383 17463 20389
rect 17405 20349 17417 20383
rect 17451 20349 17463 20383
rect 17405 20343 17463 20349
rect 19705 20383 19763 20389
rect 19705 20349 19717 20383
rect 19751 20349 19763 20383
rect 19705 20343 19763 20349
rect 11747 20284 12572 20312
rect 12989 20315 13047 20321
rect 11747 20281 11759 20284
rect 11701 20275 11759 20281
rect 12989 20281 13001 20315
rect 13035 20312 13047 20315
rect 14918 20312 14924 20324
rect 13035 20284 14924 20312
rect 13035 20281 13047 20284
rect 12989 20275 13047 20281
rect 14918 20272 14924 20284
rect 14976 20272 14982 20324
rect 15105 20315 15163 20321
rect 15105 20281 15117 20315
rect 15151 20312 15163 20315
rect 17218 20312 17224 20324
rect 15151 20284 17224 20312
rect 15151 20281 15163 20284
rect 15105 20275 15163 20281
rect 17218 20272 17224 20284
rect 17276 20272 17282 20324
rect 10594 20244 10600 20256
rect 10555 20216 10600 20244
rect 10594 20204 10600 20216
rect 10652 20204 10658 20256
rect 13722 20244 13728 20256
rect 13683 20216 13728 20244
rect 13722 20204 13728 20216
rect 13780 20204 13786 20256
rect 15194 20204 15200 20256
rect 15252 20244 15258 20256
rect 16025 20247 16083 20253
rect 16025 20244 16037 20247
rect 15252 20216 16037 20244
rect 15252 20204 15258 20216
rect 16025 20213 16037 20216
rect 16071 20213 16083 20247
rect 16025 20207 16083 20213
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 17420 20244 17448 20343
rect 17494 20272 17500 20324
rect 17552 20312 17558 20324
rect 19720 20312 19748 20343
rect 19978 20340 19984 20392
rect 20036 20380 20042 20392
rect 20717 20383 20775 20389
rect 20717 20380 20729 20383
rect 20036 20352 20729 20380
rect 20036 20340 20042 20352
rect 20717 20349 20729 20352
rect 20763 20349 20775 20383
rect 20717 20343 20775 20349
rect 21361 20383 21419 20389
rect 21361 20349 21373 20383
rect 21407 20380 21419 20383
rect 21818 20380 21824 20392
rect 21407 20352 21824 20380
rect 21407 20349 21419 20352
rect 21361 20343 21419 20349
rect 21818 20340 21824 20352
rect 21876 20340 21882 20392
rect 22002 20340 22008 20392
rect 22060 20380 22066 20392
rect 22572 20380 22600 20420
rect 23753 20417 23765 20420
rect 23799 20417 23811 20451
rect 23753 20411 23811 20417
rect 22060 20352 22600 20380
rect 22649 20383 22707 20389
rect 22060 20340 22066 20352
rect 22649 20349 22661 20383
rect 22695 20380 22707 20383
rect 24578 20380 24584 20392
rect 22695 20352 24584 20380
rect 22695 20349 22707 20352
rect 22649 20343 22707 20349
rect 24578 20340 24584 20352
rect 24636 20340 24642 20392
rect 25222 20312 25228 20324
rect 17552 20284 19748 20312
rect 19812 20284 25228 20312
rect 17552 20272 17558 20284
rect 19812 20244 19840 20284
rect 25222 20272 25228 20284
rect 25280 20272 25286 20324
rect 16632 20216 19840 20244
rect 20165 20247 20223 20253
rect 16632 20204 16638 20216
rect 20165 20213 20177 20247
rect 20211 20244 20223 20247
rect 20254 20244 20260 20256
rect 20211 20216 20260 20244
rect 20211 20213 20223 20216
rect 20165 20207 20223 20213
rect 20254 20204 20260 20216
rect 20312 20204 20318 20256
rect 22830 20244 22836 20256
rect 22791 20216 22836 20244
rect 22830 20204 22836 20216
rect 22888 20204 22894 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 10502 20040 10508 20052
rect 7064 20012 10508 20040
rect 7064 20000 7070 20012
rect 10502 20000 10508 20012
rect 10560 20000 10566 20052
rect 10965 20043 11023 20049
rect 10965 20009 10977 20043
rect 11011 20040 11023 20043
rect 12986 20040 12992 20052
rect 11011 20012 12992 20040
rect 11011 20009 11023 20012
rect 10965 20003 11023 20009
rect 12986 20000 12992 20012
rect 13044 20000 13050 20052
rect 14458 20040 14464 20052
rect 14419 20012 14464 20040
rect 14458 20000 14464 20012
rect 14516 20000 14522 20052
rect 16114 20040 16120 20052
rect 16075 20012 16120 20040
rect 16114 20000 16120 20012
rect 16172 20000 16178 20052
rect 22189 20043 22247 20049
rect 17696 20012 20116 20040
rect 8389 19975 8447 19981
rect 8389 19941 8401 19975
rect 8435 19941 8447 19975
rect 8389 19935 8447 19941
rect 9217 19975 9275 19981
rect 9217 19941 9229 19975
rect 9263 19972 9275 19975
rect 9263 19944 11192 19972
rect 9263 19941 9275 19944
rect 9217 19935 9275 19941
rect 8404 19904 8432 19935
rect 10045 19907 10103 19913
rect 10045 19904 10057 19907
rect 8404 19876 10057 19904
rect 10045 19873 10057 19876
rect 10091 19873 10103 19907
rect 10045 19867 10103 19873
rect 1762 19836 1768 19848
rect 1723 19808 1768 19836
rect 1762 19796 1768 19808
rect 1820 19796 1826 19848
rect 7834 19796 7840 19848
rect 7892 19836 7898 19848
rect 7929 19839 7987 19845
rect 7929 19836 7941 19839
rect 7892 19808 7941 19836
rect 7892 19796 7898 19808
rect 7929 19805 7941 19808
rect 7975 19805 7987 19839
rect 7929 19799 7987 19805
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19805 8631 19839
rect 8573 19799 8631 19805
rect 8588 19768 8616 19799
rect 9214 19796 9220 19848
rect 9272 19836 9278 19848
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 9272 19808 9413 19836
rect 9272 19796 9278 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9858 19836 9864 19848
rect 9819 19808 9864 19836
rect 9401 19799 9459 19805
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 11164 19845 11192 19944
rect 13262 19932 13268 19984
rect 13320 19972 13326 19984
rect 17696 19981 17724 20012
rect 20088 19981 20116 20012
rect 22189 20009 22201 20043
rect 22235 20040 22247 20043
rect 22830 20040 22836 20052
rect 22235 20012 22836 20040
rect 22235 20009 22247 20012
rect 22189 20003 22247 20009
rect 22830 20000 22836 20012
rect 22888 20000 22894 20052
rect 24578 20040 24584 20052
rect 24539 20012 24584 20040
rect 24578 20000 24584 20012
rect 24636 20000 24642 20052
rect 17681 19975 17739 19981
rect 13320 19944 17632 19972
rect 13320 19932 13326 19944
rect 13722 19864 13728 19916
rect 13780 19904 13786 19916
rect 15933 19907 15991 19913
rect 15933 19904 15945 19907
rect 13780 19876 15945 19904
rect 13780 19864 13786 19876
rect 15933 19873 15945 19876
rect 15979 19873 15991 19907
rect 17604 19904 17632 19944
rect 17681 19941 17693 19975
rect 17727 19941 17739 19975
rect 17681 19935 17739 19941
rect 18693 19975 18751 19981
rect 18693 19941 18705 19975
rect 18739 19941 18751 19975
rect 18693 19935 18751 19941
rect 20073 19975 20131 19981
rect 20073 19941 20085 19975
rect 20119 19972 20131 19975
rect 23937 19975 23995 19981
rect 23937 19972 23949 19975
rect 20119 19944 20944 19972
rect 20119 19941 20131 19944
rect 20073 19935 20131 19941
rect 18708 19904 18736 19935
rect 17604 19876 17816 19904
rect 18708 19876 20852 19904
rect 15933 19867 15991 19873
rect 11149 19839 11207 19845
rect 11149 19805 11161 19839
rect 11195 19805 11207 19839
rect 11149 19799 11207 19805
rect 11514 19796 11520 19848
rect 11572 19836 11578 19848
rect 11609 19839 11667 19845
rect 11609 19836 11621 19839
rect 11572 19808 11621 19836
rect 11572 19796 11578 19808
rect 11609 19805 11621 19808
rect 11655 19805 11667 19839
rect 11609 19799 11667 19805
rect 11790 19796 11796 19848
rect 11848 19836 11854 19848
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 11848 19808 12449 19836
rect 11848 19796 11854 19808
rect 12437 19805 12449 19808
rect 12483 19805 12495 19839
rect 12437 19799 12495 19805
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 14645 19839 14703 19845
rect 14645 19836 14657 19839
rect 13872 19808 14657 19836
rect 13872 19796 13878 19808
rect 14645 19805 14657 19808
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 15010 19796 15016 19848
rect 15068 19836 15074 19848
rect 15289 19839 15347 19845
rect 15289 19836 15301 19839
rect 15068 19808 15301 19836
rect 15068 19796 15074 19808
rect 15289 19805 15301 19808
rect 15335 19805 15347 19839
rect 15289 19799 15347 19805
rect 15470 19796 15476 19848
rect 15528 19836 15534 19848
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 15528 19808 15761 19836
rect 15528 19796 15534 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 17788 19836 17816 19876
rect 18877 19839 18935 19845
rect 18877 19836 18889 19839
rect 17788 19808 18889 19836
rect 15749 19799 15807 19805
rect 18877 19805 18889 19808
rect 18923 19836 18935 19839
rect 19334 19836 19340 19848
rect 18923 19808 19340 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 20824 19845 20852 19876
rect 20809 19839 20867 19845
rect 20809 19805 20821 19839
rect 20855 19805 20867 19839
rect 20809 19799 20867 19805
rect 7760 19740 8616 19768
rect 11701 19771 11759 19777
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 5534 19700 5540 19712
rect 1627 19672 5540 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 7760 19709 7788 19740
rect 11701 19737 11713 19771
rect 11747 19768 11759 19771
rect 12802 19768 12808 19780
rect 11747 19740 12808 19768
rect 11747 19737 11759 19740
rect 11701 19731 11759 19737
rect 12802 19728 12808 19740
rect 12860 19728 12866 19780
rect 12897 19771 12955 19777
rect 12897 19737 12909 19771
rect 12943 19768 12955 19771
rect 14274 19768 14280 19780
rect 12943 19740 14280 19768
rect 12943 19737 12955 19740
rect 12897 19731 12955 19737
rect 14274 19728 14280 19740
rect 14332 19728 14338 19780
rect 15378 19768 15384 19780
rect 14936 19740 15384 19768
rect 7745 19703 7803 19709
rect 7745 19669 7757 19703
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 7926 19660 7932 19712
rect 7984 19700 7990 19712
rect 10505 19703 10563 19709
rect 10505 19700 10517 19703
rect 7984 19672 10517 19700
rect 7984 19660 7990 19672
rect 10505 19669 10517 19672
rect 10551 19700 10563 19703
rect 10594 19700 10600 19712
rect 10551 19672 10600 19700
rect 10551 19669 10563 19672
rect 10505 19663 10563 19669
rect 10594 19660 10600 19672
rect 10652 19660 10658 19712
rect 12253 19703 12311 19709
rect 12253 19669 12265 19703
rect 12299 19700 12311 19703
rect 13446 19700 13452 19712
rect 12299 19672 13452 19700
rect 12299 19669 12311 19672
rect 12253 19663 12311 19669
rect 13446 19660 13452 19672
rect 13504 19660 13510 19712
rect 13541 19703 13599 19709
rect 13541 19669 13553 19703
rect 13587 19700 13599 19703
rect 14936 19700 14964 19740
rect 15378 19728 15384 19740
rect 15436 19728 15442 19780
rect 16666 19728 16672 19780
rect 16724 19768 16730 19780
rect 17129 19771 17187 19777
rect 17129 19768 17141 19771
rect 16724 19740 17141 19768
rect 16724 19728 16730 19740
rect 17129 19737 17141 19740
rect 17175 19737 17187 19771
rect 17129 19731 17187 19737
rect 17218 19728 17224 19780
rect 17276 19768 17282 19780
rect 17276 19740 17321 19768
rect 17276 19728 17282 19740
rect 18138 19728 18144 19780
rect 18196 19768 18202 19780
rect 19521 19771 19579 19777
rect 19521 19768 19533 19771
rect 18196 19740 19533 19768
rect 18196 19728 18202 19740
rect 19521 19737 19533 19740
rect 19567 19737 19579 19771
rect 19521 19731 19579 19737
rect 19613 19771 19671 19777
rect 19613 19737 19625 19771
rect 19659 19737 19671 19771
rect 19613 19731 19671 19737
rect 13587 19672 14964 19700
rect 15105 19703 15163 19709
rect 13587 19669 13599 19672
rect 13541 19663 13599 19669
rect 15105 19669 15117 19703
rect 15151 19700 15163 19703
rect 16758 19700 16764 19712
rect 15151 19672 16764 19700
rect 15151 19669 15163 19672
rect 15105 19663 15163 19669
rect 16758 19660 16764 19672
rect 16816 19660 16822 19712
rect 16850 19660 16856 19712
rect 16908 19700 16914 19712
rect 19628 19700 19656 19731
rect 16908 19672 19656 19700
rect 16908 19660 16914 19672
rect 20070 19660 20076 19712
rect 20128 19700 20134 19712
rect 20625 19703 20683 19709
rect 20625 19700 20637 19703
rect 20128 19672 20637 19700
rect 20128 19660 20134 19672
rect 20625 19669 20637 19672
rect 20671 19669 20683 19703
rect 20916 19700 20944 19944
rect 22066 19944 23949 19972
rect 21729 19907 21787 19913
rect 21729 19873 21741 19907
rect 21775 19904 21787 19907
rect 22066 19904 22094 19944
rect 23937 19941 23949 19944
rect 23983 19941 23995 19975
rect 23937 19935 23995 19941
rect 23198 19904 23204 19916
rect 21775 19876 22094 19904
rect 23159 19876 23204 19904
rect 21775 19873 21787 19876
rect 21729 19867 21787 19873
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 21542 19836 21548 19848
rect 21503 19808 21548 19836
rect 21542 19796 21548 19808
rect 21600 19796 21606 19848
rect 23842 19836 23848 19848
rect 23803 19808 23848 19836
rect 23842 19796 23848 19808
rect 23900 19796 23906 19848
rect 24762 19836 24768 19848
rect 24723 19808 24768 19836
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 25406 19836 25412 19848
rect 25367 19808 25412 19836
rect 25406 19796 25412 19808
rect 25464 19796 25470 19848
rect 38286 19836 38292 19848
rect 38247 19808 38292 19836
rect 38286 19796 38292 19808
rect 38344 19796 38350 19848
rect 22738 19768 22744 19780
rect 22699 19740 22744 19768
rect 22738 19728 22744 19740
rect 22796 19728 22802 19780
rect 22830 19728 22836 19780
rect 22888 19768 22894 19780
rect 22888 19740 22933 19768
rect 22888 19728 22894 19740
rect 24854 19700 24860 19712
rect 20916 19672 24860 19700
rect 20625 19663 20683 19669
rect 24854 19660 24860 19672
rect 24912 19660 24918 19712
rect 25222 19700 25228 19712
rect 25183 19672 25228 19700
rect 25222 19660 25228 19672
rect 25280 19660 25286 19712
rect 36998 19660 37004 19712
rect 37056 19700 37062 19712
rect 38105 19703 38163 19709
rect 38105 19700 38117 19703
rect 37056 19672 38117 19700
rect 37056 19660 37062 19672
rect 38105 19669 38117 19672
rect 38151 19669 38163 19703
rect 38105 19663 38163 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 7745 19499 7803 19505
rect 7745 19465 7757 19499
rect 7791 19496 7803 19499
rect 12713 19499 12771 19505
rect 7791 19468 10824 19496
rect 7791 19465 7803 19468
rect 7745 19459 7803 19465
rect 8665 19431 8723 19437
rect 8665 19397 8677 19431
rect 8711 19428 8723 19431
rect 8711 19400 10732 19428
rect 8711 19397 8723 19400
rect 8665 19391 8723 19397
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 7653 19363 7711 19369
rect 7653 19360 7665 19363
rect 5684 19332 7665 19360
rect 5684 19320 5690 19332
rect 7653 19329 7665 19332
rect 7699 19329 7711 19363
rect 7653 19323 7711 19329
rect 7742 19320 7748 19372
rect 7800 19360 7806 19372
rect 8573 19363 8631 19369
rect 8573 19360 8585 19363
rect 7800 19332 8585 19360
rect 7800 19320 7806 19332
rect 8573 19329 8585 19332
rect 8619 19329 8631 19363
rect 9214 19360 9220 19372
rect 9175 19332 9220 19360
rect 8573 19323 8631 19329
rect 9214 19320 9220 19332
rect 9272 19320 9278 19372
rect 9309 19363 9367 19369
rect 9309 19329 9321 19363
rect 9355 19360 9367 19363
rect 10594 19360 10600 19372
rect 9355 19332 10600 19360
rect 9355 19329 9367 19332
rect 9309 19323 9367 19329
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19261 9919 19295
rect 10502 19292 10508 19304
rect 10463 19264 10508 19292
rect 9861 19255 9919 19261
rect 9876 19224 9904 19255
rect 10502 19252 10508 19264
rect 10560 19252 10566 19304
rect 10704 19301 10732 19400
rect 10796 19360 10824 19468
rect 12713 19465 12725 19499
rect 12759 19496 12771 19499
rect 12759 19468 13860 19496
rect 12759 19465 12771 19468
rect 12713 19459 12771 19465
rect 11149 19431 11207 19437
rect 11149 19397 11161 19431
rect 11195 19428 11207 19431
rect 11195 19400 12572 19428
rect 11195 19397 11207 19400
rect 11149 19391 11207 19397
rect 12069 19363 12127 19369
rect 12069 19360 12081 19363
rect 10796 19332 12081 19360
rect 12069 19329 12081 19332
rect 12115 19329 12127 19363
rect 12544 19360 12572 19400
rect 12986 19388 12992 19440
rect 13044 19428 13050 19440
rect 13357 19431 13415 19437
rect 13357 19428 13369 19431
rect 13044 19400 13369 19428
rect 13044 19388 13050 19400
rect 13357 19397 13369 19400
rect 13403 19397 13415 19431
rect 13832 19428 13860 19468
rect 13906 19456 13912 19508
rect 13964 19496 13970 19508
rect 14737 19499 14795 19505
rect 14737 19496 14749 19499
rect 13964 19468 14749 19496
rect 13964 19456 13970 19468
rect 14737 19465 14749 19468
rect 14783 19465 14795 19499
rect 14737 19459 14795 19465
rect 14918 19456 14924 19508
rect 14976 19496 14982 19508
rect 16025 19499 16083 19505
rect 16025 19496 16037 19499
rect 14976 19468 16037 19496
rect 14976 19456 14982 19468
rect 16025 19465 16037 19468
rect 16071 19496 16083 19499
rect 16666 19496 16672 19508
rect 16071 19468 16672 19496
rect 16071 19465 16083 19468
rect 16025 19459 16083 19465
rect 16666 19456 16672 19468
rect 16724 19456 16730 19508
rect 16850 19496 16856 19508
rect 16811 19468 16856 19496
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 17494 19496 17500 19508
rect 17455 19468 17500 19496
rect 17494 19456 17500 19468
rect 17552 19456 17558 19508
rect 18138 19496 18144 19508
rect 18099 19468 18144 19496
rect 18138 19456 18144 19468
rect 18196 19456 18202 19508
rect 20898 19496 20904 19508
rect 19904 19468 20904 19496
rect 15286 19428 15292 19440
rect 13832 19400 14136 19428
rect 13357 19391 13415 19397
rect 13078 19360 13084 19372
rect 12544 19332 13084 19360
rect 12069 19323 12127 19329
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 14108 19360 14136 19400
rect 14844 19400 15292 19428
rect 14844 19360 14872 19400
rect 15286 19388 15292 19400
rect 15344 19388 15350 19440
rect 19904 19428 19932 19468
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 22557 19499 22615 19505
rect 22557 19465 22569 19499
rect 22603 19496 22615 19499
rect 22830 19496 22836 19508
rect 22603 19468 22836 19496
rect 22603 19465 22615 19468
rect 22557 19459 22615 19465
rect 22830 19456 22836 19468
rect 22888 19456 22894 19508
rect 24489 19499 24547 19505
rect 24489 19465 24501 19499
rect 24535 19496 24547 19499
rect 25406 19496 25412 19508
rect 24535 19468 25412 19496
rect 24535 19465 24547 19468
rect 24489 19459 24547 19465
rect 25406 19456 25412 19468
rect 25464 19456 25470 19508
rect 20070 19428 20076 19440
rect 15396 19400 19932 19428
rect 20031 19400 20076 19428
rect 14108 19332 14872 19360
rect 14918 19320 14924 19372
rect 14976 19360 14982 19372
rect 14976 19332 15021 19360
rect 14976 19320 14982 19332
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19261 10747 19295
rect 10689 19255 10747 19261
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 11112 19264 12265 19292
rect 11112 19252 11118 19264
rect 12253 19261 12265 19264
rect 12299 19261 12311 19295
rect 12253 19255 12311 19261
rect 13265 19295 13323 19301
rect 13265 19261 13277 19295
rect 13311 19292 13323 19295
rect 13814 19292 13820 19304
rect 13311 19264 13820 19292
rect 13311 19261 13323 19264
rect 13265 19255 13323 19261
rect 13814 19252 13820 19264
rect 13872 19252 13878 19304
rect 13906 19252 13912 19304
rect 13964 19292 13970 19304
rect 15396 19301 15424 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 21358 19388 21364 19440
rect 21416 19428 21422 19440
rect 22002 19428 22008 19440
rect 21416 19400 22008 19428
rect 21416 19388 21422 19400
rect 22002 19388 22008 19400
rect 22060 19428 22066 19440
rect 22060 19400 22508 19428
rect 22060 19388 22066 19400
rect 16758 19320 16764 19372
rect 16816 19360 16822 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16816 19332 17049 19360
rect 16816 19320 16822 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 17126 19320 17132 19372
rect 17184 19360 17190 19372
rect 17681 19363 17739 19369
rect 17681 19360 17693 19363
rect 17184 19332 17693 19360
rect 17184 19320 17190 19332
rect 17681 19329 17693 19332
rect 17727 19329 17739 19363
rect 18782 19360 18788 19372
rect 18743 19332 18788 19360
rect 17681 19323 17739 19329
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 19426 19360 19432 19372
rect 19387 19332 19432 19360
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 21726 19360 21732 19372
rect 21131 19332 21732 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 21726 19320 21732 19332
rect 21784 19320 21790 19372
rect 22480 19369 22508 19400
rect 22922 19388 22928 19440
rect 22980 19428 22986 19440
rect 23385 19431 23443 19437
rect 23385 19428 23397 19431
rect 22980 19400 23397 19428
rect 22980 19388 22986 19400
rect 23385 19397 23397 19400
rect 23431 19397 23443 19431
rect 23385 19391 23443 19397
rect 23477 19431 23535 19437
rect 23477 19397 23489 19431
rect 23523 19428 23535 19431
rect 25222 19428 25228 19440
rect 23523 19400 25228 19428
rect 23523 19397 23535 19400
rect 23477 19391 23535 19397
rect 25222 19388 25228 19400
rect 25280 19388 25286 19440
rect 22465 19363 22523 19369
rect 22465 19329 22477 19363
rect 22511 19329 22523 19363
rect 24670 19360 24676 19372
rect 24631 19332 24676 19360
rect 22465 19323 22523 19329
rect 24670 19320 24676 19332
rect 24728 19320 24734 19372
rect 15381 19295 15439 19301
rect 13964 19264 14009 19292
rect 13964 19252 13970 19264
rect 15381 19261 15393 19295
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19261 15623 19295
rect 18966 19292 18972 19304
rect 18927 19264 18972 19292
rect 15565 19255 15623 19261
rect 11238 19224 11244 19236
rect 9876 19196 11244 19224
rect 11238 19184 11244 19196
rect 11296 19184 11302 19236
rect 11330 19184 11336 19236
rect 11388 19224 11394 19236
rect 11388 19196 12434 19224
rect 11388 19184 11394 19196
rect 7466 19116 7472 19168
rect 7524 19156 7530 19168
rect 12250 19156 12256 19168
rect 7524 19128 12256 19156
rect 7524 19116 7530 19128
rect 12250 19116 12256 19128
rect 12308 19116 12314 19168
rect 12406 19156 12434 19196
rect 12802 19184 12808 19236
rect 12860 19224 12866 19236
rect 15580 19224 15608 19255
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19981 19295 20039 19301
rect 19981 19261 19993 19295
rect 20027 19292 20039 19295
rect 20070 19292 20076 19304
rect 20027 19264 20076 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 23658 19252 23664 19304
rect 23716 19292 23722 19304
rect 24029 19295 24087 19301
rect 24029 19292 24041 19295
rect 23716 19264 24041 19292
rect 23716 19252 23722 19264
rect 24029 19261 24041 19264
rect 24075 19292 24087 19295
rect 29730 19292 29736 19304
rect 24075 19264 29736 19292
rect 24075 19261 24087 19264
rect 24029 19255 24087 19261
rect 29730 19252 29736 19264
rect 29788 19252 29794 19304
rect 12860 19196 15608 19224
rect 12860 19184 12866 19196
rect 20438 19184 20444 19236
rect 20496 19224 20502 19236
rect 20533 19227 20591 19233
rect 20533 19224 20545 19227
rect 20496 19196 20545 19224
rect 20496 19184 20502 19196
rect 20533 19193 20545 19196
rect 20579 19224 20591 19227
rect 28718 19224 28724 19236
rect 20579 19196 28724 19224
rect 20579 19193 20591 19196
rect 20533 19187 20591 19193
rect 28718 19184 28724 19196
rect 28776 19184 28782 19236
rect 13262 19156 13268 19168
rect 12406 19128 13268 19156
rect 13262 19116 13268 19128
rect 13320 19116 13326 19168
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 14366 19156 14372 19168
rect 13412 19128 14372 19156
rect 13412 19116 13418 19128
rect 14366 19116 14372 19128
rect 14424 19156 14430 19168
rect 14918 19156 14924 19168
rect 14424 19128 14924 19156
rect 14424 19116 14430 19128
rect 14918 19116 14924 19128
rect 14976 19116 14982 19168
rect 21174 19156 21180 19168
rect 21135 19128 21180 19156
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 10594 18912 10600 18964
rect 10652 18952 10658 18964
rect 10652 18924 11928 18952
rect 10652 18912 10658 18924
rect 9766 18884 9772 18896
rect 8404 18856 9772 18884
rect 8404 18757 8432 18856
rect 9766 18844 9772 18856
rect 9824 18844 9830 18896
rect 10137 18887 10195 18893
rect 10137 18853 10149 18887
rect 10183 18884 10195 18887
rect 11793 18887 11851 18893
rect 11793 18884 11805 18887
rect 10183 18856 11805 18884
rect 10183 18853 10195 18856
rect 10137 18847 10195 18853
rect 11793 18853 11805 18856
rect 11839 18853 11851 18887
rect 11793 18847 11851 18853
rect 8481 18819 8539 18825
rect 8481 18785 8493 18819
rect 8527 18816 8539 18819
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 8527 18788 9689 18816
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 9677 18785 9689 18788
rect 9723 18785 9735 18819
rect 11609 18819 11667 18825
rect 11609 18816 11621 18819
rect 9677 18779 9735 18785
rect 9784 18788 11621 18816
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 9493 18751 9551 18757
rect 9493 18748 9505 18751
rect 8389 18711 8447 18717
rect 8496 18720 9505 18748
rect 6638 18640 6644 18692
rect 6696 18680 6702 18692
rect 8496 18680 8524 18720
rect 9493 18717 9505 18720
rect 9539 18717 9551 18751
rect 9784 18748 9812 18788
rect 11609 18785 11621 18788
rect 11655 18785 11667 18819
rect 11609 18779 11667 18785
rect 9493 18711 9551 18717
rect 9600 18720 9812 18748
rect 6696 18652 8524 18680
rect 6696 18640 6702 18652
rect 9030 18640 9036 18692
rect 9088 18680 9094 18692
rect 9600 18680 9628 18720
rect 10778 18708 10784 18760
rect 10836 18748 10842 18760
rect 10965 18751 11023 18757
rect 10965 18748 10977 18751
rect 10836 18720 10977 18748
rect 10836 18708 10842 18720
rect 10965 18717 10977 18720
rect 11011 18717 11023 18751
rect 10965 18711 11023 18717
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18717 11483 18751
rect 11425 18711 11483 18717
rect 9088 18652 9628 18680
rect 9088 18640 9094 18652
rect 9674 18640 9680 18692
rect 9732 18680 9738 18692
rect 11440 18680 11468 18711
rect 9732 18652 11468 18680
rect 9732 18640 9738 18652
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7193 18615 7251 18621
rect 7193 18612 7205 18615
rect 7156 18584 7205 18612
rect 7156 18572 7162 18584
rect 7193 18581 7205 18584
rect 7239 18581 7251 18615
rect 7193 18575 7251 18581
rect 10781 18615 10839 18621
rect 10781 18581 10793 18615
rect 10827 18612 10839 18615
rect 11698 18612 11704 18624
rect 10827 18584 11704 18612
rect 10827 18581 10839 18584
rect 10781 18575 10839 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 11808 18612 11836 18847
rect 11900 18680 11928 18924
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 16761 18955 16819 18961
rect 12308 18924 16160 18952
rect 12308 18912 12314 18924
rect 11974 18844 11980 18896
rect 12032 18884 12038 18896
rect 13354 18884 13360 18896
rect 12032 18856 13360 18884
rect 12032 18844 12038 18856
rect 13354 18844 13360 18856
rect 13412 18844 13418 18896
rect 13446 18844 13452 18896
rect 13504 18884 13510 18896
rect 13504 18856 14504 18884
rect 13504 18844 13510 18856
rect 12713 18819 12771 18825
rect 12713 18785 12725 18819
rect 12759 18816 12771 18819
rect 13725 18819 13783 18825
rect 12759 18788 13676 18816
rect 12759 18785 12771 18788
rect 12713 18779 12771 18785
rect 12805 18683 12863 18689
rect 11900 18652 12664 18680
rect 12526 18612 12532 18624
rect 11808 18584 12532 18612
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 12636 18612 12664 18652
rect 12805 18649 12817 18683
rect 12851 18649 12863 18683
rect 13648 18680 13676 18788
rect 13725 18785 13737 18819
rect 13771 18816 13783 18819
rect 13998 18816 14004 18828
rect 13771 18788 14004 18816
rect 13771 18785 13783 18788
rect 13725 18779 13783 18785
rect 13998 18776 14004 18788
rect 14056 18776 14062 18828
rect 14274 18816 14280 18828
rect 14235 18788 14280 18816
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 14476 18825 14504 18856
rect 14461 18819 14519 18825
rect 14461 18785 14473 18819
rect 14507 18785 14519 18819
rect 14461 18779 14519 18785
rect 15654 18748 15660 18760
rect 15615 18720 15660 18748
rect 15654 18708 15660 18720
rect 15712 18708 15718 18760
rect 16132 18757 16160 18924
rect 16761 18921 16773 18955
rect 16807 18952 16819 18955
rect 17126 18952 17132 18964
rect 16807 18924 17132 18952
rect 16807 18921 16819 18924
rect 16761 18915 16819 18921
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 17310 18912 17316 18964
rect 17368 18952 17374 18964
rect 17405 18955 17463 18961
rect 17405 18952 17417 18955
rect 17368 18924 17417 18952
rect 17368 18912 17374 18924
rect 17405 18921 17417 18924
rect 17451 18921 17463 18955
rect 17405 18915 17463 18921
rect 22281 18955 22339 18961
rect 22281 18921 22293 18955
rect 22327 18952 22339 18955
rect 24762 18952 24768 18964
rect 22327 18924 24768 18952
rect 22327 18921 22339 18924
rect 22281 18915 22339 18921
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 18877 18887 18935 18893
rect 18877 18853 18889 18887
rect 18923 18884 18935 18887
rect 20254 18884 20260 18896
rect 18923 18856 20260 18884
rect 18923 18853 18935 18856
rect 18877 18847 18935 18853
rect 20254 18844 20260 18856
rect 20312 18844 20318 18896
rect 20438 18884 20444 18896
rect 20399 18856 20444 18884
rect 20438 18844 20444 18856
rect 20496 18844 20502 18896
rect 30558 18884 30564 18896
rect 21008 18856 30564 18884
rect 16209 18819 16267 18825
rect 16209 18785 16221 18819
rect 16255 18816 16267 18819
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 16255 18788 18429 18816
rect 16255 18785 16267 18788
rect 16209 18779 16267 18785
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 19889 18819 19947 18825
rect 19889 18785 19901 18819
rect 19935 18816 19947 18819
rect 20162 18816 20168 18828
rect 19935 18788 20168 18816
rect 19935 18785 19947 18788
rect 19889 18779 19947 18785
rect 20162 18776 20168 18788
rect 20220 18776 20226 18828
rect 21008 18825 21036 18856
rect 30558 18844 30564 18856
rect 30616 18844 30622 18896
rect 20993 18819 21051 18825
rect 20993 18785 21005 18819
rect 21039 18785 21051 18819
rect 21174 18816 21180 18828
rect 21135 18788 21180 18816
rect 20993 18779 21051 18785
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 23658 18816 23664 18828
rect 23619 18788 23664 18816
rect 23658 18776 23664 18788
rect 23716 18776 23722 18828
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18748 16175 18751
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 16163 18720 16957 18748
rect 16163 18717 16175 18720
rect 16117 18711 16175 18717
rect 16945 18717 16957 18720
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17126 18708 17132 18760
rect 17184 18748 17190 18760
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 17184 18720 17601 18748
rect 17184 18708 17190 18720
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 18230 18748 18236 18760
rect 18191 18720 18236 18748
rect 17589 18711 17647 18717
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 22465 18751 22523 18757
rect 22465 18717 22477 18751
rect 22511 18717 22523 18751
rect 22465 18711 22523 18717
rect 33045 18751 33103 18757
rect 33045 18717 33057 18751
rect 33091 18748 33103 18751
rect 36998 18748 37004 18760
rect 33091 18720 37004 18748
rect 33091 18717 33103 18720
rect 33045 18711 33103 18717
rect 19981 18683 20039 18689
rect 13648 18652 19012 18680
rect 12805 18643 12863 18649
rect 12820 18612 12848 18643
rect 12636 18584 12848 18612
rect 13814 18572 13820 18624
rect 13872 18612 13878 18624
rect 14921 18615 14979 18621
rect 14921 18612 14933 18615
rect 13872 18584 14933 18612
rect 13872 18572 13878 18584
rect 14921 18581 14933 18584
rect 14967 18581 14979 18615
rect 14921 18575 14979 18581
rect 15473 18615 15531 18621
rect 15473 18581 15485 18615
rect 15519 18612 15531 18615
rect 17862 18612 17868 18624
rect 15519 18584 17868 18612
rect 15519 18581 15531 18584
rect 15473 18575 15531 18581
rect 17862 18572 17868 18584
rect 17920 18572 17926 18624
rect 18984 18612 19012 18652
rect 19981 18649 19993 18683
rect 20027 18680 20039 18683
rect 20622 18680 20628 18692
rect 20027 18652 20628 18680
rect 20027 18649 20039 18652
rect 19981 18643 20039 18649
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 21174 18612 21180 18624
rect 18984 18584 21180 18612
rect 21174 18572 21180 18584
rect 21232 18612 21238 18624
rect 21637 18615 21695 18621
rect 21637 18612 21649 18615
rect 21232 18584 21649 18612
rect 21232 18572 21238 18584
rect 21637 18581 21649 18584
rect 21683 18581 21695 18615
rect 22480 18612 22508 18711
rect 36998 18708 37004 18720
rect 37056 18708 37062 18760
rect 38286 18748 38292 18760
rect 38247 18720 38292 18748
rect 38286 18708 38292 18720
rect 38344 18708 38350 18760
rect 23014 18680 23020 18692
rect 22975 18652 23020 18680
rect 23014 18640 23020 18652
rect 23072 18640 23078 18692
rect 23106 18640 23112 18692
rect 23164 18680 23170 18692
rect 23164 18652 23209 18680
rect 23164 18640 23170 18652
rect 23842 18612 23848 18624
rect 22480 18584 23848 18612
rect 21637 18575 21695 18581
rect 23842 18572 23848 18584
rect 23900 18572 23906 18624
rect 33134 18612 33140 18624
rect 33095 18584 33140 18612
rect 33134 18572 33140 18584
rect 33192 18572 33198 18624
rect 34514 18572 34520 18624
rect 34572 18612 34578 18624
rect 38105 18615 38163 18621
rect 38105 18612 38117 18615
rect 34572 18584 38117 18612
rect 34572 18572 34578 18584
rect 38105 18581 38117 18584
rect 38151 18581 38163 18615
rect 38105 18575 38163 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 7650 18368 7656 18420
rect 7708 18368 7714 18420
rect 9030 18408 9036 18420
rect 8991 18380 9036 18408
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9674 18408 9680 18420
rect 9635 18380 9680 18408
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 13354 18408 13360 18420
rect 10520 18380 13360 18408
rect 7098 18340 7104 18352
rect 7059 18312 7104 18340
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 7190 18300 7196 18352
rect 7248 18340 7254 18352
rect 7668 18340 7696 18368
rect 7745 18343 7803 18349
rect 7745 18340 7757 18343
rect 7248 18312 7293 18340
rect 7668 18312 7757 18340
rect 7248 18300 7254 18312
rect 7745 18309 7757 18312
rect 7791 18340 7803 18343
rect 8662 18340 8668 18352
rect 7791 18312 8668 18340
rect 7791 18309 7803 18312
rect 7745 18303 7803 18309
rect 8662 18300 8668 18312
rect 8720 18300 8726 18352
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 8570 18272 8576 18284
rect 8531 18244 8576 18272
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 9214 18272 9220 18284
rect 9175 18244 9220 18272
rect 9214 18232 9220 18244
rect 9272 18232 9278 18284
rect 10520 18281 10548 18380
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 14185 18411 14243 18417
rect 14185 18377 14197 18411
rect 14231 18408 14243 18411
rect 18325 18411 18383 18417
rect 14231 18380 17080 18408
rect 14231 18377 14243 18380
rect 14185 18371 14243 18377
rect 11330 18340 11336 18352
rect 10704 18312 11336 18340
rect 10505 18275 10563 18281
rect 10505 18272 10517 18275
rect 9646 18244 10517 18272
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 9646 18204 9674 18244
rect 10505 18241 10517 18244
rect 10551 18241 10563 18275
rect 10505 18235 10563 18241
rect 7800 18176 9674 18204
rect 7800 18164 7806 18176
rect 10704 18136 10732 18312
rect 11330 18300 11336 18312
rect 11388 18300 11394 18352
rect 17052 18349 17080 18380
rect 18325 18377 18337 18411
rect 18371 18408 18383 18411
rect 18966 18408 18972 18420
rect 18371 18380 18972 18408
rect 18371 18377 18383 18380
rect 18325 18371 18383 18377
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 21174 18408 21180 18420
rect 21135 18380 21180 18408
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 23106 18368 23112 18420
rect 23164 18408 23170 18420
rect 23661 18411 23719 18417
rect 23661 18408 23673 18411
rect 23164 18380 23673 18408
rect 23164 18368 23170 18380
rect 23661 18377 23673 18380
rect 23707 18377 23719 18411
rect 23661 18371 23719 18377
rect 11885 18343 11943 18349
rect 11885 18309 11897 18343
rect 11931 18340 11943 18343
rect 15657 18343 15715 18349
rect 15657 18340 15669 18343
rect 11931 18312 13860 18340
rect 11931 18309 11943 18312
rect 11885 18303 11943 18309
rect 11149 18275 11207 18281
rect 11149 18272 11161 18275
rect 8312 18108 10732 18136
rect 10796 18244 11161 18272
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 3050 18028 3056 18080
rect 3108 18068 3114 18080
rect 3970 18068 3976 18080
rect 3108 18040 3976 18068
rect 3108 18028 3114 18040
rect 3970 18028 3976 18040
rect 4028 18068 4034 18080
rect 8312 18068 8340 18108
rect 4028 18040 8340 18068
rect 8389 18071 8447 18077
rect 4028 18028 4034 18040
rect 8389 18037 8401 18071
rect 8435 18068 8447 18071
rect 8938 18068 8944 18080
rect 8435 18040 8944 18068
rect 8435 18037 8447 18040
rect 8389 18031 8447 18037
rect 8938 18028 8944 18040
rect 8996 18028 9002 18080
rect 10321 18071 10379 18077
rect 10321 18037 10333 18071
rect 10367 18068 10379 18071
rect 10796 18068 10824 18244
rect 11149 18241 11161 18244
rect 11195 18241 11207 18275
rect 11790 18272 11796 18284
rect 11751 18244 11796 18272
rect 11149 18235 11207 18241
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 12621 18275 12679 18281
rect 12621 18241 12633 18275
rect 12667 18272 12679 18275
rect 12986 18272 12992 18284
rect 12667 18244 12992 18272
rect 12667 18241 12679 18244
rect 12621 18235 12679 18241
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 13832 18272 13860 18312
rect 14016 18312 15669 18340
rect 14016 18272 14044 18312
rect 15657 18309 15669 18312
rect 15703 18309 15715 18343
rect 15657 18303 15715 18309
rect 17037 18343 17095 18349
rect 17037 18309 17049 18343
rect 17083 18309 17095 18343
rect 17037 18303 17095 18309
rect 18524 18312 22094 18340
rect 14366 18272 14372 18284
rect 13832 18244 14044 18272
rect 14327 18244 14372 18272
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18272 15071 18275
rect 15059 18244 15148 18272
rect 15059 18241 15071 18244
rect 15013 18235 15071 18241
rect 11238 18164 11244 18216
rect 11296 18204 11302 18216
rect 13081 18207 13139 18213
rect 13081 18204 13093 18207
rect 11296 18176 13093 18204
rect 11296 18164 11302 18176
rect 13081 18173 13093 18176
rect 13127 18173 13139 18207
rect 13081 18167 13139 18173
rect 13265 18207 13323 18213
rect 13265 18173 13277 18207
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 10965 18139 11023 18145
rect 10965 18105 10977 18139
rect 11011 18136 11023 18139
rect 12250 18136 12256 18148
rect 11011 18108 12256 18136
rect 11011 18105 11023 18108
rect 10965 18099 11023 18105
rect 12250 18096 12256 18108
rect 12308 18096 12314 18148
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 12437 18139 12495 18145
rect 12437 18136 12449 18139
rect 12400 18108 12449 18136
rect 12400 18096 12406 18108
rect 12437 18105 12449 18108
rect 12483 18105 12495 18139
rect 12437 18099 12495 18105
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 13280 18136 13308 18167
rect 13354 18164 13360 18216
rect 13412 18204 13418 18216
rect 15120 18204 15148 18244
rect 17586 18232 17592 18284
rect 17644 18272 17650 18284
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 17644 18244 18245 18272
rect 17644 18232 17650 18244
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 13412 18176 15148 18204
rect 13412 18164 13418 18176
rect 12584 18108 13308 18136
rect 12584 18096 12590 18108
rect 10367 18040 10824 18068
rect 10367 18037 10379 18040
rect 10321 18031 10379 18037
rect 13078 18028 13084 18080
rect 13136 18068 13142 18080
rect 13725 18071 13783 18077
rect 13725 18068 13737 18071
rect 13136 18040 13737 18068
rect 13136 18028 13142 18040
rect 13725 18037 13737 18040
rect 13771 18068 13783 18071
rect 14090 18068 14096 18080
rect 13771 18040 14096 18068
rect 13771 18037 13783 18040
rect 13725 18031 13783 18037
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 14826 18068 14832 18080
rect 14787 18040 14832 18068
rect 14826 18028 14832 18040
rect 14884 18028 14890 18080
rect 15120 18068 15148 18176
rect 15286 18164 15292 18216
rect 15344 18204 15350 18216
rect 15565 18207 15623 18213
rect 15565 18204 15577 18207
rect 15344 18176 15577 18204
rect 15344 18164 15350 18176
rect 15565 18173 15577 18176
rect 15611 18173 15623 18207
rect 16942 18204 16948 18216
rect 16903 18176 16948 18204
rect 15565 18167 15623 18173
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17405 18207 17463 18213
rect 17405 18173 17417 18207
rect 17451 18204 17463 18207
rect 18524 18204 18552 18312
rect 18877 18275 18935 18281
rect 18877 18241 18889 18275
rect 18923 18272 18935 18275
rect 21542 18272 21548 18284
rect 18923 18244 21548 18272
rect 18923 18241 18935 18244
rect 18877 18235 18935 18241
rect 21542 18232 21548 18244
rect 21600 18232 21606 18284
rect 19058 18204 19064 18216
rect 17451 18176 18552 18204
rect 19019 18176 19064 18204
rect 17451 18173 17463 18176
rect 17405 18167 17463 18173
rect 16117 18139 16175 18145
rect 16117 18105 16129 18139
rect 16163 18136 16175 18139
rect 17420 18136 17448 18167
rect 19058 18164 19064 18176
rect 19116 18164 19122 18216
rect 20533 18207 20591 18213
rect 20533 18173 20545 18207
rect 20579 18173 20591 18207
rect 20714 18204 20720 18216
rect 20675 18176 20720 18204
rect 20533 18167 20591 18173
rect 16163 18108 17448 18136
rect 16163 18105 16175 18108
rect 16117 18099 16175 18105
rect 18138 18068 18144 18080
rect 15120 18040 18144 18068
rect 18138 18028 18144 18040
rect 18196 18028 18202 18080
rect 19521 18071 19579 18077
rect 19521 18037 19533 18071
rect 19567 18068 19579 18071
rect 20346 18068 20352 18080
rect 19567 18040 20352 18068
rect 19567 18037 19579 18040
rect 19521 18031 19579 18037
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 20548 18068 20576 18167
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 22066 18136 22094 18312
rect 22465 18275 22523 18281
rect 22465 18241 22477 18275
rect 22511 18272 22523 18275
rect 22511 18244 23520 18272
rect 22511 18241 22523 18244
rect 22465 18235 22523 18241
rect 22646 18204 22652 18216
rect 22607 18176 22652 18204
rect 22646 18164 22652 18176
rect 22704 18164 22710 18216
rect 23492 18204 23520 18244
rect 23566 18232 23572 18284
rect 23624 18272 23630 18284
rect 24394 18272 24400 18284
rect 23624 18244 23669 18272
rect 24355 18244 24400 18272
rect 23624 18232 23630 18244
rect 24394 18232 24400 18244
rect 24452 18232 24458 18284
rect 33318 18204 33324 18216
rect 23492 18176 33324 18204
rect 33318 18164 33324 18176
rect 33376 18164 33382 18216
rect 29638 18136 29644 18148
rect 22066 18108 29644 18136
rect 29638 18096 29644 18108
rect 29696 18096 29702 18148
rect 21634 18068 21640 18080
rect 20548 18040 21640 18068
rect 21634 18028 21640 18040
rect 21692 18028 21698 18080
rect 22738 18028 22744 18080
rect 22796 18068 22802 18080
rect 22833 18071 22891 18077
rect 22833 18068 22845 18071
rect 22796 18040 22845 18068
rect 22796 18028 22802 18040
rect 22833 18037 22845 18040
rect 22879 18037 22891 18071
rect 24210 18068 24216 18080
rect 24171 18040 24216 18068
rect 22833 18031 22891 18037
rect 24210 18028 24216 18040
rect 24268 18028 24274 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 7101 17867 7159 17873
rect 7101 17833 7113 17867
rect 7147 17864 7159 17867
rect 7190 17864 7196 17876
rect 7147 17836 7196 17864
rect 7147 17833 7159 17836
rect 7101 17827 7159 17833
rect 7190 17824 7196 17836
rect 7248 17824 7254 17876
rect 9214 17824 9220 17876
rect 9272 17864 9278 17876
rect 9493 17867 9551 17873
rect 9493 17864 9505 17867
rect 9272 17836 9505 17864
rect 9272 17824 9278 17836
rect 9493 17833 9505 17836
rect 9539 17833 9551 17867
rect 9493 17827 9551 17833
rect 13725 17867 13783 17873
rect 13725 17833 13737 17867
rect 13771 17864 13783 17867
rect 13814 17864 13820 17876
rect 13771 17836 13820 17864
rect 13771 17833 13783 17836
rect 13725 17827 13783 17833
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 16942 17864 16948 17876
rect 16903 17836 16948 17864
rect 16942 17824 16948 17836
rect 17000 17824 17006 17876
rect 18230 17864 18236 17876
rect 17604 17836 18236 17864
rect 10134 17756 10140 17808
rect 10192 17756 10198 17808
rect 11885 17799 11943 17805
rect 11885 17765 11897 17799
rect 11931 17796 11943 17799
rect 14458 17796 14464 17808
rect 11931 17768 14464 17796
rect 11931 17765 11943 17768
rect 11885 17759 11943 17765
rect 14458 17756 14464 17768
rect 14516 17756 14522 17808
rect 14645 17799 14703 17805
rect 14645 17765 14657 17799
rect 14691 17796 14703 17799
rect 16114 17796 16120 17808
rect 14691 17768 16120 17796
rect 14691 17765 14703 17768
rect 14645 17759 14703 17765
rect 16114 17756 16120 17768
rect 16172 17756 16178 17808
rect 16298 17756 16304 17808
rect 16356 17796 16362 17808
rect 16356 17768 17172 17796
rect 16356 17756 16362 17768
rect 7834 17728 7840 17740
rect 7747 17700 7840 17728
rect 1949 17663 2007 17669
rect 1949 17629 1961 17663
rect 1995 17660 2007 17663
rect 2314 17660 2320 17672
rect 1995 17632 2320 17660
rect 1995 17629 2007 17632
rect 1949 17623 2007 17629
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17660 2467 17663
rect 2774 17660 2780 17672
rect 2455 17632 2780 17660
rect 2455 17629 2467 17632
rect 2409 17623 2467 17629
rect 2774 17620 2780 17632
rect 2832 17620 2838 17672
rect 3234 17660 3240 17672
rect 3195 17632 3240 17660
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 5166 17660 5172 17672
rect 5127 17632 5172 17660
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17660 6699 17663
rect 7006 17660 7012 17672
rect 6687 17632 7012 17660
rect 6687 17629 6699 17632
rect 6641 17623 6699 17629
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 7760 17669 7788 17700
rect 7834 17688 7840 17700
rect 7892 17728 7898 17740
rect 8846 17728 8852 17740
rect 7892 17700 8852 17728
rect 7892 17688 7898 17700
rect 8846 17688 8852 17700
rect 8904 17688 8910 17740
rect 9766 17728 9772 17740
rect 9679 17700 9772 17728
rect 9692 17669 9720 17700
rect 9766 17688 9772 17700
rect 9824 17728 9830 17740
rect 10152 17728 10180 17756
rect 10870 17728 10876 17740
rect 9824 17700 10180 17728
rect 10831 17700 10876 17728
rect 9824 17688 9830 17700
rect 10870 17688 10876 17700
rect 10928 17688 10934 17740
rect 12986 17728 12992 17740
rect 11808 17700 12992 17728
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 7745 17663 7803 17669
rect 7745 17629 7757 17663
rect 7791 17629 7803 17663
rect 7745 17623 7803 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 7300 17592 7328 17623
rect 6472 17564 7328 17592
rect 8588 17592 8616 17623
rect 10962 17620 10968 17672
rect 11020 17660 11026 17672
rect 11808 17669 11836 17700
rect 12986 17688 12992 17700
rect 13044 17688 13050 17740
rect 13081 17731 13139 17737
rect 13081 17697 13093 17731
rect 13127 17728 13139 17731
rect 13538 17728 13544 17740
rect 13127 17700 13544 17728
rect 13127 17697 13139 17700
rect 13081 17691 13139 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 15378 17728 15384 17740
rect 15339 17700 15384 17728
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 16022 17728 16028 17740
rect 15983 17700 16028 17728
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11020 17632 11805 17660
rect 11020 17620 11026 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 12342 17620 12348 17672
rect 12400 17660 12406 17672
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 12400 17632 12633 17660
rect 12400 17620 12406 17632
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 12710 17620 12716 17672
rect 12768 17660 12774 17672
rect 13265 17663 13323 17669
rect 13265 17660 13277 17663
rect 12768 17632 13277 17660
rect 12768 17620 12774 17632
rect 13265 17629 13277 17632
rect 13311 17629 13323 17663
rect 14826 17660 14832 17672
rect 14787 17632 14832 17660
rect 13265 17623 13323 17629
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 16482 17660 16488 17672
rect 16443 17632 16488 17660
rect 16482 17620 16488 17632
rect 16540 17620 16546 17672
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17629 16727 17663
rect 17144 17660 17172 17768
rect 17604 17737 17632 17836
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 18693 17867 18751 17873
rect 18693 17833 18705 17867
rect 18739 17864 18751 17867
rect 19058 17864 19064 17876
rect 18739 17836 19064 17864
rect 18739 17833 18751 17836
rect 18693 17827 18751 17833
rect 19058 17824 19064 17836
rect 19116 17824 19122 17876
rect 19812 17836 20668 17864
rect 19812 17737 19840 17836
rect 17589 17731 17647 17737
rect 17589 17697 17601 17731
rect 17635 17697 17647 17731
rect 17589 17691 17647 17697
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 20441 17731 20499 17737
rect 20441 17697 20453 17731
rect 20487 17697 20499 17731
rect 20640 17728 20668 17836
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 20901 17867 20959 17873
rect 20901 17864 20913 17867
rect 20772 17836 20913 17864
rect 20772 17824 20778 17836
rect 20901 17833 20913 17836
rect 20947 17833 20959 17867
rect 20901 17827 20959 17833
rect 21545 17867 21603 17873
rect 21545 17833 21557 17867
rect 21591 17833 21603 17867
rect 21545 17827 21603 17833
rect 21174 17728 21180 17740
rect 20640 17700 21180 17728
rect 20441 17691 20499 17697
rect 17773 17663 17831 17669
rect 17773 17660 17785 17663
rect 17144 17632 17785 17660
rect 16669 17623 16727 17629
rect 17773 17629 17785 17632
rect 17819 17629 17831 17663
rect 17773 17623 17831 17629
rect 9766 17592 9772 17604
rect 8588 17564 9772 17592
rect 1765 17527 1823 17533
rect 1765 17493 1777 17527
rect 1811 17524 1823 17527
rect 1854 17524 1860 17536
rect 1811 17496 1860 17524
rect 1811 17493 1823 17496
rect 1765 17487 1823 17493
rect 1854 17484 1860 17496
rect 1912 17484 1918 17536
rect 2498 17524 2504 17536
rect 2459 17496 2504 17524
rect 2498 17484 2504 17496
rect 2556 17484 2562 17536
rect 2590 17484 2596 17536
rect 2648 17524 2654 17536
rect 3053 17527 3111 17533
rect 3053 17524 3065 17527
rect 2648 17496 3065 17524
rect 2648 17484 2654 17496
rect 3053 17493 3065 17496
rect 3099 17493 3111 17527
rect 3053 17487 3111 17493
rect 4706 17484 4712 17536
rect 4764 17524 4770 17536
rect 6472 17533 6500 17564
rect 9766 17552 9772 17564
rect 9824 17552 9830 17604
rect 10226 17592 10232 17604
rect 10187 17564 10232 17592
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 10321 17595 10379 17601
rect 10321 17561 10333 17595
rect 10367 17561 10379 17595
rect 10321 17555 10379 17561
rect 12452 17564 15332 17592
rect 4985 17527 5043 17533
rect 4985 17524 4997 17527
rect 4764 17496 4997 17524
rect 4764 17484 4770 17496
rect 4985 17493 4997 17496
rect 5031 17493 5043 17527
rect 4985 17487 5043 17493
rect 6457 17527 6515 17533
rect 6457 17493 6469 17527
rect 6503 17493 6515 17527
rect 6457 17487 6515 17493
rect 7837 17527 7895 17533
rect 7837 17493 7849 17527
rect 7883 17524 7895 17527
rect 8294 17524 8300 17536
rect 7883 17496 8300 17524
rect 7883 17493 7895 17496
rect 7837 17487 7895 17493
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 8389 17527 8447 17533
rect 8389 17493 8401 17527
rect 8435 17524 8447 17527
rect 10336 17524 10364 17555
rect 12452 17533 12480 17564
rect 8435 17496 10364 17524
rect 12437 17527 12495 17533
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 12437 17493 12449 17527
rect 12483 17493 12495 17527
rect 15304 17524 15332 17564
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 15528 17564 15573 17592
rect 15528 17552 15534 17564
rect 16684 17524 16712 17623
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 18877 17663 18935 17669
rect 18877 17660 18889 17663
rect 17920 17632 18889 17660
rect 17920 17620 17926 17632
rect 18877 17629 18889 17632
rect 18923 17629 18935 17663
rect 18877 17623 18935 17629
rect 16850 17552 16856 17604
rect 16908 17592 16914 17604
rect 19889 17595 19947 17601
rect 19889 17592 19901 17595
rect 16908 17564 19901 17592
rect 16908 17552 16914 17564
rect 19889 17561 19901 17564
rect 19935 17561 19947 17595
rect 19889 17555 19947 17561
rect 20456 17592 20484 17691
rect 21174 17688 21180 17700
rect 21232 17688 21238 17740
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17660 21143 17663
rect 21560 17660 21588 17827
rect 21634 17824 21640 17876
rect 21692 17864 21698 17876
rect 21692 17836 22232 17864
rect 21692 17824 21698 17836
rect 22204 17737 22232 17836
rect 22646 17824 22652 17876
rect 22704 17864 22710 17876
rect 23385 17867 23443 17873
rect 23385 17864 23397 17867
rect 22704 17836 23397 17864
rect 22704 17824 22710 17836
rect 23385 17833 23397 17836
rect 23431 17833 23443 17867
rect 23385 17827 23443 17833
rect 22738 17796 22744 17808
rect 22699 17768 22744 17796
rect 22738 17756 22744 17768
rect 22796 17756 22802 17808
rect 22189 17731 22247 17737
rect 22189 17697 22201 17731
rect 22235 17728 22247 17731
rect 22278 17728 22284 17740
rect 22235 17700 22284 17728
rect 22235 17697 22247 17700
rect 22189 17691 22247 17697
rect 22278 17688 22284 17700
rect 22336 17688 22342 17740
rect 22373 17731 22431 17737
rect 22373 17697 22385 17731
rect 22419 17728 22431 17731
rect 24210 17728 24216 17740
rect 22419 17700 24216 17728
rect 22419 17697 22431 17700
rect 22373 17691 22431 17697
rect 24210 17688 24216 17700
rect 24268 17688 24274 17740
rect 38102 17728 38108 17740
rect 31496 17700 38108 17728
rect 21726 17660 21732 17672
rect 21131 17632 21588 17660
rect 21687 17632 21732 17660
rect 21131 17629 21143 17632
rect 21085 17623 21143 17629
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 23290 17660 23296 17672
rect 23251 17632 23296 17660
rect 23290 17620 23296 17632
rect 23348 17620 23354 17672
rect 31496 17669 31524 17700
rect 38102 17688 38108 17700
rect 38160 17688 38166 17740
rect 31481 17663 31539 17669
rect 31481 17629 31493 17663
rect 31527 17629 31539 17663
rect 31481 17623 31539 17629
rect 33137 17663 33195 17669
rect 33137 17629 33149 17663
rect 33183 17660 33195 17663
rect 34514 17660 34520 17672
rect 33183 17632 34520 17660
rect 33183 17629 33195 17632
rect 33137 17623 33195 17629
rect 34514 17620 34520 17632
rect 34572 17620 34578 17672
rect 29086 17592 29092 17604
rect 20456 17564 29092 17592
rect 20456 17536 20484 17564
rect 29086 17552 29092 17564
rect 29144 17552 29150 17604
rect 18230 17524 18236 17536
rect 15304 17496 16712 17524
rect 18191 17496 18236 17524
rect 12437 17487 12495 17493
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 20438 17484 20444 17536
rect 20496 17484 20502 17536
rect 31570 17524 31576 17536
rect 31531 17496 31576 17524
rect 31570 17484 31576 17496
rect 31628 17484 31634 17536
rect 33226 17524 33232 17536
rect 33187 17496 33232 17524
rect 33226 17484 33232 17496
rect 33284 17484 33290 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 8570 17320 8576 17332
rect 8531 17292 8576 17320
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10321 17323 10379 17329
rect 10321 17320 10333 17323
rect 10284 17292 10333 17320
rect 10284 17280 10290 17292
rect 10321 17289 10333 17292
rect 10367 17289 10379 17323
rect 11054 17320 11060 17332
rect 11015 17292 11060 17320
rect 10321 17283 10379 17289
rect 11054 17280 11060 17292
rect 11112 17280 11118 17332
rect 12897 17323 12955 17329
rect 12897 17289 12909 17323
rect 12943 17289 12955 17323
rect 12897 17283 12955 17289
rect 13541 17323 13599 17329
rect 13541 17289 13553 17323
rect 13587 17320 13599 17323
rect 16482 17320 16488 17332
rect 13587 17292 16488 17320
rect 13587 17289 13599 17292
rect 13541 17283 13599 17289
rect 4706 17252 4712 17264
rect 4667 17224 4712 17252
rect 4706 17212 4712 17224
rect 4764 17212 4770 17264
rect 11790 17212 11796 17264
rect 11848 17252 11854 17264
rect 12912 17252 12940 17283
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 16942 17280 16948 17332
rect 17000 17320 17006 17332
rect 17497 17323 17555 17329
rect 17497 17320 17509 17323
rect 17000 17292 17509 17320
rect 17000 17280 17006 17292
rect 17497 17289 17509 17292
rect 17543 17289 17555 17323
rect 17497 17283 17555 17289
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 19978 17320 19984 17332
rect 19484 17292 19984 17320
rect 19484 17280 19490 17292
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 20993 17323 21051 17329
rect 20993 17320 21005 17323
rect 20864 17292 21005 17320
rect 20864 17280 20870 17292
rect 20993 17289 21005 17292
rect 21039 17289 21051 17323
rect 20993 17283 21051 17289
rect 22649 17323 22707 17329
rect 22649 17289 22661 17323
rect 22695 17320 22707 17323
rect 23014 17320 23020 17332
rect 22695 17292 23020 17320
rect 22695 17289 22707 17292
rect 22649 17283 22707 17289
rect 23014 17280 23020 17292
rect 23072 17280 23078 17332
rect 23109 17323 23167 17329
rect 23109 17289 23121 17323
rect 23155 17320 23167 17323
rect 24394 17320 24400 17332
rect 23155 17292 24400 17320
rect 23155 17289 23167 17292
rect 23109 17283 23167 17289
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 14366 17252 14372 17264
rect 11848 17224 12664 17252
rect 12912 17224 14372 17252
rect 11848 17212 11854 17224
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 2406 17184 2412 17196
rect 1903 17156 2412 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 2593 17187 2651 17193
rect 2593 17153 2605 17187
rect 2639 17184 2651 17187
rect 2774 17184 2780 17196
rect 2639 17156 2780 17184
rect 2639 17153 2651 17156
rect 2593 17147 2651 17153
rect 2774 17144 2780 17156
rect 2832 17184 2838 17196
rect 3142 17184 3148 17196
rect 2832 17156 3148 17184
rect 2832 17144 2838 17156
rect 3142 17144 3148 17156
rect 3200 17184 3206 17196
rect 3237 17187 3295 17193
rect 3237 17184 3249 17187
rect 3200 17156 3249 17184
rect 3200 17144 3206 17156
rect 3237 17153 3249 17156
rect 3283 17153 3295 17187
rect 3237 17147 3295 17153
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 7282 17184 7288 17196
rect 5859 17156 7288 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 8846 17184 8852 17196
rect 8803 17156 8852 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 8846 17144 8852 17156
rect 8904 17144 8910 17196
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9401 17187 9459 17193
rect 9401 17184 9413 17187
rect 8996 17156 9413 17184
rect 8996 17144 9002 17156
rect 9401 17153 9413 17156
rect 9447 17153 9459 17187
rect 10962 17184 10968 17196
rect 10923 17156 10968 17184
rect 9401 17147 9459 17153
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12636 17184 12664 17224
rect 14366 17212 14372 17224
rect 14424 17212 14430 17264
rect 14829 17255 14887 17261
rect 14829 17221 14841 17255
rect 14875 17252 14887 17255
rect 15286 17252 15292 17264
rect 14875 17224 15292 17252
rect 14875 17221 14887 17224
rect 14829 17215 14887 17221
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 15473 17255 15531 17261
rect 15473 17221 15485 17255
rect 15519 17252 15531 17255
rect 18877 17255 18935 17261
rect 15519 17224 18276 17252
rect 15519 17221 15531 17224
rect 15473 17215 15531 17221
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12492 17156 12537 17184
rect 12636 17156 13093 17184
rect 12492 17144 12498 17156
rect 13081 17153 13093 17156
rect 13127 17184 13139 17187
rect 13262 17184 13268 17196
rect 13127 17156 13268 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 16758 17184 16764 17196
rect 16347 17156 16764 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 17218 17184 17224 17196
rect 16899 17156 17224 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 17218 17144 17224 17156
rect 17276 17144 17282 17196
rect 18248 17193 18276 17224
rect 18877 17221 18889 17255
rect 18923 17252 18935 17255
rect 20070 17252 20076 17264
rect 18923 17224 20076 17252
rect 18923 17221 18935 17224
rect 18877 17215 18935 17221
rect 20070 17212 20076 17224
rect 20128 17252 20134 17264
rect 20254 17252 20260 17264
rect 20128 17224 20260 17252
rect 20128 17212 20134 17224
rect 20254 17212 20260 17224
rect 20312 17212 20318 17264
rect 31570 17252 31576 17264
rect 20364 17224 31576 17252
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 18966 17144 18972 17196
rect 19024 17184 19030 17196
rect 20364 17184 20392 17224
rect 31570 17212 31576 17224
rect 31628 17212 31634 17264
rect 19024 17156 20392 17184
rect 21177 17187 21235 17193
rect 19024 17144 19030 17156
rect 21177 17153 21189 17187
rect 21223 17184 21235 17187
rect 23106 17184 23112 17196
rect 21223 17156 23112 17184
rect 21223 17153 21235 17156
rect 21177 17147 21235 17153
rect 23106 17144 23112 17156
rect 23164 17144 23170 17196
rect 23290 17184 23296 17196
rect 23251 17156 23296 17184
rect 23290 17144 23296 17156
rect 23348 17144 23354 17196
rect 23842 17144 23848 17196
rect 23900 17184 23906 17196
rect 23937 17187 23995 17193
rect 23937 17184 23949 17187
rect 23900 17156 23949 17184
rect 23900 17144 23906 17156
rect 23937 17153 23949 17156
rect 23983 17153 23995 17187
rect 24578 17184 24584 17196
rect 24539 17156 24584 17184
rect 23937 17147 23995 17153
rect 24578 17144 24584 17156
rect 24636 17144 24642 17196
rect 35894 17144 35900 17196
rect 35952 17184 35958 17196
rect 38013 17187 38071 17193
rect 38013 17184 38025 17187
rect 35952 17156 38025 17184
rect 35952 17144 35958 17156
rect 38013 17153 38025 17156
rect 38059 17153 38071 17187
rect 38013 17147 38071 17153
rect 4614 17116 4620 17128
rect 4575 17088 4620 17116
rect 4614 17076 4620 17088
rect 4672 17076 4678 17128
rect 4798 17076 4804 17128
rect 4856 17116 4862 17128
rect 4893 17119 4951 17125
rect 4893 17116 4905 17119
rect 4856 17088 4905 17116
rect 4856 17076 4862 17088
rect 4893 17085 4905 17088
rect 4939 17085 4951 17119
rect 4893 17079 4951 17085
rect 6733 17119 6791 17125
rect 6733 17085 6745 17119
rect 6779 17116 6791 17119
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 6779 17088 7389 17116
rect 6779 17085 6791 17088
rect 6733 17079 6791 17085
rect 7377 17085 7389 17088
rect 7423 17085 7435 17119
rect 7558 17116 7564 17128
rect 7519 17088 7564 17116
rect 7377 17079 7435 17085
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 9217 17119 9275 17125
rect 9217 17085 9229 17119
rect 9263 17116 9275 17119
rect 9306 17116 9312 17128
rect 9263 17088 9312 17116
rect 9263 17085 9275 17088
rect 9217 17079 9275 17085
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 14185 17119 14243 17125
rect 14185 17085 14197 17119
rect 14231 17116 14243 17119
rect 14274 17116 14280 17128
rect 14231 17088 14280 17116
rect 14231 17085 14243 17088
rect 14185 17079 14243 17085
rect 14274 17076 14280 17088
rect 14332 17076 14338 17128
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17085 14427 17119
rect 14369 17079 14427 17085
rect 3326 17048 3332 17060
rect 3287 17020 3332 17048
rect 3326 17008 3332 17020
rect 3384 17008 3390 17060
rect 9324 17048 9352 17076
rect 11422 17048 11428 17060
rect 9324 17020 11428 17048
rect 11422 17008 11428 17020
rect 11480 17008 11486 17060
rect 11606 17008 11612 17060
rect 11664 17048 11670 17060
rect 14384 17048 14412 17079
rect 14458 17076 14464 17128
rect 14516 17116 14522 17128
rect 17037 17119 17095 17125
rect 14516 17088 16068 17116
rect 14516 17076 14522 17088
rect 15470 17048 15476 17060
rect 11664 17020 14412 17048
rect 14476 17020 15476 17048
rect 11664 17008 11670 17020
rect 1949 16983 2007 16989
rect 1949 16949 1961 16983
rect 1995 16980 2007 16983
rect 2130 16980 2136 16992
rect 1995 16952 2136 16980
rect 1995 16949 2007 16952
rect 1949 16943 2007 16949
rect 2130 16940 2136 16952
rect 2188 16940 2194 16992
rect 2682 16980 2688 16992
rect 2643 16952 2688 16980
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 5905 16983 5963 16989
rect 5905 16949 5917 16983
rect 5951 16980 5963 16983
rect 6454 16980 6460 16992
rect 5951 16952 6460 16980
rect 5951 16949 5963 16952
rect 5905 16943 5963 16949
rect 6454 16940 6460 16952
rect 6512 16940 6518 16992
rect 6914 16940 6920 16992
rect 6972 16980 6978 16992
rect 7745 16983 7803 16989
rect 7745 16980 7757 16983
rect 6972 16952 7757 16980
rect 6972 16940 6978 16952
rect 7745 16949 7757 16952
rect 7791 16949 7803 16983
rect 9674 16980 9680 16992
rect 9635 16952 9680 16980
rect 7745 16943 7803 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 12253 16983 12311 16989
rect 12253 16949 12265 16983
rect 12299 16980 12311 16983
rect 14476 16980 14504 17020
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 16040 17048 16068 17088
rect 17037 17085 17049 17119
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17085 18475 17119
rect 19334 17116 19340 17128
rect 19295 17088 19340 17116
rect 18417 17079 18475 17085
rect 17052 17048 17080 17079
rect 16040 17020 17080 17048
rect 18432 17048 18460 17079
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 19521 17119 19579 17125
rect 19521 17116 19533 17119
rect 19484 17088 19533 17116
rect 19484 17076 19490 17088
rect 19521 17085 19533 17088
rect 19567 17085 19579 17119
rect 22002 17116 22008 17128
rect 21963 17088 22008 17116
rect 19521 17079 19579 17085
rect 22002 17076 22008 17088
rect 22060 17076 22066 17128
rect 22189 17119 22247 17125
rect 22189 17085 22201 17119
rect 22235 17116 22247 17119
rect 22830 17116 22836 17128
rect 22235 17088 22836 17116
rect 22235 17085 22247 17088
rect 22189 17079 22247 17085
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 24397 17051 24455 17057
rect 24397 17048 24409 17051
rect 18432 17020 24409 17048
rect 24397 17017 24409 17020
rect 24443 17017 24455 17051
rect 38194 17048 38200 17060
rect 38155 17020 38200 17048
rect 24397 17011 24455 17017
rect 38194 17008 38200 17020
rect 38252 17008 38258 17060
rect 12299 16952 14504 16980
rect 16117 16983 16175 16989
rect 12299 16949 12311 16952
rect 12253 16943 12311 16949
rect 16117 16949 16129 16983
rect 16163 16980 16175 16983
rect 16850 16980 16856 16992
rect 16163 16952 16856 16980
rect 16163 16949 16175 16952
rect 16117 16943 16175 16949
rect 16850 16940 16856 16952
rect 16908 16940 16914 16992
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 22002 16980 22008 16992
rect 17368 16952 22008 16980
rect 17368 16940 17374 16952
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 23474 16940 23480 16992
rect 23532 16980 23538 16992
rect 23753 16983 23811 16989
rect 23753 16980 23765 16983
rect 23532 16952 23765 16980
rect 23532 16940 23538 16952
rect 23753 16949 23765 16952
rect 23799 16949 23811 16983
rect 23753 16943 23811 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 11606 16776 11612 16788
rect 11567 16748 11612 16776
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 12897 16779 12955 16785
rect 12897 16776 12909 16779
rect 12492 16748 12909 16776
rect 12492 16736 12498 16748
rect 12897 16745 12909 16748
rect 12943 16745 12955 16779
rect 16758 16776 16764 16788
rect 16719 16748 16764 16776
rect 12897 16739 12955 16745
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 22830 16736 22836 16788
rect 22888 16776 22894 16788
rect 22888 16748 22933 16776
rect 22888 16736 22894 16748
rect 8478 16708 8484 16720
rect 8439 16680 8484 16708
rect 8478 16668 8484 16680
rect 8536 16668 8542 16720
rect 10965 16711 11023 16717
rect 10965 16677 10977 16711
rect 11011 16708 11023 16711
rect 13354 16708 13360 16720
rect 11011 16680 13360 16708
rect 11011 16677 11023 16680
rect 10965 16671 11023 16677
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 16022 16708 16028 16720
rect 15983 16680 16028 16708
rect 16022 16668 16028 16680
rect 16080 16668 16086 16720
rect 20073 16711 20131 16717
rect 20073 16677 20085 16711
rect 20119 16708 20131 16711
rect 20438 16708 20444 16720
rect 20119 16680 20444 16708
rect 20119 16677 20131 16680
rect 20073 16671 20131 16677
rect 20438 16668 20444 16680
rect 20496 16668 20502 16720
rect 20898 16708 20904 16720
rect 20640 16680 20904 16708
rect 2424 16612 4016 16640
rect 2424 16584 2452 16612
rect 1581 16575 1639 16581
rect 1581 16541 1593 16575
rect 1627 16572 1639 16575
rect 1670 16572 1676 16584
rect 1627 16544 1676 16572
rect 1627 16541 1639 16544
rect 1581 16535 1639 16541
rect 1670 16532 1676 16544
rect 1728 16532 1734 16584
rect 2317 16575 2375 16581
rect 2317 16541 2329 16575
rect 2363 16572 2375 16575
rect 2406 16572 2412 16584
rect 2363 16544 2412 16572
rect 2363 16541 2375 16544
rect 2317 16535 2375 16541
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 2958 16572 2964 16584
rect 2919 16544 2964 16572
rect 2958 16532 2964 16544
rect 3016 16532 3022 16584
rect 3988 16581 4016 16612
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 4709 16643 4767 16649
rect 4709 16640 4721 16643
rect 4672 16612 4721 16640
rect 4672 16600 4678 16612
rect 4709 16609 4721 16612
rect 4755 16609 4767 16643
rect 4709 16603 4767 16609
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 6270 16640 6276 16652
rect 5592 16612 5672 16640
rect 6231 16612 6276 16640
rect 5592 16600 5598 16612
rect 5644 16581 5672 16612
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 6454 16640 6460 16652
rect 6415 16612 6460 16640
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 7926 16640 7932 16652
rect 7887 16612 7932 16640
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 9309 16643 9367 16649
rect 9309 16640 9321 16643
rect 8352 16612 9321 16640
rect 8352 16600 8358 16612
rect 9309 16609 9321 16612
rect 9355 16609 9367 16643
rect 12710 16640 12716 16652
rect 9309 16603 9367 16609
rect 9416 16612 12716 16640
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16541 4031 16575
rect 3973 16535 4031 16541
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16541 5687 16575
rect 5629 16535 5687 16541
rect 9030 16532 9036 16584
rect 9088 16572 9094 16584
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 9088 16544 9137 16572
rect 9088 16532 9094 16544
rect 9125 16541 9137 16544
rect 9171 16572 9183 16575
rect 9416 16572 9444 16612
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16640 15531 16643
rect 17402 16640 17408 16652
rect 15519 16612 17408 16640
rect 15519 16609 15531 16612
rect 15473 16603 15531 16609
rect 17402 16600 17408 16612
rect 17460 16600 17466 16652
rect 18506 16600 18512 16652
rect 18564 16640 18570 16652
rect 20640 16649 20668 16680
rect 20898 16668 20904 16680
rect 20956 16668 20962 16720
rect 23477 16711 23535 16717
rect 23477 16708 23489 16711
rect 21928 16680 23489 16708
rect 19521 16643 19579 16649
rect 19521 16640 19533 16643
rect 18564 16612 19533 16640
rect 18564 16600 18570 16612
rect 19521 16609 19533 16612
rect 19567 16609 19579 16643
rect 19521 16603 19579 16609
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16609 20683 16643
rect 20625 16603 20683 16609
rect 20809 16643 20867 16649
rect 20809 16609 20821 16643
rect 20855 16640 20867 16643
rect 21266 16640 21272 16652
rect 20855 16612 21272 16640
rect 20855 16609 20867 16612
rect 20809 16603 20867 16609
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 21729 16643 21787 16649
rect 21729 16609 21741 16643
rect 21775 16640 21787 16643
rect 21775 16612 21864 16640
rect 21775 16609 21787 16612
rect 21729 16603 21787 16609
rect 9171 16544 9444 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 10410 16532 10416 16584
rect 10468 16572 10474 16584
rect 10505 16575 10563 16581
rect 10505 16572 10517 16575
rect 10468 16544 10517 16572
rect 10468 16532 10474 16544
rect 10505 16541 10517 16544
rect 10551 16541 10563 16575
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 10505 16535 10563 16541
rect 10888 16544 11161 16572
rect 2774 16464 2780 16516
rect 2832 16504 2838 16516
rect 3053 16507 3111 16513
rect 3053 16504 3065 16507
rect 2832 16476 3065 16504
rect 2832 16464 2838 16476
rect 3053 16473 3065 16476
rect 3099 16473 3111 16507
rect 3053 16467 3111 16473
rect 8021 16507 8079 16513
rect 8021 16473 8033 16507
rect 8067 16473 8079 16507
rect 8021 16467 8079 16473
rect 1762 16436 1768 16448
rect 1723 16408 1768 16436
rect 1762 16396 1768 16408
rect 1820 16396 1826 16448
rect 2409 16439 2467 16445
rect 2409 16405 2421 16439
rect 2455 16436 2467 16439
rect 2866 16436 2872 16448
rect 2455 16408 2872 16436
rect 2455 16405 2467 16408
rect 2409 16399 2467 16405
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 4065 16439 4123 16445
rect 4065 16436 4077 16439
rect 3384 16408 4077 16436
rect 3384 16396 3390 16408
rect 4065 16405 4077 16408
rect 4111 16405 4123 16439
rect 5718 16436 5724 16448
rect 5679 16408 5724 16436
rect 4065 16399 4123 16405
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 6914 16436 6920 16448
rect 6875 16408 6920 16436
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 7190 16396 7196 16448
rect 7248 16436 7254 16448
rect 8036 16436 8064 16467
rect 7248 16408 8064 16436
rect 7248 16396 7254 16408
rect 9674 16396 9680 16448
rect 9732 16436 9738 16448
rect 9769 16439 9827 16445
rect 9769 16436 9781 16439
rect 9732 16408 9781 16436
rect 9732 16396 9738 16408
rect 9769 16405 9781 16408
rect 9815 16405 9827 16439
rect 9769 16399 9827 16405
rect 10321 16439 10379 16445
rect 10321 16405 10333 16439
rect 10367 16436 10379 16439
rect 10888 16436 10916 16544
rect 11149 16541 11161 16544
rect 11195 16541 11207 16575
rect 11790 16572 11796 16584
rect 11751 16544 11796 16572
rect 11149 16535 11207 16541
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 13078 16572 13084 16584
rect 13039 16544 13084 16572
rect 12437 16535 12495 16541
rect 12452 16504 12480 16535
rect 13078 16532 13084 16544
rect 13136 16532 13142 16584
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 13725 16575 13783 16581
rect 13725 16572 13737 16575
rect 13688 16544 13737 16572
rect 13688 16532 13694 16544
rect 13725 16541 13737 16544
rect 13771 16541 13783 16575
rect 13725 16535 13783 16541
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 12986 16504 12992 16516
rect 12452 16476 12992 16504
rect 12986 16464 12992 16476
rect 13044 16464 13050 16516
rect 14936 16504 14964 16535
rect 16850 16532 16856 16584
rect 16908 16572 16914 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16908 16544 16957 16572
rect 16908 16532 16914 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 17586 16572 17592 16584
rect 16945 16535 17003 16541
rect 17052 16544 17592 16572
rect 13556 16476 14964 16504
rect 10367 16408 10916 16436
rect 10367 16405 10379 16408
rect 10321 16399 10379 16405
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 13556 16445 13584 16476
rect 15562 16464 15568 16516
rect 15620 16504 15626 16516
rect 15620 16476 15665 16504
rect 15620 16464 15626 16476
rect 15746 16464 15752 16516
rect 15804 16504 15810 16516
rect 16758 16504 16764 16516
rect 15804 16476 16764 16504
rect 15804 16464 15810 16476
rect 16758 16464 16764 16476
rect 16816 16504 16822 16516
rect 17052 16504 17080 16544
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 18693 16575 18751 16581
rect 18693 16541 18705 16575
rect 18739 16572 18751 16575
rect 19334 16572 19340 16584
rect 18739 16544 19340 16572
rect 18739 16541 18751 16544
rect 18693 16535 18751 16541
rect 18248 16504 18276 16535
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 16816 16476 17080 16504
rect 17420 16476 18276 16504
rect 19613 16507 19671 16513
rect 16816 16464 16822 16476
rect 12253 16439 12311 16445
rect 12253 16436 12265 16439
rect 11848 16408 12265 16436
rect 11848 16396 11854 16408
rect 12253 16405 12265 16408
rect 12299 16405 12311 16439
rect 12253 16399 12311 16405
rect 13541 16439 13599 16445
rect 13541 16405 13553 16439
rect 13587 16405 13599 16439
rect 14734 16436 14740 16448
rect 14695 16408 14740 16436
rect 13541 16399 13599 16405
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 17420 16445 17448 16476
rect 19613 16473 19625 16507
rect 19659 16473 19671 16507
rect 21836 16504 21864 16612
rect 21928 16581 21956 16680
rect 23477 16677 23489 16680
rect 23523 16677 23535 16711
rect 23477 16671 23535 16677
rect 22848 16640 23060 16652
rect 33226 16640 33232 16652
rect 22112 16624 33232 16640
rect 22112 16612 22876 16624
rect 23032 16612 33232 16624
rect 21913 16575 21971 16581
rect 21913 16541 21925 16575
rect 21959 16541 21971 16575
rect 22112 16572 22140 16612
rect 33226 16600 33232 16612
rect 33284 16600 33290 16652
rect 21913 16535 21971 16541
rect 22066 16544 22140 16572
rect 23017 16575 23075 16581
rect 22066 16504 22094 16544
rect 23017 16541 23029 16575
rect 23063 16572 23075 16575
rect 23474 16572 23480 16584
rect 23063 16544 23480 16572
rect 23063 16541 23075 16544
rect 23017 16535 23075 16541
rect 23474 16532 23480 16544
rect 23532 16532 23538 16584
rect 23658 16572 23664 16584
rect 23619 16544 23664 16572
rect 23658 16532 23664 16544
rect 23716 16532 23722 16584
rect 21836 16476 22094 16504
rect 19613 16467 19671 16473
rect 17405 16439 17463 16445
rect 17405 16405 17417 16439
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 18049 16439 18107 16445
rect 18049 16405 18061 16439
rect 18095 16436 18107 16439
rect 19426 16436 19432 16448
rect 18095 16408 19432 16436
rect 18095 16405 18107 16408
rect 18049 16399 18107 16405
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 19628 16436 19656 16467
rect 20070 16436 20076 16448
rect 19628 16408 20076 16436
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20898 16396 20904 16448
rect 20956 16436 20962 16448
rect 21269 16439 21327 16445
rect 21269 16436 21281 16439
rect 20956 16408 21281 16436
rect 20956 16396 20962 16408
rect 21269 16405 21281 16408
rect 21315 16436 21327 16439
rect 22373 16439 22431 16445
rect 22373 16436 22385 16439
rect 21315 16408 22385 16436
rect 21315 16405 21327 16408
rect 21269 16399 21327 16405
rect 22373 16405 22385 16408
rect 22419 16405 22431 16439
rect 22373 16399 22431 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 5166 16192 5172 16244
rect 5224 16232 5230 16244
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 5224 16204 5365 16232
rect 5224 16192 5230 16204
rect 5353 16201 5365 16204
rect 5399 16201 5411 16235
rect 5353 16195 5411 16201
rect 5718 16192 5724 16244
rect 5776 16232 5782 16244
rect 9677 16235 9735 16241
rect 5776 16204 9076 16232
rect 5776 16192 5782 16204
rect 2958 16124 2964 16176
rect 3016 16164 3022 16176
rect 5258 16164 5264 16176
rect 3016 16136 5264 16164
rect 3016 16124 3022 16136
rect 1949 16099 2007 16105
rect 1949 16065 1961 16099
rect 1995 16096 2007 16099
rect 2038 16096 2044 16108
rect 1995 16068 2044 16096
rect 1995 16065 2007 16068
rect 1949 16059 2007 16065
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 2406 16056 2412 16108
rect 2464 16096 2470 16108
rect 3160 16105 3188 16136
rect 5258 16124 5264 16136
rect 5316 16124 5322 16176
rect 7006 16124 7012 16176
rect 7064 16164 7070 16176
rect 7745 16167 7803 16173
rect 7064 16136 7696 16164
rect 7064 16124 7070 16136
rect 2501 16099 2559 16105
rect 2501 16096 2513 16099
rect 2464 16068 2513 16096
rect 2464 16056 2470 16068
rect 2501 16065 2513 16068
rect 2547 16065 2559 16099
rect 2501 16059 2559 16065
rect 3145 16099 3203 16105
rect 3145 16065 3157 16099
rect 3191 16065 3203 16099
rect 4430 16096 4436 16108
rect 4391 16068 4436 16096
rect 3145 16059 3203 16065
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 5534 16096 5540 16108
rect 5495 16068 5540 16096
rect 5534 16056 5540 16068
rect 5592 16056 5598 16108
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16096 7251 16099
rect 7282 16096 7288 16108
rect 7239 16068 7288 16096
rect 7239 16065 7251 16068
rect 7193 16059 7251 16065
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 7668 16105 7696 16136
rect 7745 16133 7757 16167
rect 7791 16164 7803 16167
rect 8481 16167 8539 16173
rect 8481 16164 8493 16167
rect 7791 16136 8493 16164
rect 7791 16133 7803 16136
rect 7745 16127 7803 16133
rect 8481 16133 8493 16136
rect 8527 16133 8539 16167
rect 8481 16127 8539 16133
rect 7653 16099 7711 16105
rect 7653 16065 7665 16099
rect 7699 16096 7711 16099
rect 7834 16096 7840 16108
rect 7699 16068 7840 16096
rect 7699 16065 7711 16068
rect 7653 16059 7711 16065
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 3789 16031 3847 16037
rect 3789 15997 3801 16031
rect 3835 16028 3847 16031
rect 3970 16028 3976 16040
rect 3835 16000 3976 16028
rect 3835 15997 3847 16000
rect 3789 15991 3847 15997
rect 3970 15988 3976 16000
rect 4028 15988 4034 16040
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 16028 8447 16031
rect 8435 16000 8616 16028
rect 8435 15997 8447 16000
rect 8389 15991 8447 15997
rect 1486 15852 1492 15904
rect 1544 15892 1550 15904
rect 1765 15895 1823 15901
rect 1765 15892 1777 15895
rect 1544 15864 1777 15892
rect 1544 15852 1550 15864
rect 1765 15861 1777 15864
rect 1811 15861 1823 15895
rect 1765 15855 1823 15861
rect 2593 15895 2651 15901
rect 2593 15861 2605 15895
rect 2639 15892 2651 15895
rect 2682 15892 2688 15904
rect 2639 15864 2688 15892
rect 2639 15861 2651 15864
rect 2593 15855 2651 15861
rect 2682 15852 2688 15864
rect 2740 15852 2746 15904
rect 3237 15895 3295 15901
rect 3237 15861 3249 15895
rect 3283 15892 3295 15895
rect 3510 15892 3516 15904
rect 3283 15864 3516 15892
rect 3283 15861 3295 15864
rect 3237 15855 3295 15861
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 4525 15895 4583 15901
rect 4525 15861 4537 15895
rect 4571 15892 4583 15895
rect 5626 15892 5632 15904
rect 4571 15864 5632 15892
rect 4571 15861 4583 15864
rect 4525 15855 4583 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 7009 15895 7067 15901
rect 7009 15861 7021 15895
rect 7055 15892 7067 15895
rect 8018 15892 8024 15904
rect 7055 15864 8024 15892
rect 7055 15861 7067 15864
rect 7009 15855 7067 15861
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 8588 15892 8616 16000
rect 8662 15988 8668 16040
rect 8720 16028 8726 16040
rect 8720 16000 8765 16028
rect 8720 15988 8726 16000
rect 9048 15960 9076 16204
rect 9677 16201 9689 16235
rect 9723 16232 9735 16235
rect 9766 16232 9772 16244
rect 9723 16204 9772 16232
rect 9723 16201 9735 16204
rect 9677 16195 9735 16201
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 10778 16192 10784 16244
rect 10836 16232 10842 16244
rect 10836 16204 12434 16232
rect 10836 16192 10842 16204
rect 9306 16124 9312 16176
rect 9364 16164 9370 16176
rect 10597 16167 10655 16173
rect 10597 16164 10609 16167
rect 9364 16136 10609 16164
rect 9364 16124 9370 16136
rect 10597 16133 10609 16136
rect 10643 16133 10655 16167
rect 10597 16127 10655 16133
rect 10870 16124 10876 16176
rect 10928 16164 10934 16176
rect 11149 16167 11207 16173
rect 11149 16164 11161 16167
rect 10928 16136 11161 16164
rect 10928 16124 10934 16136
rect 11149 16133 11161 16136
rect 11195 16133 11207 16167
rect 12406 16164 12434 16204
rect 12618 16192 12624 16244
rect 12676 16232 12682 16244
rect 12713 16235 12771 16241
rect 12713 16232 12725 16235
rect 12676 16204 12725 16232
rect 12676 16192 12682 16204
rect 12713 16201 12725 16204
rect 12759 16201 12771 16235
rect 21174 16232 21180 16244
rect 12713 16195 12771 16201
rect 13280 16204 20760 16232
rect 21135 16204 21180 16232
rect 13280 16164 13308 16204
rect 12406 16136 13308 16164
rect 14921 16167 14979 16173
rect 11149 16127 11207 16133
rect 9858 16096 9864 16108
rect 9819 16068 9864 16096
rect 9858 16056 9864 16068
rect 9916 16056 9922 16108
rect 12342 16096 12348 16108
rect 12303 16068 12348 16096
rect 12342 16056 12348 16068
rect 12400 16056 12406 16108
rect 12636 16105 12664 16136
rect 14921 16133 14933 16167
rect 14967 16164 14979 16167
rect 18693 16167 18751 16173
rect 18693 16164 18705 16167
rect 14967 16136 18705 16164
rect 14967 16133 14979 16136
rect 14921 16127 14979 16133
rect 18693 16133 18705 16136
rect 18739 16133 18751 16167
rect 18693 16127 18751 16133
rect 19613 16167 19671 16173
rect 19613 16133 19625 16167
rect 19659 16164 19671 16167
rect 20622 16164 20628 16176
rect 19659 16136 20628 16164
rect 19659 16133 19671 16136
rect 19613 16127 19671 16133
rect 20622 16124 20628 16136
rect 20680 16124 20686 16176
rect 20732 16164 20760 16204
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 22741 16235 22799 16241
rect 22741 16201 22753 16235
rect 22787 16232 22799 16235
rect 23014 16232 23020 16244
rect 22787 16204 23020 16232
rect 22787 16201 22799 16204
rect 22741 16195 22799 16201
rect 23014 16192 23020 16204
rect 23072 16192 23078 16244
rect 23106 16192 23112 16244
rect 23164 16232 23170 16244
rect 23201 16235 23259 16241
rect 23201 16232 23213 16235
rect 23164 16204 23213 16232
rect 23164 16192 23170 16204
rect 23201 16201 23213 16204
rect 23247 16201 23259 16235
rect 23201 16195 23259 16201
rect 21726 16164 21732 16176
rect 20732 16136 21732 16164
rect 21726 16124 21732 16136
rect 21784 16124 21790 16176
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16065 12679 16099
rect 12621 16059 12679 16065
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13633 16099 13691 16105
rect 13633 16096 13645 16099
rect 13412 16068 13645 16096
rect 13412 16056 13418 16068
rect 13633 16065 13645 16068
rect 13679 16065 13691 16099
rect 13633 16059 13691 16065
rect 14829 16099 14887 16105
rect 14829 16065 14841 16099
rect 14875 16065 14887 16099
rect 15654 16096 15660 16108
rect 15615 16068 15660 16096
rect 14829 16059 14887 16065
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 16028 10563 16031
rect 11606 16028 11612 16040
rect 10551 16000 11612 16028
rect 10551 15997 10563 16000
rect 10505 15991 10563 15997
rect 11606 15988 11612 16000
rect 11664 15988 11670 16040
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 16028 13231 16031
rect 13446 16028 13452 16040
rect 13219 16000 13452 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 14844 16028 14872 16059
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 17862 16096 17868 16108
rect 16163 16068 17868 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 17862 16056 17868 16068
rect 17920 16056 17926 16108
rect 20898 16096 20904 16108
rect 19536 16068 20904 16096
rect 13648 16000 14872 16028
rect 16853 16031 16911 16037
rect 13648 15972 13676 16000
rect 16853 15997 16865 16031
rect 16899 16028 16911 16031
rect 16942 16028 16948 16040
rect 16899 16000 16948 16028
rect 16899 15997 16911 16000
rect 16853 15991 16911 15997
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 17037 16031 17095 16037
rect 17037 15997 17049 16031
rect 17083 16028 17095 16031
rect 18601 16031 18659 16037
rect 17083 16000 17172 16028
rect 17083 15997 17095 16000
rect 17037 15991 17095 15997
rect 12434 15960 12440 15972
rect 9048 15932 12440 15960
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 13630 15920 13636 15972
rect 13688 15920 13694 15972
rect 15473 15963 15531 15969
rect 15473 15929 15485 15963
rect 15519 15960 15531 15963
rect 16666 15960 16672 15972
rect 15519 15932 16672 15960
rect 15519 15929 15531 15932
rect 15473 15923 15531 15929
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 17144 15960 17172 16000
rect 18601 15997 18613 16031
rect 18647 16028 18659 16031
rect 19536 16028 19564 16068
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 21542 16056 21548 16108
rect 21600 16096 21606 16108
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 21600 16068 23397 16096
rect 21600 16056 21606 16068
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23842 16096 23848 16108
rect 23803 16068 23848 16096
rect 23385 16059 23443 16065
rect 23842 16056 23848 16068
rect 23900 16056 23906 16108
rect 34149 16099 34207 16105
rect 34149 16065 34161 16099
rect 34195 16096 34207 16099
rect 38102 16096 38108 16108
rect 34195 16068 38108 16096
rect 34195 16065 34207 16068
rect 34149 16059 34207 16065
rect 38102 16056 38108 16068
rect 38160 16056 38166 16108
rect 18647 16000 19564 16028
rect 20073 16031 20131 16037
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 20073 15997 20085 16031
rect 20119 15997 20131 16031
rect 20073 15991 20131 15997
rect 20257 16031 20315 16037
rect 20257 15997 20269 16031
rect 20303 16028 20315 16031
rect 20806 16028 20812 16040
rect 20303 16000 20812 16028
rect 20303 15997 20315 16000
rect 20257 15991 20315 15997
rect 16776 15932 17172 15960
rect 9950 15892 9956 15904
rect 8588 15864 9956 15892
rect 9950 15852 9956 15864
rect 10008 15892 10014 15904
rect 10686 15892 10692 15904
rect 10008 15864 10692 15892
rect 10008 15852 10014 15864
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 12161 15895 12219 15901
rect 12161 15861 12173 15895
rect 12207 15892 12219 15895
rect 12618 15892 12624 15904
rect 12207 15864 12624 15892
rect 12207 15861 12219 15864
rect 12161 15855 12219 15861
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 13170 15852 13176 15904
rect 13228 15892 13234 15904
rect 13817 15895 13875 15901
rect 13817 15892 13829 15895
rect 13228 15864 13829 15892
rect 13228 15852 13234 15864
rect 13817 15861 13829 15864
rect 13863 15861 13875 15895
rect 13817 15855 13875 15861
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 16776 15892 16804 15932
rect 17494 15920 17500 15972
rect 17552 15960 17558 15972
rect 19610 15960 19616 15972
rect 17552 15932 19616 15960
rect 17552 15920 17558 15932
rect 19610 15920 19616 15932
rect 19668 15920 19674 15972
rect 20088 15960 20116 15991
rect 20806 15988 20812 16000
rect 20864 15988 20870 16040
rect 22097 16031 22155 16037
rect 22097 15997 22109 16031
rect 22143 15997 22155 16031
rect 22097 15991 22155 15997
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 16028 22339 16031
rect 23937 16031 23995 16037
rect 23937 16028 23949 16031
rect 22327 16000 23949 16028
rect 22327 15997 22339 16000
rect 22281 15991 22339 15997
rect 23937 15997 23949 16000
rect 23983 15997 23995 16031
rect 23937 15991 23995 15997
rect 22112 15960 22140 15991
rect 34241 15963 34299 15969
rect 34241 15960 34253 15963
rect 20088 15932 21128 15960
rect 22112 15932 34253 15960
rect 17218 15892 17224 15904
rect 14608 15864 16804 15892
rect 17179 15864 17224 15892
rect 14608 15852 14614 15864
rect 17218 15852 17224 15864
rect 17276 15852 17282 15904
rect 20438 15892 20444 15904
rect 20399 15864 20444 15892
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 21100 15892 21128 15932
rect 34241 15929 34253 15932
rect 34287 15929 34299 15963
rect 34241 15923 34299 15929
rect 23106 15892 23112 15904
rect 21100 15864 23112 15892
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 7190 15688 7196 15700
rect 7151 15660 7196 15688
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 9306 15688 9312 15700
rect 9267 15660 9312 15688
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 10744 15660 11069 15688
rect 10744 15648 10750 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 11057 15651 11115 15657
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 12621 15691 12679 15697
rect 12621 15688 12633 15691
rect 12584 15660 12633 15688
rect 12584 15648 12590 15660
rect 12621 15657 12633 15660
rect 12667 15688 12679 15691
rect 13170 15688 13176 15700
rect 12667 15660 13176 15688
rect 12667 15657 12679 15660
rect 12621 15651 12679 15657
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 14553 15691 14611 15697
rect 14553 15657 14565 15691
rect 14599 15688 14611 15691
rect 15562 15688 15568 15700
rect 14599 15660 15568 15688
rect 14599 15657 14611 15660
rect 14553 15651 14611 15657
rect 15562 15648 15568 15660
rect 15620 15648 15626 15700
rect 17129 15691 17187 15697
rect 17129 15657 17141 15691
rect 17175 15688 17187 15691
rect 17218 15688 17224 15700
rect 17175 15660 17224 15688
rect 17175 15657 17187 15660
rect 17129 15651 17187 15657
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 22833 15691 22891 15697
rect 17328 15660 22094 15688
rect 1581 15623 1639 15629
rect 1581 15589 1593 15623
rect 1627 15620 1639 15623
rect 7098 15620 7104 15632
rect 1627 15592 7104 15620
rect 1627 15589 1639 15592
rect 1581 15583 1639 15589
rect 7098 15580 7104 15592
rect 7156 15580 7162 15632
rect 8478 15620 8484 15632
rect 8439 15592 8484 15620
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 13446 15580 13452 15632
rect 13504 15620 13510 15632
rect 17328 15620 17356 15660
rect 21450 15620 21456 15632
rect 13504 15592 17356 15620
rect 19536 15592 21456 15620
rect 13504 15580 13510 15592
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15552 7987 15555
rect 9674 15552 9680 15564
rect 7975 15524 9680 15552
rect 7975 15521 7987 15524
rect 7929 15515 7987 15521
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15552 10011 15555
rect 12161 15555 12219 15561
rect 12161 15552 12173 15555
rect 9999 15524 12173 15552
rect 9999 15521 10011 15524
rect 9953 15515 10011 15521
rect 12161 15521 12173 15524
rect 12207 15521 12219 15555
rect 12161 15515 12219 15521
rect 12618 15512 12624 15564
rect 12676 15552 12682 15564
rect 13265 15555 13323 15561
rect 13265 15552 13277 15555
rect 12676 15524 13277 15552
rect 12676 15512 12682 15524
rect 13265 15521 13277 15524
rect 13311 15521 13323 15555
rect 13265 15515 13323 15521
rect 15010 15512 15016 15564
rect 15068 15552 15074 15564
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 15068 15524 15301 15552
rect 15068 15512 15074 15524
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 16206 15512 16212 15564
rect 16264 15552 16270 15564
rect 19536 15561 19564 15592
rect 21450 15580 21456 15592
rect 21508 15580 21514 15632
rect 22066 15620 22094 15660
rect 22833 15657 22845 15691
rect 22879 15688 22891 15691
rect 23658 15688 23664 15700
rect 22879 15660 23664 15688
rect 22879 15657 22891 15660
rect 22833 15651 22891 15657
rect 23658 15648 23664 15660
rect 23716 15648 23722 15700
rect 35069 15691 35127 15697
rect 35069 15657 35081 15691
rect 35115 15688 35127 15691
rect 35894 15688 35900 15700
rect 35115 15660 35900 15688
rect 35115 15657 35127 15660
rect 35069 15651 35127 15657
rect 35894 15648 35900 15660
rect 35952 15648 35958 15700
rect 38102 15688 38108 15700
rect 38063 15660 38108 15688
rect 38102 15648 38108 15660
rect 38160 15648 38166 15700
rect 32398 15620 32404 15632
rect 22066 15592 32404 15620
rect 32398 15580 32404 15592
rect 32456 15580 32462 15632
rect 18325 15555 18383 15561
rect 18325 15552 18337 15555
rect 16264 15524 18337 15552
rect 16264 15512 16270 15524
rect 18325 15521 18337 15524
rect 18371 15521 18383 15555
rect 18325 15515 18383 15521
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15521 19579 15555
rect 19521 15515 19579 15521
rect 19610 15512 19616 15564
rect 19668 15552 19674 15564
rect 21085 15555 21143 15561
rect 19668 15524 20668 15552
rect 19668 15512 19674 15524
rect 1762 15484 1768 15496
rect 1723 15456 1768 15484
rect 1762 15444 1768 15456
rect 1820 15444 1826 15496
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 2590 15484 2596 15496
rect 2455 15456 2596 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 3237 15487 3295 15493
rect 3237 15453 3249 15487
rect 3283 15484 3295 15487
rect 3602 15484 3608 15496
rect 3283 15456 3608 15484
rect 3283 15453 3295 15456
rect 3237 15447 3295 15453
rect 3602 15444 3608 15456
rect 3660 15444 3666 15496
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15484 4583 15487
rect 5166 15484 5172 15496
rect 4571 15456 5172 15484
rect 4571 15453 4583 15456
rect 4525 15447 4583 15453
rect 5166 15444 5172 15456
rect 5224 15444 5230 15496
rect 5350 15484 5356 15496
rect 5311 15456 5356 15484
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 6181 15487 6239 15493
rect 6181 15453 6193 15487
rect 6227 15484 6239 15487
rect 7006 15484 7012 15496
rect 6227 15456 7012 15484
rect 6227 15453 6239 15456
rect 6181 15447 6239 15453
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 7374 15484 7380 15496
rect 7335 15456 7380 15484
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15484 9275 15487
rect 9766 15484 9772 15496
rect 9263 15456 9772 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15484 9919 15487
rect 10410 15484 10416 15496
rect 9907 15456 10416 15484
rect 9907 15453 9919 15456
rect 9861 15447 9919 15453
rect 8021 15419 8079 15425
rect 8021 15385 8033 15419
rect 8067 15416 8079 15419
rect 8386 15416 8392 15428
rect 8067 15388 8392 15416
rect 8067 15385 8079 15388
rect 8021 15379 8079 15385
rect 8386 15376 8392 15388
rect 8444 15376 8450 15428
rect 9674 15376 9680 15428
rect 9732 15416 9738 15428
rect 9876 15416 9904 15447
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 9732 15388 9904 15416
rect 10520 15416 10548 15447
rect 10594 15444 10600 15496
rect 10652 15484 10658 15496
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10652 15456 10701 15484
rect 10652 15444 10658 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 11977 15487 12035 15493
rect 11977 15453 11989 15487
rect 12023 15484 12035 15487
rect 12066 15484 12072 15496
rect 12023 15456 12072 15484
rect 12023 15453 12035 15456
rect 11977 15447 12035 15453
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 12710 15444 12716 15496
rect 12768 15484 12774 15496
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 12768 15456 13093 15484
rect 12768 15444 12774 15456
rect 13081 15453 13093 15456
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 13170 15444 13176 15496
rect 13228 15484 13234 15496
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 13228 15456 14473 15484
rect 13228 15444 13234 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 15105 15487 15163 15493
rect 15105 15484 15117 15487
rect 14461 15447 14519 15453
rect 14660 15456 15117 15484
rect 14660 15416 14688 15456
rect 15105 15453 15117 15456
rect 15151 15484 15163 15487
rect 16298 15484 16304 15496
rect 15151 15456 16304 15484
rect 15151 15453 15163 15456
rect 15105 15447 15163 15453
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 16482 15484 16488 15496
rect 16443 15456 16488 15484
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 16666 15484 16672 15496
rect 16627 15456 16672 15484
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 16942 15444 16948 15496
rect 17000 15484 17006 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 17000 15456 18153 15484
rect 17000 15444 17006 15456
rect 18141 15453 18153 15456
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 10520 15388 14688 15416
rect 9732 15376 9738 15388
rect 14734 15376 14740 15428
rect 14792 15416 14798 15428
rect 19613 15419 19671 15425
rect 19613 15416 19625 15419
rect 14792 15388 19625 15416
rect 14792 15376 14798 15388
rect 19613 15385 19625 15388
rect 19659 15385 19671 15419
rect 19613 15379 19671 15385
rect 20533 15419 20591 15425
rect 20533 15385 20545 15419
rect 20579 15385 20591 15419
rect 20640 15416 20668 15524
rect 21085 15521 21097 15555
rect 21131 15552 21143 15555
rect 22189 15555 22247 15561
rect 22189 15552 22201 15555
rect 21131 15524 22201 15552
rect 21131 15521 21143 15524
rect 21085 15515 21143 15521
rect 22189 15521 22201 15524
rect 22235 15521 22247 15555
rect 22189 15515 22247 15521
rect 22554 15512 22560 15564
rect 22612 15552 22618 15564
rect 22612 15524 23060 15552
rect 22612 15512 22618 15524
rect 21269 15487 21327 15493
rect 21269 15453 21281 15487
rect 21315 15484 21327 15487
rect 22922 15484 22928 15496
rect 21315 15456 22928 15484
rect 21315 15453 21327 15456
rect 21269 15447 21327 15453
rect 22922 15444 22928 15456
rect 22980 15444 22986 15496
rect 23032 15493 23060 15524
rect 23106 15512 23112 15564
rect 23164 15552 23170 15564
rect 33134 15552 33140 15564
rect 23164 15524 33140 15552
rect 23164 15512 23170 15524
rect 33134 15512 33140 15524
rect 33192 15512 33198 15564
rect 23017 15487 23075 15493
rect 23017 15453 23029 15487
rect 23063 15484 23075 15487
rect 23661 15487 23719 15493
rect 23661 15484 23673 15487
rect 23063 15456 23673 15484
rect 23063 15453 23075 15456
rect 23017 15447 23075 15453
rect 23661 15453 23673 15456
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 31938 15444 31944 15496
rect 31996 15484 32002 15496
rect 35253 15487 35311 15493
rect 35253 15484 35265 15487
rect 31996 15456 35265 15484
rect 31996 15444 32002 15456
rect 35253 15453 35265 15456
rect 35299 15453 35311 15487
rect 38286 15484 38292 15496
rect 38247 15456 38292 15484
rect 35253 15447 35311 15453
rect 38286 15444 38292 15456
rect 38344 15444 38350 15496
rect 24578 15416 24584 15428
rect 20640 15388 24584 15416
rect 20533 15379 20591 15385
rect 2501 15351 2559 15357
rect 2501 15317 2513 15351
rect 2547 15348 2559 15351
rect 2682 15348 2688 15360
rect 2547 15320 2688 15348
rect 2547 15317 2559 15320
rect 2501 15311 2559 15317
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 3050 15348 3056 15360
rect 3011 15320 3056 15348
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 4614 15348 4620 15360
rect 4575 15320 4620 15348
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 4798 15308 4804 15360
rect 4856 15348 4862 15360
rect 5169 15351 5227 15357
rect 5169 15348 5181 15351
rect 4856 15320 5181 15348
rect 4856 15308 4862 15320
rect 5169 15317 5181 15320
rect 5215 15317 5227 15351
rect 6270 15348 6276 15360
rect 6231 15320 6276 15348
rect 5169 15311 5227 15317
rect 6270 15308 6276 15320
rect 6328 15308 6334 15360
rect 7834 15308 7840 15360
rect 7892 15348 7898 15360
rect 11330 15348 11336 15360
rect 7892 15320 11336 15348
rect 7892 15308 7898 15320
rect 11330 15308 11336 15320
rect 11388 15308 11394 15360
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 13630 15348 13636 15360
rect 13228 15320 13636 15348
rect 13228 15308 13234 15320
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 13725 15351 13783 15357
rect 13725 15317 13737 15351
rect 13771 15348 13783 15351
rect 15749 15351 15807 15357
rect 15749 15348 15761 15351
rect 13771 15320 15761 15348
rect 13771 15317 13783 15320
rect 13725 15311 13783 15317
rect 15749 15317 15761 15320
rect 15795 15348 15807 15351
rect 17034 15348 17040 15360
rect 15795 15320 17040 15348
rect 15795 15317 15807 15320
rect 15749 15311 15807 15317
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 18785 15351 18843 15357
rect 18785 15317 18797 15351
rect 18831 15348 18843 15351
rect 20254 15348 20260 15360
rect 18831 15320 20260 15348
rect 18831 15317 18843 15320
rect 18785 15311 18843 15317
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 20548 15348 20576 15379
rect 24578 15376 24584 15388
rect 24636 15376 24642 15428
rect 20622 15348 20628 15360
rect 20548 15320 20628 15348
rect 20622 15308 20628 15320
rect 20680 15308 20686 15360
rect 23474 15348 23480 15360
rect 23435 15320 23480 15348
rect 23474 15308 23480 15320
rect 23532 15308 23538 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 3145 15147 3203 15153
rect 3145 15113 3157 15147
rect 3191 15113 3203 15147
rect 3145 15107 3203 15113
rect 5077 15147 5135 15153
rect 5077 15113 5089 15147
rect 5123 15144 5135 15147
rect 5350 15144 5356 15156
rect 5123 15116 5356 15144
rect 5123 15113 5135 15116
rect 5077 15107 5135 15113
rect 3160 15076 3188 15107
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 7193 15147 7251 15153
rect 7193 15113 7205 15147
rect 7239 15144 7251 15147
rect 7374 15144 7380 15156
rect 7239 15116 7380 15144
rect 7239 15113 7251 15116
rect 7193 15107 7251 15113
rect 7374 15104 7380 15116
rect 7432 15104 7438 15156
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7616 15116 7849 15144
rect 7616 15104 7622 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 8386 15104 8392 15156
rect 8444 15144 8450 15156
rect 8573 15147 8631 15153
rect 8573 15144 8585 15147
rect 8444 15116 8585 15144
rect 8444 15104 8450 15116
rect 8573 15113 8585 15116
rect 8619 15113 8631 15147
rect 12526 15144 12532 15156
rect 8573 15107 8631 15113
rect 10428 15116 12532 15144
rect 6270 15076 6276 15088
rect 3160 15048 4016 15076
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 1857 15011 1915 15017
rect 1857 15008 1869 15011
rect 1636 14980 1869 15008
rect 1636 14968 1642 14980
rect 1857 14977 1869 14980
rect 1903 14977 1915 15011
rect 1857 14971 1915 14977
rect 2130 14968 2136 15020
rect 2188 15008 2194 15020
rect 2685 15011 2743 15017
rect 2685 15008 2697 15011
rect 2188 14980 2697 15008
rect 2188 14968 2194 14980
rect 2685 14977 2697 14980
rect 2731 14977 2743 15011
rect 2685 14971 2743 14977
rect 3142 14968 3148 15020
rect 3200 15008 3206 15020
rect 3988 15017 4016 15048
rect 4632 15048 6276 15076
rect 4632 15017 4660 15048
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 3329 15011 3387 15017
rect 3329 15008 3341 15011
rect 3200 14980 3341 15008
rect 3200 14968 3206 14980
rect 3329 14977 3341 14980
rect 3375 14977 3387 15011
rect 3329 14971 3387 14977
rect 3973 15011 4031 15017
rect 3973 14977 3985 15011
rect 4019 14977 4031 15011
rect 3973 14971 4031 14977
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 5166 14968 5172 15020
rect 5224 15008 5230 15020
rect 5261 15011 5319 15017
rect 5261 15008 5273 15011
rect 5224 14980 5273 15008
rect 5224 14968 5230 14980
rect 5261 14977 5273 14980
rect 5307 14977 5319 15011
rect 5261 14971 5319 14977
rect 5534 14968 5540 15020
rect 5592 15008 5598 15020
rect 5721 15011 5779 15017
rect 5721 15008 5733 15011
rect 5592 14980 5733 15008
rect 5592 14968 5598 14980
rect 5721 14977 5733 14980
rect 5767 14977 5779 15011
rect 5721 14971 5779 14977
rect 5736 14940 5764 14971
rect 5810 14968 5816 15020
rect 5868 15008 5874 15020
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 5868 14980 6745 15008
rect 5868 14968 5874 14980
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 8018 15008 8024 15020
rect 7979 14980 8024 15008
rect 7377 14971 7435 14977
rect 6270 14940 6276 14952
rect 5736 14912 6276 14940
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 7392 14940 7420 14971
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 8481 15011 8539 15017
rect 8481 14977 8493 15011
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 15008 9275 15011
rect 10428 15008 10456 15116
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 14550 15144 14556 15156
rect 13403 15116 14556 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 16206 15144 16212 15156
rect 16167 15116 16212 15144
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 16390 15104 16396 15156
rect 16448 15144 16454 15156
rect 16448 15116 17253 15144
rect 16448 15104 16454 15116
rect 11698 15036 11704 15088
rect 11756 15076 11762 15088
rect 14093 15079 14151 15085
rect 14093 15076 14105 15079
rect 11756 15048 14105 15076
rect 11756 15036 11762 15048
rect 14093 15045 14105 15048
rect 14139 15045 14151 15079
rect 17225 15076 17253 15116
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 20165 15147 20223 15153
rect 20165 15144 20177 15147
rect 19392 15116 20177 15144
rect 19392 15104 19398 15116
rect 20165 15113 20177 15116
rect 20211 15144 20223 15147
rect 20438 15144 20444 15156
rect 20211 15116 20444 15144
rect 20211 15113 20223 15116
rect 20165 15107 20223 15113
rect 20438 15104 20444 15116
rect 20496 15104 20502 15156
rect 21266 15144 21272 15156
rect 21227 15116 21272 15144
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 22922 15104 22928 15156
rect 22980 15144 22986 15156
rect 23109 15147 23167 15153
rect 23109 15144 23121 15147
rect 22980 15116 23121 15144
rect 22980 15104 22986 15116
rect 23109 15113 23121 15116
rect 23155 15113 23167 15147
rect 23109 15107 23167 15113
rect 17290 15079 17348 15085
rect 17290 15076 17302 15079
rect 17225 15048 17302 15076
rect 14093 15039 14151 15045
rect 17290 15045 17302 15048
rect 17336 15045 17348 15079
rect 17290 15039 17348 15045
rect 17494 15036 17500 15088
rect 17552 15076 17558 15088
rect 20714 15076 20720 15088
rect 17552 15048 20720 15076
rect 17552 15036 17558 15048
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 22554 15076 22560 15088
rect 21192 15048 22560 15076
rect 9263 14980 10456 15008
rect 10505 15011 10563 15017
rect 9263 14977 9275 14980
rect 9217 14971 9275 14977
rect 10505 14977 10517 15011
rect 10551 15008 10563 15011
rect 11149 15011 11207 15017
rect 10551 14980 11100 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 8496 14940 8524 14971
rect 9398 14940 9404 14952
rect 7392 14912 8524 14940
rect 9359 14912 9404 14940
rect 8496 14872 8524 14912
rect 9398 14900 9404 14912
rect 9456 14900 9462 14952
rect 10686 14940 10692 14952
rect 10647 14912 10692 14940
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 11072 14940 11100 14980
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 12805 15011 12863 15017
rect 12805 15008 12817 15011
rect 11195 14980 12817 15008
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 12805 14977 12817 14980
rect 12851 14977 12863 15011
rect 12805 14971 12863 14977
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 15008 13323 15011
rect 13814 15008 13820 15020
rect 13311 14980 13820 15008
rect 13311 14977 13323 14980
rect 13265 14971 13323 14977
rect 11882 14940 11888 14952
rect 11072 14912 11888 14940
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 12158 14940 12164 14952
rect 12119 14912 12164 14940
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 12314 14943 12372 14949
rect 12314 14909 12326 14943
rect 12360 14909 12372 14943
rect 12820 14940 12848 14971
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 15654 15008 15660 15020
rect 15567 14980 15660 15008
rect 15654 14968 15660 14980
rect 15712 15008 15718 15020
rect 16117 15011 16175 15017
rect 16117 15008 16129 15011
rect 15712 14980 16129 15008
rect 15712 14968 15718 14980
rect 16117 14977 16129 14980
rect 16163 15008 16175 15011
rect 16298 15008 16304 15020
rect 16163 14980 16304 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 18601 15011 18659 15017
rect 17920 14980 18552 15008
rect 17920 14968 17926 14980
rect 14001 14943 14059 14949
rect 14001 14940 14013 14943
rect 12820 14912 14013 14940
rect 12314 14903 12372 14909
rect 14001 14909 14013 14912
rect 14047 14909 14059 14943
rect 14001 14903 14059 14909
rect 10962 14872 10968 14884
rect 8496 14844 10968 14872
rect 10962 14832 10968 14844
rect 11020 14832 11026 14884
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 12329 14872 12357 14903
rect 17218 14900 17224 14952
rect 17276 14940 17282 14952
rect 18414 14940 18420 14952
rect 17276 14912 17321 14940
rect 18375 14912 18420 14940
rect 17276 14900 17282 14912
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 18524 14940 18552 14980
rect 18601 14977 18613 15011
rect 18647 15008 18659 15011
rect 20254 15008 20260 15020
rect 18647 14980 20260 15008
rect 18647 14977 18659 14980
rect 18601 14971 18659 14977
rect 20254 14968 20260 14980
rect 20312 14968 20318 15020
rect 21192 15017 21220 15048
rect 22554 15036 22560 15048
rect 22612 15036 22618 15088
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 14977 21235 15011
rect 21177 14971 21235 14977
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 15008 22063 15011
rect 23293 15011 23351 15017
rect 22051 14980 23244 15008
rect 22051 14977 22063 14980
rect 22005 14971 22063 14977
rect 19521 14943 19579 14949
rect 19521 14940 19533 14943
rect 18524 14912 19533 14940
rect 19521 14909 19533 14912
rect 19567 14909 19579 14943
rect 19521 14903 19579 14909
rect 19705 14943 19763 14949
rect 19705 14909 19717 14943
rect 19751 14940 19763 14943
rect 19978 14940 19984 14952
rect 19751 14912 19984 14940
rect 19751 14909 19763 14912
rect 19705 14903 19763 14909
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 22189 14943 22247 14949
rect 22189 14909 22201 14943
rect 22235 14940 22247 14943
rect 22646 14940 22652 14952
rect 22235 14912 22652 14940
rect 22235 14909 22247 14912
rect 22189 14903 22247 14909
rect 22646 14900 22652 14912
rect 22704 14900 22710 14952
rect 23216 14940 23244 14980
rect 23293 14977 23305 15011
rect 23339 15008 23351 15011
rect 23474 15008 23480 15020
rect 23339 14980 23480 15008
rect 23339 14977 23351 14980
rect 23293 14971 23351 14977
rect 23474 14968 23480 14980
rect 23532 14968 23538 15020
rect 33410 14940 33416 14952
rect 23216 14912 33416 14940
rect 33410 14900 33416 14912
rect 33468 14900 33474 14952
rect 11112 14844 12357 14872
rect 14553 14875 14611 14881
rect 11112 14832 11118 14844
rect 14553 14841 14565 14875
rect 14599 14872 14611 14875
rect 16574 14872 16580 14884
rect 14599 14844 16580 14872
rect 14599 14841 14611 14844
rect 14553 14835 14611 14841
rect 16574 14832 16580 14844
rect 16632 14832 16638 14884
rect 17678 14832 17684 14884
rect 17736 14872 17742 14884
rect 17773 14875 17831 14881
rect 17773 14872 17785 14875
rect 17736 14844 17785 14872
rect 17736 14832 17742 14844
rect 17773 14841 17785 14844
rect 17819 14841 17831 14875
rect 17773 14835 17831 14841
rect 19061 14875 19119 14881
rect 19061 14841 19073 14875
rect 19107 14872 19119 14875
rect 19426 14872 19432 14884
rect 19107 14844 19432 14872
rect 19107 14841 19119 14844
rect 19061 14835 19119 14841
rect 19426 14832 19432 14844
rect 19484 14872 19490 14884
rect 20162 14872 20168 14884
rect 19484 14844 20168 14872
rect 19484 14832 19490 14844
rect 20162 14832 20168 14844
rect 20220 14832 20226 14884
rect 21450 14832 21456 14884
rect 21508 14872 21514 14884
rect 22373 14875 22431 14881
rect 22373 14872 22385 14875
rect 21508 14844 22385 14872
rect 21508 14832 21514 14844
rect 22373 14841 22385 14844
rect 22419 14841 22431 14875
rect 22373 14835 22431 14841
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 2501 14807 2559 14813
rect 2501 14773 2513 14807
rect 2547 14804 2559 14807
rect 3418 14804 3424 14816
rect 2547 14776 3424 14804
rect 2547 14773 2559 14776
rect 2501 14767 2559 14773
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 3786 14804 3792 14816
rect 3747 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 4433 14807 4491 14813
rect 4433 14773 4445 14807
rect 4479 14804 4491 14807
rect 4706 14804 4712 14816
rect 4479 14776 4712 14804
rect 4479 14773 4491 14776
rect 4433 14767 4491 14773
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 5813 14807 5871 14813
rect 5813 14804 5825 14807
rect 5408 14776 5825 14804
rect 5408 14764 5414 14776
rect 5813 14773 5825 14776
rect 5859 14773 5871 14807
rect 5813 14767 5871 14773
rect 6549 14807 6607 14813
rect 6549 14773 6561 14807
rect 6595 14804 6607 14807
rect 6730 14804 6736 14816
rect 6595 14776 6736 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 8570 14764 8576 14816
rect 8628 14804 8634 14816
rect 9585 14807 9643 14813
rect 9585 14804 9597 14807
rect 8628 14776 9597 14804
rect 8628 14764 8634 14776
rect 9585 14773 9597 14776
rect 9631 14773 9643 14807
rect 9585 14767 9643 14773
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 12158 14804 12164 14816
rect 11204 14776 12164 14804
rect 11204 14764 11210 14776
rect 12158 14764 12164 14776
rect 12216 14764 12222 14816
rect 15473 14807 15531 14813
rect 15473 14773 15485 14807
rect 15519 14804 15531 14807
rect 17862 14804 17868 14816
rect 15519 14776 17868 14804
rect 15519 14773 15531 14776
rect 15473 14767 15531 14773
rect 17862 14764 17868 14776
rect 17920 14764 17926 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 2314 14560 2320 14612
rect 2372 14600 2378 14612
rect 2593 14603 2651 14609
rect 2593 14600 2605 14603
rect 2372 14572 2605 14600
rect 2372 14560 2378 14572
rect 2593 14569 2605 14572
rect 2639 14569 2651 14603
rect 2593 14563 2651 14569
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 10321 14603 10379 14609
rect 4580 14572 8708 14600
rect 4580 14560 4586 14572
rect 2682 14492 2688 14544
rect 2740 14532 2746 14544
rect 8478 14532 8484 14544
rect 2740 14504 4016 14532
rect 2740 14492 2746 14504
rect 3050 14464 3056 14476
rect 1596 14436 3056 14464
rect 1596 14405 1624 14436
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 3988 14473 4016 14504
rect 4080 14504 8484 14532
rect 3973 14467 4031 14473
rect 3973 14433 3985 14467
rect 4019 14433 4031 14467
rect 3973 14427 4031 14433
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14365 1639 14399
rect 1581 14359 1639 14365
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14365 2559 14399
rect 3418 14396 3424 14408
rect 3379 14368 3424 14396
rect 2501 14359 2559 14365
rect 2516 14328 2544 14359
rect 3418 14356 3424 14368
rect 3476 14356 3482 14408
rect 4080 14328 4108 14504
rect 8478 14492 8484 14504
rect 8536 14492 8542 14544
rect 8680 14532 8708 14572
rect 10321 14569 10333 14603
rect 10367 14600 10379 14603
rect 10686 14600 10692 14612
rect 10367 14572 10692 14600
rect 10367 14569 10379 14572
rect 10321 14563 10379 14569
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 11054 14600 11060 14612
rect 11015 14572 11060 14600
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11698 14600 11704 14612
rect 11659 14572 11704 14600
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 12253 14603 12311 14609
rect 12253 14569 12265 14603
rect 12299 14600 12311 14603
rect 12342 14600 12348 14612
rect 12299 14572 12348 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 12897 14603 12955 14609
rect 12897 14569 12909 14603
rect 12943 14600 12955 14603
rect 14826 14600 14832 14612
rect 12943 14572 14832 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 14826 14560 14832 14572
rect 14884 14560 14890 14612
rect 15010 14600 15016 14612
rect 14971 14572 15016 14600
rect 15010 14560 15016 14572
rect 15068 14560 15074 14612
rect 15102 14560 15108 14612
rect 15160 14600 15166 14612
rect 16850 14600 16856 14612
rect 15160 14572 16856 14600
rect 15160 14560 15166 14572
rect 16850 14560 16856 14572
rect 16908 14600 16914 14612
rect 17586 14600 17592 14612
rect 16908 14572 17592 14600
rect 16908 14560 16914 14572
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 17681 14603 17739 14609
rect 17681 14569 17693 14603
rect 17727 14600 17739 14603
rect 20070 14600 20076 14612
rect 17727 14572 20076 14600
rect 17727 14569 17739 14572
rect 17681 14563 17739 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20806 14600 20812 14612
rect 20767 14572 20812 14600
rect 20806 14560 20812 14572
rect 20864 14560 20870 14612
rect 22646 14600 22652 14612
rect 22607 14572 22652 14600
rect 22646 14560 22652 14572
rect 22704 14560 22710 14612
rect 28445 14603 28503 14609
rect 28445 14569 28457 14603
rect 28491 14600 28503 14603
rect 31938 14600 31944 14612
rect 28491 14572 31944 14600
rect 28491 14569 28503 14572
rect 28445 14563 28503 14569
rect 31938 14560 31944 14572
rect 31996 14560 32002 14612
rect 8680 14504 23244 14532
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14464 4215 14467
rect 4614 14464 4620 14476
rect 4203 14436 4620 14464
rect 4203 14433 4215 14436
rect 4157 14427 4215 14433
rect 4614 14424 4620 14436
rect 4672 14424 4678 14476
rect 4890 14424 4896 14476
rect 4948 14464 4954 14476
rect 5537 14467 5595 14473
rect 5537 14464 5549 14467
rect 4948 14436 5549 14464
rect 4948 14424 4954 14436
rect 5537 14433 5549 14436
rect 5583 14433 5595 14467
rect 8570 14464 8576 14476
rect 5537 14427 5595 14433
rect 7300 14436 8576 14464
rect 7300 14405 7328 14436
rect 8570 14424 8576 14436
rect 8628 14424 8634 14476
rect 12710 14464 12716 14476
rect 9876 14436 10732 14464
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 7285 14399 7343 14405
rect 7285 14365 7297 14399
rect 7331 14365 7343 14399
rect 7926 14396 7932 14408
rect 7887 14368 7932 14396
rect 7285 14359 7343 14365
rect 2516 14300 4108 14328
rect 4617 14331 4675 14337
rect 4617 14297 4629 14331
rect 4663 14328 4675 14331
rect 4890 14328 4896 14340
rect 4663 14300 4896 14328
rect 4663 14297 4675 14300
rect 4617 14291 4675 14297
rect 4890 14288 4896 14300
rect 4948 14328 4954 14340
rect 5261 14331 5319 14337
rect 5261 14328 5273 14331
rect 4948 14300 5273 14328
rect 4948 14288 4954 14300
rect 5261 14297 5273 14300
rect 5307 14297 5319 14331
rect 5261 14291 5319 14297
rect 5350 14288 5356 14340
rect 5408 14328 5414 14340
rect 6840 14328 6868 14359
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8110 14396 8116 14408
rect 8071 14368 8116 14396
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 9876 14405 9904 14436
rect 10704 14408 10732 14436
rect 12452 14436 12716 14464
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 9582 14328 9588 14340
rect 5408 14300 5453 14328
rect 6840 14300 9588 14328
rect 5408 14288 5414 14300
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 10520 14328 10548 14359
rect 10686 14356 10692 14408
rect 10744 14396 10750 14408
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 10744 14368 10977 14396
rect 10744 14356 10750 14368
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 11514 14356 11520 14408
rect 11572 14396 11578 14408
rect 12452 14405 12480 14436
rect 12710 14424 12716 14436
rect 12768 14464 12774 14476
rect 15565 14467 15623 14473
rect 12768 14436 14964 14464
rect 12768 14424 12774 14436
rect 14936 14408 14964 14436
rect 15565 14433 15577 14467
rect 15611 14464 15623 14467
rect 16482 14464 16488 14476
rect 15611 14436 16488 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 16632 14436 16957 14464
rect 16632 14424 16638 14436
rect 16945 14433 16957 14436
rect 16991 14464 17003 14467
rect 16991 14436 17724 14464
rect 16991 14433 17003 14436
rect 16945 14427 17003 14433
rect 11609 14399 11667 14405
rect 11609 14396 11621 14399
rect 11572 14368 11621 14396
rect 11572 14356 11578 14368
rect 11609 14365 11621 14368
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14365 12495 14399
rect 12437 14359 12495 14365
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14365 13139 14399
rect 13081 14359 13139 14365
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13906 14396 13912 14408
rect 13587 14368 13912 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 9692 14300 10548 14328
rect 13096 14328 13124 14359
rect 13906 14356 13912 14368
rect 13964 14396 13970 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 13964 14368 14473 14396
rect 13964 14356 13970 14368
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14918 14396 14924 14408
rect 14879 14368 14924 14396
rect 14461 14359 14519 14365
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 17586 14396 17592 14408
rect 17547 14368 17592 14396
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 17696 14396 17724 14436
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 18012 14436 18429 14464
rect 18012 14424 18018 14436
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 19613 14467 19671 14473
rect 19613 14433 19625 14467
rect 19659 14464 19671 14467
rect 19886 14464 19892 14476
rect 19659 14436 19892 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 19886 14424 19892 14436
rect 19944 14424 19950 14476
rect 20070 14464 20076 14476
rect 20031 14436 20076 14464
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 20990 14424 20996 14476
rect 21048 14464 21054 14476
rect 21453 14467 21511 14473
rect 21453 14464 21465 14467
rect 21048 14436 21465 14464
rect 21048 14424 21054 14436
rect 21453 14433 21465 14436
rect 21499 14433 21511 14467
rect 21453 14427 21511 14433
rect 23216 14464 23244 14504
rect 23750 14464 23756 14476
rect 23216 14436 23756 14464
rect 18046 14396 18052 14408
rect 17696 14368 18052 14396
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 19334 14396 19340 14408
rect 18279 14368 19340 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19426 14356 19432 14408
rect 19484 14356 19490 14408
rect 20714 14396 20720 14408
rect 20675 14368 20720 14396
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 21634 14396 21640 14408
rect 21595 14368 21640 14396
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 22554 14396 22560 14408
rect 22515 14368 22560 14396
rect 22554 14356 22560 14368
rect 22612 14356 22618 14408
rect 23216 14405 23244 14436
rect 23750 14424 23756 14436
rect 23808 14424 23814 14476
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14365 23259 14399
rect 23201 14359 23259 14365
rect 23474 14356 23480 14408
rect 23532 14396 23538 14408
rect 28353 14399 28411 14405
rect 28353 14396 28365 14399
rect 23532 14368 28365 14396
rect 23532 14356 23538 14368
rect 28353 14365 28365 14368
rect 28399 14365 28411 14399
rect 28353 14359 28411 14365
rect 13814 14328 13820 14340
rect 13096 14300 13820 14328
rect 1762 14260 1768 14272
rect 1723 14232 1768 14260
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 3237 14263 3295 14269
rect 3237 14229 3249 14263
rect 3283 14260 3295 14263
rect 4062 14260 4068 14272
rect 3283 14232 4068 14260
rect 3283 14229 3295 14232
rect 3237 14223 3295 14229
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 6546 14220 6552 14272
rect 6604 14260 6610 14272
rect 6641 14263 6699 14269
rect 6641 14260 6653 14263
rect 6604 14232 6653 14260
rect 6604 14220 6610 14232
rect 6641 14229 6653 14232
rect 6687 14229 6699 14263
rect 7374 14260 7380 14272
rect 7335 14232 7380 14260
rect 6641 14223 6699 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 9692 14269 9720 14300
rect 13814 14288 13820 14300
rect 13872 14328 13878 14340
rect 13998 14328 14004 14340
rect 13872 14300 14004 14328
rect 13872 14288 13878 14300
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 16302 14331 16360 14337
rect 16302 14297 16314 14331
rect 16348 14297 16360 14331
rect 16302 14291 16360 14297
rect 16393 14331 16451 14337
rect 16393 14297 16405 14331
rect 16439 14328 16451 14331
rect 16574 14328 16580 14340
rect 16439 14300 16580 14328
rect 16439 14297 16451 14300
rect 16393 14291 16451 14297
rect 9677 14263 9735 14269
rect 9677 14229 9689 14263
rect 9723 14229 9735 14263
rect 13630 14260 13636 14272
rect 13591 14232 13636 14260
rect 9677 14223 9735 14229
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 14277 14263 14335 14269
rect 14277 14229 14289 14263
rect 14323 14260 14335 14263
rect 15010 14260 15016 14272
rect 14323 14232 15016 14260
rect 14323 14229 14335 14232
rect 14277 14223 14335 14229
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 16317 14260 16345 14291
rect 16574 14288 16580 14300
rect 16632 14288 16638 14340
rect 18598 14328 18604 14340
rect 17696 14300 18604 14328
rect 17696 14260 17724 14300
rect 18598 14288 18604 14300
rect 18656 14288 18662 14340
rect 19444 14328 19472 14356
rect 19352 14300 19472 14328
rect 19705 14331 19763 14337
rect 19352 14272 19380 14300
rect 19705 14297 19717 14331
rect 19751 14297 19763 14331
rect 19705 14291 19763 14297
rect 16317 14232 17724 14260
rect 17770 14220 17776 14272
rect 17828 14260 17834 14272
rect 18877 14263 18935 14269
rect 18877 14260 18889 14263
rect 17828 14232 18889 14260
rect 17828 14220 17834 14232
rect 18877 14229 18889 14232
rect 18923 14229 18935 14263
rect 18877 14223 18935 14229
rect 19334 14220 19340 14272
rect 19392 14220 19398 14272
rect 19426 14220 19432 14272
rect 19484 14260 19490 14272
rect 19720 14260 19748 14291
rect 19484 14232 19748 14260
rect 22097 14263 22155 14269
rect 19484 14220 19490 14232
rect 22097 14229 22109 14263
rect 22143 14260 22155 14263
rect 22370 14260 22376 14272
rect 22143 14232 22376 14260
rect 22143 14229 22155 14232
rect 22097 14223 22155 14229
rect 22370 14220 22376 14232
rect 22428 14220 22434 14272
rect 22462 14220 22468 14272
rect 22520 14260 22526 14272
rect 23293 14263 23351 14269
rect 23293 14260 23305 14263
rect 22520 14232 23305 14260
rect 22520 14220 22526 14232
rect 23293 14229 23305 14232
rect 23339 14229 23351 14263
rect 23293 14223 23351 14229
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 1728 14028 4997 14056
rect 1728 14016 1734 14028
rect 4985 14025 4997 14028
rect 5031 14025 5043 14059
rect 4985 14019 5043 14025
rect 5994 14016 6000 14068
rect 6052 14056 6058 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6052 14028 6837 14056
rect 6052 14016 6058 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 6825 14019 6883 14025
rect 7926 14016 7932 14068
rect 7984 14056 7990 14068
rect 8113 14059 8171 14065
rect 8113 14056 8125 14059
rect 7984 14028 8125 14056
rect 7984 14016 7990 14028
rect 8113 14025 8125 14028
rect 8159 14025 8171 14059
rect 8113 14019 8171 14025
rect 9125 14059 9183 14065
rect 9125 14025 9137 14059
rect 9171 14056 9183 14059
rect 9398 14056 9404 14068
rect 9171 14028 9404 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 10594 14056 10600 14068
rect 9815 14028 10600 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 13630 14016 13636 14068
rect 13688 14056 13694 14068
rect 13688 14028 17080 14056
rect 13688 14016 13694 14028
rect 1857 13991 1915 13997
rect 1857 13957 1869 13991
rect 1903 13988 1915 13991
rect 2130 13988 2136 14000
rect 1903 13960 2136 13988
rect 1903 13957 1915 13960
rect 1857 13951 1915 13957
rect 2130 13948 2136 13960
rect 2188 13948 2194 14000
rect 2866 13948 2872 14000
rect 2924 13948 2930 14000
rect 7374 13988 7380 14000
rect 5184 13960 7380 13988
rect 4062 13920 4068 13932
rect 4023 13892 4068 13920
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 5184 13929 5212 13960
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 8478 13988 8484 14000
rect 7484 13960 8484 13988
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5408 13892 5825 13920
rect 5408 13880 5414 13892
rect 5813 13889 5825 13892
rect 5859 13920 5871 13923
rect 6178 13920 6184 13932
rect 5859 13892 6184 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 7282 13920 7288 13932
rect 7055 13892 7288 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7282 13880 7288 13892
rect 7340 13920 7346 13932
rect 7484 13920 7512 13960
rect 8478 13948 8484 13960
rect 8536 13948 8542 14000
rect 13814 13988 13820 14000
rect 12406 13960 13820 13988
rect 7340 13892 7512 13920
rect 7653 13923 7711 13929
rect 7340 13880 7346 13892
rect 7653 13889 7665 13923
rect 7699 13920 7711 13923
rect 8570 13920 8576 13932
rect 7699 13892 8576 13920
rect 7699 13889 7711 13892
rect 7653 13883 7711 13889
rect 8570 13880 8576 13892
rect 8628 13920 8634 13932
rect 9033 13923 9091 13929
rect 9033 13920 9045 13923
rect 8628 13892 9045 13920
rect 8628 13880 8634 13892
rect 9033 13889 9045 13892
rect 9079 13889 9091 13923
rect 9033 13883 9091 13889
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 9677 13923 9735 13929
rect 9677 13920 9689 13923
rect 9640 13892 9689 13920
rect 9640 13880 9646 13892
rect 9677 13889 9689 13892
rect 9723 13920 9735 13923
rect 9766 13920 9772 13932
rect 9723 13892 9772 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 10594 13920 10600 13932
rect 10551 13892 10600 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 10962 13920 10968 13932
rect 10923 13892 10968 13920
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 12406 13920 12434 13960
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 14090 13988 14096 14000
rect 14016 13960 14096 13988
rect 12299 13892 12434 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 1946 13812 1952 13864
rect 2004 13852 2010 13864
rect 3881 13855 3939 13861
rect 3881 13852 3893 13855
rect 2004 13824 3893 13852
rect 2004 13812 2010 13824
rect 3881 13821 3893 13824
rect 3927 13821 3939 13855
rect 3881 13815 3939 13821
rect 5905 13855 5963 13861
rect 5905 13821 5917 13855
rect 5951 13852 5963 13855
rect 8018 13852 8024 13864
rect 5951 13824 8024 13852
rect 5951 13821 5963 13824
rect 5905 13815 5963 13821
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 10134 13812 10140 13864
rect 10192 13852 10198 13864
rect 10980 13852 11008 13880
rect 10192 13824 11008 13852
rect 10192 13812 10198 13824
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 12492 13824 12725 13852
rect 12492 13812 12498 13824
rect 12713 13821 12725 13824
rect 12759 13821 12771 13855
rect 12894 13852 12900 13864
rect 12855 13824 12900 13852
rect 12713 13815 12771 13821
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 14016 13861 14044 13960
rect 14090 13948 14096 13960
rect 14148 13948 14154 14000
rect 15010 13948 15016 14000
rect 15068 13988 15074 14000
rect 17052 13997 17080 14028
rect 18230 14016 18236 14068
rect 18288 14056 18294 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 18288 14028 18889 14056
rect 18288 14016 18294 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 19978 14056 19984 14068
rect 19843 14028 19984 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 28810 14056 28816 14068
rect 20088 14028 28816 14056
rect 17037 13991 17095 13997
rect 15068 13960 16252 13988
rect 15068 13948 15074 13960
rect 14826 13880 14832 13932
rect 14884 13920 14890 13932
rect 15657 13923 15715 13929
rect 15657 13920 15669 13923
rect 14884 13892 15669 13920
rect 14884 13880 14890 13892
rect 15657 13889 15669 13892
rect 15703 13889 15715 13923
rect 16224 13918 16252 13960
rect 17037 13957 17049 13991
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 17589 13991 17647 13997
rect 17589 13957 17601 13991
rect 17635 13988 17647 13991
rect 17678 13988 17684 14000
rect 17635 13960 17684 13988
rect 17635 13957 17647 13960
rect 17589 13951 17647 13957
rect 17678 13948 17684 13960
rect 17736 13988 17742 14000
rect 20088 13988 20116 14028
rect 28810 14016 28816 14028
rect 28868 14016 28874 14068
rect 17736 13960 20116 13988
rect 21453 13991 21511 13997
rect 17736 13948 17742 13960
rect 21453 13957 21465 13991
rect 21499 13988 21511 13991
rect 23198 13988 23204 14000
rect 21499 13960 23204 13988
rect 21499 13957 21511 13960
rect 21453 13951 21511 13957
rect 23198 13948 23204 13960
rect 23256 13988 23262 14000
rect 23753 13991 23811 13997
rect 23753 13988 23765 13991
rect 23256 13960 23765 13988
rect 23256 13948 23262 13960
rect 23753 13957 23765 13960
rect 23799 13957 23811 13991
rect 23753 13951 23811 13957
rect 16301 13923 16359 13929
rect 16301 13918 16313 13923
rect 16224 13890 16313 13918
rect 15657 13883 15715 13889
rect 16301 13889 16313 13890
rect 16347 13889 16359 13923
rect 16666 13920 16672 13932
rect 16301 13883 16359 13889
rect 16401 13892 16672 13920
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 14001 13855 14059 13861
rect 13403 13824 13952 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 5500 13756 11192 13784
rect 5500 13744 5506 13756
rect 3142 13676 3148 13728
rect 3200 13716 3206 13728
rect 3329 13719 3387 13725
rect 3329 13716 3341 13719
rect 3200 13688 3341 13716
rect 3200 13676 3206 13688
rect 3329 13685 3341 13688
rect 3375 13685 3387 13719
rect 3329 13679 3387 13685
rect 4525 13719 4583 13725
rect 4525 13685 4537 13719
rect 4571 13716 4583 13719
rect 5074 13716 5080 13728
rect 4571 13688 5080 13716
rect 4571 13685 4583 13688
rect 4525 13679 4583 13685
rect 5074 13676 5080 13688
rect 5132 13676 5138 13728
rect 7469 13719 7527 13725
rect 7469 13685 7481 13719
rect 7515 13716 7527 13719
rect 8202 13716 8208 13728
rect 7515 13688 8208 13716
rect 7515 13685 7527 13688
rect 7469 13679 7527 13685
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 10318 13716 10324 13728
rect 10279 13688 10324 13716
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 11054 13716 11060 13728
rect 11015 13688 11060 13716
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 11164 13716 11192 13756
rect 11422 13744 11428 13796
rect 11480 13784 11486 13796
rect 11698 13784 11704 13796
rect 11480 13756 11704 13784
rect 11480 13744 11486 13756
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 12066 13784 12072 13796
rect 12027 13756 12072 13784
rect 12066 13744 12072 13756
rect 12124 13744 12130 13796
rect 13262 13744 13268 13796
rect 13320 13784 13326 13796
rect 13722 13784 13728 13796
rect 13320 13756 13728 13784
rect 13320 13744 13326 13756
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 13924 13784 13952 13824
rect 14001 13821 14013 13855
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 14090 13812 14096 13864
rect 14148 13852 14154 13864
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 14148 13824 14197 13852
rect 14148 13812 14154 13824
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 14185 13815 14243 13821
rect 14645 13855 14703 13861
rect 14645 13821 14657 13855
rect 14691 13852 14703 13855
rect 15378 13852 15384 13864
rect 14691 13824 15384 13852
rect 14691 13821 14703 13824
rect 14645 13815 14703 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 16401 13852 16429 13892
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 18233 13923 18291 13929
rect 18233 13889 18245 13923
rect 18279 13920 18291 13923
rect 19978 13920 19984 13932
rect 18279 13892 19840 13920
rect 19939 13892 19984 13920
rect 18279 13889 18291 13892
rect 18233 13883 18291 13889
rect 15488 13824 16429 13852
rect 15286 13784 15292 13796
rect 13924 13756 15292 13784
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 15488 13793 15516 13824
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16540 13824 16957 13852
rect 16540 13812 16546 13824
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 18414 13852 18420 13864
rect 18375 13824 18420 13852
rect 16945 13815 17003 13821
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 19812 13852 19840 13892
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 20993 13923 21051 13929
rect 20993 13889 21005 13923
rect 21039 13920 21051 13923
rect 22462 13920 22468 13932
rect 21039 13892 22468 13920
rect 21039 13889 21051 13892
rect 20993 13883 21051 13889
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 23109 13923 23167 13929
rect 23109 13889 23121 13923
rect 23155 13920 23167 13923
rect 23155 13892 24348 13920
rect 23155 13889 23167 13892
rect 23109 13883 23167 13889
rect 20438 13852 20444 13864
rect 19812 13824 20444 13852
rect 20438 13812 20444 13824
rect 20496 13852 20502 13864
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 20496 13824 20821 13852
rect 20496 13812 20502 13824
rect 20809 13821 20821 13824
rect 20855 13852 20867 13855
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 20855 13824 22017 13852
rect 20855 13821 20867 13824
rect 20809 13815 20867 13821
rect 22005 13821 22017 13824
rect 22051 13821 22063 13855
rect 22186 13852 22192 13864
rect 22147 13824 22192 13852
rect 22005 13815 22063 13821
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 23293 13855 23351 13861
rect 23293 13821 23305 13855
rect 23339 13852 23351 13855
rect 24320 13852 24348 13892
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 24452 13892 24497 13920
rect 24452 13880 24458 13892
rect 34238 13880 34244 13932
rect 34296 13920 34302 13932
rect 38013 13923 38071 13929
rect 38013 13920 38025 13923
rect 34296 13892 38025 13920
rect 34296 13880 34302 13892
rect 38013 13889 38025 13892
rect 38059 13889 38071 13923
rect 38013 13883 38071 13889
rect 34698 13852 34704 13864
rect 23339 13824 24256 13852
rect 24320 13824 34704 13852
rect 23339 13821 23351 13824
rect 23293 13815 23351 13821
rect 15473 13787 15531 13793
rect 15473 13753 15485 13787
rect 15519 13753 15531 13787
rect 15473 13747 15531 13753
rect 16117 13787 16175 13793
rect 16117 13753 16129 13787
rect 16163 13784 16175 13787
rect 16390 13784 16396 13796
rect 16163 13756 16396 13784
rect 16163 13753 16175 13756
rect 16117 13747 16175 13753
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 22370 13784 22376 13796
rect 22331 13756 22376 13784
rect 22370 13744 22376 13756
rect 22428 13744 22434 13796
rect 24228 13793 24256 13824
rect 34698 13812 34704 13824
rect 34756 13812 34762 13864
rect 24213 13787 24271 13793
rect 24213 13753 24225 13787
rect 24259 13753 24271 13787
rect 24213 13747 24271 13753
rect 12158 13716 12164 13728
rect 11164 13688 12164 13716
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 14550 13676 14556 13728
rect 14608 13716 14614 13728
rect 16574 13716 16580 13728
rect 14608 13688 16580 13716
rect 14608 13676 14614 13688
rect 16574 13676 16580 13688
rect 16632 13676 16638 13728
rect 38194 13716 38200 13728
rect 38155 13688 38200 13716
rect 38194 13676 38200 13688
rect 38252 13676 38258 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 4341 13515 4399 13521
rect 4341 13481 4353 13515
rect 4387 13512 4399 13515
rect 5810 13512 5816 13524
rect 4387 13484 5816 13512
rect 4387 13481 4399 13484
rect 4341 13475 4399 13481
rect 5810 13472 5816 13484
rect 5868 13472 5874 13524
rect 8021 13515 8079 13521
rect 8021 13481 8033 13515
rect 8067 13512 8079 13515
rect 8110 13512 8116 13524
rect 8067 13484 8116 13512
rect 8067 13481 8079 13484
rect 8021 13475 8079 13481
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 9674 13512 9680 13524
rect 8680 13484 9680 13512
rect 7558 13404 7564 13456
rect 7616 13444 7622 13456
rect 8680 13444 8708 13484
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 10689 13515 10747 13521
rect 10689 13481 10701 13515
rect 10735 13512 10747 13515
rect 12894 13512 12900 13524
rect 10735 13484 12900 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13630 13512 13636 13524
rect 13320 13484 13636 13512
rect 13320 13472 13326 13484
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 14369 13515 14427 13521
rect 14369 13481 14381 13515
rect 14415 13512 14427 13515
rect 14550 13512 14556 13524
rect 14415 13484 14556 13512
rect 14415 13481 14427 13484
rect 14369 13475 14427 13481
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15436 13484 16037 13512
rect 15436 13472 15442 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 16025 13475 16083 13481
rect 17681 13515 17739 13521
rect 17681 13481 17693 13515
rect 17727 13512 17739 13515
rect 17770 13512 17776 13524
rect 17727 13484 17776 13512
rect 17727 13481 17739 13484
rect 17681 13475 17739 13481
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 18598 13512 18604 13524
rect 18559 13484 18604 13512
rect 18598 13472 18604 13484
rect 18656 13472 18662 13524
rect 19978 13472 19984 13524
rect 20036 13512 20042 13524
rect 20625 13515 20683 13521
rect 20625 13512 20637 13515
rect 20036 13484 20637 13512
rect 20036 13472 20042 13484
rect 20625 13481 20637 13484
rect 20671 13481 20683 13515
rect 20625 13475 20683 13481
rect 21634 13472 21640 13524
rect 21692 13512 21698 13524
rect 21821 13515 21879 13521
rect 21821 13512 21833 13515
rect 21692 13484 21833 13512
rect 21692 13472 21698 13484
rect 21821 13481 21833 13484
rect 21867 13481 21879 13515
rect 21821 13475 21879 13481
rect 23569 13515 23627 13521
rect 23569 13481 23581 13515
rect 23615 13512 23627 13515
rect 24394 13512 24400 13524
rect 23615 13484 24400 13512
rect 23615 13481 23627 13484
rect 23569 13475 23627 13481
rect 24394 13472 24400 13484
rect 24452 13472 24458 13524
rect 33410 13512 33416 13524
rect 33371 13484 33416 13512
rect 33410 13472 33416 13484
rect 33468 13472 33474 13524
rect 7616 13416 8708 13444
rect 7616 13404 7622 13416
rect 8754 13404 8760 13456
rect 8812 13444 8818 13456
rect 11146 13444 11152 13456
rect 8812 13416 11152 13444
rect 8812 13404 8818 13416
rect 11146 13404 11152 13416
rect 11204 13404 11210 13456
rect 11241 13447 11299 13453
rect 11241 13413 11253 13447
rect 11287 13444 11299 13447
rect 14458 13444 14464 13456
rect 11287 13416 14464 13444
rect 11287 13413 11299 13416
rect 11241 13407 11299 13413
rect 14458 13404 14464 13416
rect 14516 13404 14522 13456
rect 15654 13404 15660 13456
rect 15712 13444 15718 13456
rect 18230 13444 18236 13456
rect 15712 13416 18236 13444
rect 15712 13404 15718 13416
rect 18230 13404 18236 13416
rect 18288 13404 18294 13456
rect 20070 13444 20076 13456
rect 20031 13416 20076 13444
rect 20070 13404 20076 13416
rect 20128 13404 20134 13456
rect 22370 13404 22376 13456
rect 22428 13404 22434 13456
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 5350 13376 5356 13388
rect 4540 13348 5356 13376
rect 4540 13317 4568 13348
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 6512 13348 6745 13376
rect 6512 13336 6518 13348
rect 6733 13345 6745 13348
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 10870 13376 10876 13388
rect 9272 13348 10876 13376
rect 9272 13336 9278 13348
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11112 13348 12081 13376
rect 11112 13336 11118 13348
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 14918 13376 14924 13388
rect 12492 13348 14924 13376
rect 12492 13336 12498 13348
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 17034 13376 17040 13388
rect 15028 13348 16344 13376
rect 16995 13348 17040 13376
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13277 4583 13311
rect 4982 13308 4988 13320
rect 4943 13280 4988 13308
rect 4525 13271 4583 13277
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 7098 13268 7104 13320
rect 7156 13308 7162 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7156 13280 7389 13308
rect 7156 13268 7162 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 8202 13308 8208 13320
rect 8163 13280 8208 13308
rect 7377 13271 7435 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 9490 13308 9496 13320
rect 9451 13280 9496 13308
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 10468 13280 10609 13308
rect 10468 13268 10474 13280
rect 10597 13277 10609 13280
rect 10643 13277 10655 13311
rect 11422 13308 11428 13320
rect 11383 13280 11428 13308
rect 10597 13271 10655 13277
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 11698 13268 11704 13320
rect 11756 13308 11762 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11756 13280 11897 13308
rect 11756 13268 11762 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 12032 13280 13737 13308
rect 12032 13268 12038 13280
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 1857 13243 1915 13249
rect 1857 13209 1869 13243
rect 1903 13240 1915 13243
rect 1946 13240 1952 13252
rect 1903 13212 1952 13240
rect 1903 13209 1915 13212
rect 1857 13203 1915 13209
rect 1946 13200 1952 13212
rect 2004 13200 2010 13252
rect 3694 13240 3700 13252
rect 3082 13212 3700 13240
rect 3694 13200 3700 13212
rect 3752 13200 3758 13252
rect 5261 13243 5319 13249
rect 5261 13209 5273 13243
rect 5307 13209 5319 13243
rect 7469 13243 7527 13249
rect 5261 13203 5319 13209
rect 5644 13212 5750 13240
rect 3329 13175 3387 13181
rect 3329 13141 3341 13175
rect 3375 13172 3387 13175
rect 4430 13172 4436 13184
rect 3375 13144 4436 13172
rect 3375 13141 3387 13144
rect 3329 13135 3387 13141
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 5276 13172 5304 13203
rect 5644 13184 5672 13212
rect 7469 13209 7481 13243
rect 7515 13240 7527 13243
rect 10226 13240 10232 13252
rect 7515 13212 10232 13240
rect 7515 13209 7527 13212
rect 7469 13203 7527 13209
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 14568 13240 14596 13271
rect 15028 13240 15056 13348
rect 15102 13268 15108 13320
rect 15160 13308 15166 13320
rect 15197 13311 15255 13317
rect 15197 13308 15209 13311
rect 15160 13280 15209 13308
rect 15160 13268 15166 13280
rect 15197 13277 15209 13280
rect 15243 13277 15255 13311
rect 15654 13308 15660 13320
rect 15615 13280 15660 13308
rect 15197 13271 15255 13277
rect 15654 13268 15660 13280
rect 15712 13268 15718 13320
rect 15838 13308 15844 13320
rect 15799 13280 15844 13308
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 13556 13212 14596 13240
rect 14660 13212 15056 13240
rect 16316 13240 16344 13348
rect 17034 13336 17040 13348
rect 17092 13336 17098 13388
rect 19521 13379 19579 13385
rect 19521 13345 19533 13379
rect 19567 13376 19579 13379
rect 20346 13376 20352 13388
rect 19567 13348 20352 13376
rect 19567 13345 19579 13348
rect 19521 13339 19579 13345
rect 20346 13336 20352 13348
rect 20404 13376 20410 13388
rect 20622 13376 20628 13388
rect 20404 13348 20628 13376
rect 20404 13336 20410 13348
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 22388 13376 22416 13404
rect 22465 13379 22523 13385
rect 22465 13376 22477 13379
rect 22388 13348 22477 13376
rect 22465 13345 22477 13348
rect 22511 13345 22523 13379
rect 22465 13339 22523 13345
rect 23109 13379 23167 13385
rect 23109 13345 23121 13379
rect 23155 13376 23167 13379
rect 23474 13376 23480 13388
rect 23155 13348 23480 13376
rect 23155 13345 23167 13348
rect 23109 13339 23167 13345
rect 23474 13336 23480 13348
rect 23532 13376 23538 13388
rect 24026 13376 24032 13388
rect 23532 13348 24032 13376
rect 23532 13336 23538 13348
rect 24026 13336 24032 13348
rect 24084 13336 24090 13388
rect 17218 13308 17224 13320
rect 17179 13280 17224 13308
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 18230 13308 18236 13320
rect 18191 13280 18236 13308
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 18417 13311 18475 13317
rect 18417 13308 18429 13311
rect 18380 13280 18429 13308
rect 18380 13268 18386 13280
rect 18417 13277 18429 13280
rect 18463 13277 18475 13311
rect 18417 13271 18475 13277
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 20772 13280 20821 13308
rect 20772 13268 20778 13280
rect 20809 13277 20821 13280
rect 20855 13277 20867 13311
rect 21726 13308 21732 13320
rect 21687 13280 21732 13308
rect 20809 13271 20867 13277
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 23750 13308 23756 13320
rect 23711 13280 23756 13308
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 33321 13311 33379 13317
rect 33321 13277 33333 13311
rect 33367 13308 33379 13311
rect 34606 13308 34612 13320
rect 33367 13280 34612 13308
rect 33367 13277 33379 13280
rect 33321 13271 33379 13277
rect 34606 13268 34612 13280
rect 34664 13268 34670 13320
rect 19613 13243 19671 13249
rect 16316 13212 17908 13240
rect 5350 13172 5356 13184
rect 5276 13144 5356 13172
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 5626 13132 5632 13184
rect 5684 13132 5690 13184
rect 9306 13172 9312 13184
rect 9267 13144 9312 13172
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 9953 13175 10011 13181
rect 9953 13141 9965 13175
rect 9999 13172 10011 13175
rect 10502 13172 10508 13184
rect 9999 13144 10508 13172
rect 9999 13141 10011 13144
rect 9953 13135 10011 13141
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 11054 13172 11060 13184
rect 10744 13144 11060 13172
rect 10744 13132 10750 13144
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11330 13172 11336 13184
rect 11204 13144 11336 13172
rect 11204 13132 11210 13144
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 11514 13132 11520 13184
rect 11572 13172 11578 13184
rect 11974 13172 11980 13184
rect 11572 13144 11980 13172
rect 11572 13132 11578 13144
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 12158 13132 12164 13184
rect 12216 13172 12222 13184
rect 12434 13172 12440 13184
rect 12216 13144 12440 13172
rect 12216 13132 12222 13144
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12618 13172 12624 13184
rect 12575 13144 12624 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 13556 13181 13584 13212
rect 13541 13175 13599 13181
rect 13541 13141 13553 13175
rect 13587 13141 13599 13175
rect 13541 13135 13599 13141
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 14660 13172 14688 13212
rect 13688 13144 14688 13172
rect 15013 13175 15071 13181
rect 13688 13132 13694 13144
rect 15013 13141 15025 13175
rect 15059 13172 15071 13175
rect 17770 13172 17776 13184
rect 15059 13144 17776 13172
rect 15059 13141 15071 13144
rect 15013 13135 15071 13141
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 17880 13172 17908 13212
rect 19613 13209 19625 13243
rect 19659 13240 19671 13243
rect 19978 13240 19984 13252
rect 19659 13212 19984 13240
rect 19659 13209 19671 13212
rect 19613 13203 19671 13209
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 22554 13200 22560 13252
rect 22612 13240 22618 13252
rect 22612 13212 22657 13240
rect 22612 13200 22618 13212
rect 21634 13172 21640 13184
rect 17880 13144 21640 13172
rect 21634 13132 21640 13144
rect 21692 13132 21698 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 3421 12971 3479 12977
rect 3421 12937 3433 12971
rect 3467 12937 3479 12971
rect 3421 12931 3479 12937
rect 3326 12900 3332 12912
rect 3174 12872 3332 12900
rect 3326 12860 3332 12872
rect 3384 12860 3390 12912
rect 3436 12900 3464 12931
rect 3878 12928 3884 12980
rect 3936 12968 3942 12980
rect 4982 12968 4988 12980
rect 3936 12940 4988 12968
rect 3936 12928 3942 12940
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 5074 12928 5080 12980
rect 5132 12968 5138 12980
rect 8938 12968 8944 12980
rect 5132 12940 5488 12968
rect 5132 12928 5138 12940
rect 4154 12900 4160 12912
rect 3436 12872 4160 12900
rect 4154 12860 4160 12872
rect 4212 12860 4218 12912
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 1673 12835 1731 12841
rect 1673 12832 1685 12835
rect 1636 12804 1685 12832
rect 1636 12792 1642 12804
rect 1673 12801 1685 12804
rect 1719 12801 1731 12835
rect 3878 12832 3884 12844
rect 3839 12804 3884 12832
rect 1673 12795 1731 12801
rect 3878 12792 3884 12804
rect 3936 12792 3942 12844
rect 5258 12792 5264 12844
rect 5316 12792 5322 12844
rect 5460 12832 5488 12940
rect 7944 12940 8944 12968
rect 5718 12860 5724 12912
rect 5776 12900 5782 12912
rect 7098 12900 7104 12912
rect 5776 12872 7104 12900
rect 5776 12860 5782 12872
rect 7098 12860 7104 12872
rect 7156 12900 7162 12912
rect 7466 12900 7472 12912
rect 7156 12872 7472 12900
rect 7156 12860 7162 12872
rect 7466 12860 7472 12872
rect 7524 12860 7530 12912
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 5460 12804 6561 12832
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 7944 12832 7972 12940
rect 8938 12928 8944 12940
rect 8996 12968 9002 12980
rect 9490 12968 9496 12980
rect 8996 12940 9496 12968
rect 8996 12928 9002 12940
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 10965 12971 11023 12977
rect 10965 12937 10977 12971
rect 11011 12968 11023 12971
rect 11793 12971 11851 12977
rect 11011 12940 11468 12968
rect 11011 12937 11023 12940
rect 10965 12931 11023 12937
rect 8113 12903 8171 12909
rect 8113 12869 8125 12903
rect 8159 12900 8171 12903
rect 11330 12900 11336 12912
rect 8159 12872 11336 12900
rect 8159 12869 8171 12872
rect 8113 12863 8171 12869
rect 11330 12860 11336 12872
rect 11388 12860 11394 12912
rect 11440 12900 11468 12940
rect 11793 12937 11805 12971
rect 11839 12968 11851 12971
rect 15013 12971 15071 12977
rect 11839 12940 14504 12968
rect 11839 12937 11851 12940
rect 11793 12931 11851 12937
rect 11440 12872 12020 12900
rect 6549 12795 6607 12801
rect 6656 12804 7972 12832
rect 8021 12835 8079 12841
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 3418 12764 3424 12776
rect 1995 12736 3424 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 3418 12724 3424 12736
rect 3476 12764 3482 12776
rect 4522 12764 4528 12776
rect 3476 12736 4528 12764
rect 3476 12724 3482 12736
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 4706 12724 4712 12776
rect 4764 12764 4770 12776
rect 5166 12764 5172 12776
rect 4764 12736 5172 12764
rect 4764 12724 4770 12736
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 6656 12764 6684 12804
rect 8021 12801 8033 12835
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 5408 12736 6684 12764
rect 6733 12767 6791 12773
rect 5408 12724 5414 12736
rect 6733 12733 6745 12767
rect 6779 12733 6791 12767
rect 6733 12727 6791 12733
rect 3344 12668 3556 12696
rect 1670 12588 1676 12640
rect 1728 12628 1734 12640
rect 3344 12628 3372 12668
rect 1728 12600 3372 12628
rect 3528 12628 3556 12668
rect 3694 12656 3700 12708
rect 3752 12696 3758 12708
rect 3878 12696 3884 12708
rect 3752 12668 3884 12696
rect 3752 12656 3758 12668
rect 3878 12656 3884 12668
rect 3936 12656 3942 12708
rect 6748 12696 6776 12727
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 7834 12764 7840 12776
rect 7524 12736 7840 12764
rect 7524 12724 7530 12736
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 5184 12668 6776 12696
rect 8036 12696 8064 12795
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8849 12835 8907 12841
rect 8849 12832 8861 12835
rect 8352 12804 8861 12832
rect 8352 12792 8358 12804
rect 8849 12801 8861 12804
rect 8895 12801 8907 12835
rect 10502 12832 10508 12844
rect 10463 12804 10508 12832
rect 8849 12795 8907 12801
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 8665 12767 8723 12773
rect 8665 12733 8677 12767
rect 8711 12764 8723 12767
rect 8754 12764 8760 12776
rect 8711 12736 8760 12764
rect 8711 12733 8723 12736
rect 8665 12727 8723 12733
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 10410 12724 10416 12776
rect 10468 12764 10474 12776
rect 11164 12764 11192 12795
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 11882 12832 11888 12844
rect 11756 12804 11888 12832
rect 11756 12792 11762 12804
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 11992 12841 12020 12872
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 12621 12903 12679 12909
rect 12621 12900 12633 12903
rect 12584 12872 12633 12900
rect 12584 12860 12590 12872
rect 12621 12869 12633 12872
rect 12667 12869 12679 12903
rect 14476 12900 14504 12940
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 15286 12968 15292 12980
rect 15059 12940 15292 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 15930 12928 15936 12980
rect 15988 12968 15994 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 15988 12940 16221 12968
rect 15988 12928 15994 12940
rect 16209 12937 16221 12940
rect 16255 12968 16267 12971
rect 16482 12968 16488 12980
rect 16255 12940 16488 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12968 18199 12971
rect 18414 12968 18420 12980
rect 18187 12940 18420 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 19392 12940 19441 12968
rect 19392 12928 19398 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 19429 12931 19487 12937
rect 19889 12971 19947 12977
rect 19889 12937 19901 12971
rect 19935 12968 19947 12971
rect 20254 12968 20260 12980
rect 19935 12940 20260 12968
rect 19935 12937 19947 12940
rect 19889 12931 19947 12937
rect 20254 12928 20260 12940
rect 20312 12928 20318 12980
rect 21269 12971 21327 12977
rect 21269 12937 21281 12971
rect 21315 12968 21327 12971
rect 22005 12971 22063 12977
rect 21315 12940 21864 12968
rect 21315 12937 21327 12940
rect 21269 12931 21327 12937
rect 17034 12900 17040 12912
rect 14476 12872 14596 12900
rect 12621 12863 12679 12869
rect 14568 12841 14596 12872
rect 16224 12872 17040 12900
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 13909 12835 13967 12841
rect 13909 12801 13921 12835
rect 13955 12832 13967 12835
rect 14553 12835 14611 12841
rect 13955 12804 14504 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 10468 12736 11192 12764
rect 12529 12767 12587 12773
rect 10468 12724 10474 12736
rect 12529 12733 12541 12767
rect 12575 12764 12587 12767
rect 12802 12764 12808 12776
rect 12575 12736 12808 12764
rect 12575 12733 12587 12736
rect 12529 12727 12587 12733
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12764 13231 12767
rect 13262 12764 13268 12776
rect 13219 12736 13268 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14274 12764 14280 12776
rect 14148 12736 14280 12764
rect 14148 12724 14154 12736
rect 14274 12724 14280 12736
rect 14332 12764 14338 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14332 12736 14381 12764
rect 14332 12724 14338 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14476 12764 14504 12804
rect 14553 12801 14565 12835
rect 14599 12801 14611 12835
rect 15746 12832 15752 12844
rect 15707 12804 15752 12832
rect 14553 12795 14611 12801
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 15102 12764 15108 12776
rect 14476 12736 15108 12764
rect 14369 12727 14427 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12764 15623 12767
rect 16114 12764 16120 12776
rect 15611 12736 16120 12764
rect 15611 12733 15623 12736
rect 15565 12727 15623 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 8036 12668 10824 12696
rect 5184 12628 5212 12668
rect 3528 12600 5212 12628
rect 5629 12631 5687 12637
rect 1728 12588 1734 12600
rect 5629 12597 5641 12631
rect 5675 12628 5687 12631
rect 5718 12628 5724 12640
rect 5675 12600 5724 12628
rect 5675 12597 5687 12600
rect 5629 12591 5687 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 6917 12631 6975 12637
rect 6917 12628 6929 12631
rect 6880 12600 6929 12628
rect 6880 12588 6886 12600
rect 6917 12597 6929 12600
rect 6963 12597 6975 12631
rect 6917 12591 6975 12597
rect 9309 12631 9367 12637
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9582 12628 9588 12640
rect 9355 12600 9588 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 10321 12631 10379 12637
rect 10321 12597 10333 12631
rect 10367 12628 10379 12631
rect 10686 12628 10692 12640
rect 10367 12600 10692 12628
rect 10367 12597 10379 12600
rect 10321 12591 10379 12597
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 10796 12628 10824 12668
rect 10870 12656 10876 12708
rect 10928 12696 10934 12708
rect 13630 12696 13636 12708
rect 10928 12668 13636 12696
rect 10928 12656 10934 12668
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 13725 12699 13783 12705
rect 13725 12665 13737 12699
rect 13771 12696 13783 12699
rect 16224 12696 16252 12872
rect 17034 12860 17040 12872
rect 17092 12860 17098 12912
rect 17862 12860 17868 12912
rect 17920 12900 17926 12912
rect 20990 12900 20996 12912
rect 17920 12872 20116 12900
rect 17920 12860 17926 12872
rect 18046 12832 18052 12844
rect 18007 12804 18052 12832
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 20088 12841 20116 12872
rect 20180 12872 20996 12900
rect 20073 12835 20131 12841
rect 18156 12804 19472 12832
rect 16666 12724 16672 12776
rect 16724 12764 16730 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 16724 12736 16865 12764
rect 16724 12724 16730 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 17034 12764 17040 12776
rect 16995 12736 17040 12764
rect 16853 12727 16911 12733
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 18156 12696 18184 12804
rect 18782 12764 18788 12776
rect 18743 12736 18788 12764
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 18969 12767 19027 12773
rect 18969 12733 18981 12767
rect 19015 12764 19027 12767
rect 19334 12764 19340 12776
rect 19015 12736 19340 12764
rect 19015 12733 19027 12736
rect 18969 12727 19027 12733
rect 19334 12724 19340 12736
rect 19392 12724 19398 12776
rect 19444 12764 19472 12804
rect 20073 12801 20085 12835
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 20180 12764 20208 12872
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 21726 12900 21732 12912
rect 21468 12872 21732 12900
rect 21468 12841 21496 12872
rect 21726 12860 21732 12872
rect 21784 12860 21790 12912
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12801 20775 12835
rect 20717 12795 20775 12801
rect 21453 12835 21511 12841
rect 21453 12801 21465 12835
rect 21499 12801 21511 12835
rect 21453 12795 21511 12801
rect 19444 12736 20208 12764
rect 13771 12668 16252 12696
rect 16316 12668 18184 12696
rect 13771 12665 13783 12668
rect 13725 12659 13783 12665
rect 16316 12628 16344 12668
rect 18690 12656 18696 12708
rect 18748 12696 18754 12708
rect 20732 12696 20760 12795
rect 21744 12764 21772 12860
rect 21836 12832 21864 12940
rect 22005 12937 22017 12971
rect 22051 12968 22063 12971
rect 22186 12968 22192 12980
rect 22051 12940 22192 12968
rect 22051 12937 22063 12940
rect 22005 12931 22063 12937
rect 22186 12928 22192 12940
rect 22244 12928 22250 12980
rect 22094 12860 22100 12912
rect 22152 12900 22158 12912
rect 23201 12903 23259 12909
rect 23201 12900 23213 12903
rect 22152 12872 23213 12900
rect 22152 12860 22158 12872
rect 23201 12869 23213 12872
rect 23247 12869 23259 12903
rect 23201 12863 23259 12869
rect 23382 12860 23388 12912
rect 23440 12900 23446 12912
rect 23440 12872 24440 12900
rect 23440 12860 23446 12872
rect 24412 12841 24440 12872
rect 22189 12835 22247 12841
rect 21836 12830 22140 12832
rect 22189 12830 22201 12835
rect 21836 12804 22201 12830
rect 22112 12802 22201 12804
rect 22189 12801 22201 12802
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12801 24455 12835
rect 31386 12832 31392 12844
rect 31347 12804 31392 12832
rect 24397 12795 24455 12801
rect 31386 12792 31392 12804
rect 31444 12792 31450 12844
rect 23109 12767 23167 12773
rect 21744 12736 22232 12764
rect 22204 12708 22232 12736
rect 23109 12733 23121 12767
rect 23155 12764 23167 12767
rect 23198 12764 23204 12776
rect 23155 12736 23204 12764
rect 23155 12733 23167 12736
rect 23109 12727 23167 12733
rect 23198 12724 23204 12736
rect 23256 12724 23262 12776
rect 23750 12764 23756 12776
rect 23711 12736 23756 12764
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 18748 12668 20760 12696
rect 18748 12656 18754 12668
rect 22186 12656 22192 12708
rect 22244 12696 22250 12708
rect 23382 12696 23388 12708
rect 22244 12668 23388 12696
rect 22244 12656 22250 12668
rect 23382 12656 23388 12668
rect 23440 12656 23446 12708
rect 31481 12699 31539 12705
rect 31481 12696 31493 12699
rect 23492 12668 31493 12696
rect 10796 12600 16344 12628
rect 16390 12588 16396 12640
rect 16448 12628 16454 12640
rect 17221 12631 17279 12637
rect 17221 12628 17233 12631
rect 16448 12600 17233 12628
rect 16448 12588 16454 12600
rect 17221 12597 17233 12600
rect 17267 12597 17279 12631
rect 17221 12591 17279 12597
rect 19978 12588 19984 12640
rect 20036 12628 20042 12640
rect 20533 12631 20591 12637
rect 20533 12628 20545 12631
rect 20036 12600 20545 12628
rect 20036 12588 20042 12600
rect 20533 12597 20545 12600
rect 20579 12597 20591 12631
rect 20533 12591 20591 12597
rect 20622 12588 20628 12640
rect 20680 12628 20686 12640
rect 22278 12628 22284 12640
rect 20680 12600 22284 12628
rect 20680 12588 20686 12600
rect 22278 12588 22284 12600
rect 22336 12628 22342 12640
rect 23492 12628 23520 12668
rect 31481 12665 31493 12668
rect 31527 12665 31539 12699
rect 31481 12659 31539 12665
rect 22336 12600 23520 12628
rect 22336 12588 22342 12600
rect 23566 12588 23572 12640
rect 23624 12628 23630 12640
rect 24213 12631 24271 12637
rect 24213 12628 24225 12631
rect 23624 12600 24225 12628
rect 23624 12588 23630 12600
rect 24213 12597 24225 12600
rect 24259 12597 24271 12631
rect 24213 12591 24271 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 6822 12424 6828 12436
rect 5868 12396 6828 12424
rect 5868 12384 5874 12396
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 9861 12427 9919 12433
rect 6932 12396 8248 12424
rect 4338 12316 4344 12368
rect 4396 12356 4402 12368
rect 5258 12356 5264 12368
rect 4396 12328 5264 12356
rect 4396 12316 4402 12328
rect 5258 12316 5264 12328
rect 5316 12356 5322 12368
rect 5316 12328 5580 12356
rect 5316 12316 5322 12328
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12288 4583 12291
rect 4798 12288 4804 12300
rect 4571 12260 4804 12288
rect 4571 12257 4583 12260
rect 4525 12251 4583 12257
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 4982 12248 4988 12300
rect 5040 12288 5046 12300
rect 5445 12291 5503 12297
rect 5445 12288 5457 12291
rect 5040 12260 5457 12288
rect 5040 12248 5046 12260
rect 5445 12257 5457 12260
rect 5491 12257 5503 12291
rect 5552 12288 5580 12328
rect 6932 12288 6960 12396
rect 7190 12316 7196 12368
rect 7248 12356 7254 12368
rect 8110 12356 8116 12368
rect 7248 12328 8116 12356
rect 7248 12316 7254 12328
rect 8110 12316 8116 12328
rect 8168 12316 8174 12368
rect 8220 12356 8248 12396
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 9950 12424 9956 12436
rect 9907 12396 9956 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 10781 12427 10839 12433
rect 10781 12393 10793 12427
rect 10827 12424 10839 12427
rect 12434 12424 12440 12436
rect 10827 12396 12440 12424
rect 10827 12393 10839 12396
rect 10781 12387 10839 12393
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 14918 12384 14924 12436
rect 14976 12424 14982 12436
rect 17681 12427 17739 12433
rect 14976 12396 17632 12424
rect 14976 12384 14982 12396
rect 8220 12328 11100 12356
rect 5552 12260 6960 12288
rect 7837 12291 7895 12297
rect 5445 12251 5503 12257
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 8018 12288 8024 12300
rect 7883 12260 8024 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 9490 12288 9496 12300
rect 9263 12260 9496 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10410 12288 10416 12300
rect 9916 12260 10416 12288
rect 9916 12248 9922 12260
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 1670 12220 1676 12232
rect 1631 12192 1676 12220
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 4154 12220 4160 12232
rect 3844 12192 4160 12220
rect 3844 12180 3850 12192
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12220 4399 12223
rect 5166 12220 5172 12232
rect 4387 12192 5172 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 7653 12223 7711 12229
rect 7653 12189 7665 12223
rect 7699 12189 7711 12223
rect 7653 12183 7711 12189
rect 1949 12155 2007 12161
rect 1949 12121 1961 12155
rect 1995 12121 2007 12155
rect 4062 12152 4068 12164
rect 3174 12124 4068 12152
rect 1949 12115 2007 12121
rect 1964 12084 1992 12115
rect 4062 12112 4068 12124
rect 4120 12112 4126 12164
rect 4890 12112 4896 12164
rect 4948 12152 4954 12164
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 4948 12124 4997 12152
rect 4948 12112 4954 12124
rect 4985 12121 4997 12124
rect 5031 12121 5043 12155
rect 5718 12152 5724 12164
rect 5679 12124 5724 12152
rect 4985 12115 5043 12121
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 5828 12124 6210 12152
rect 2958 12084 2964 12096
rect 1964 12056 2964 12084
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 3234 12044 3240 12096
rect 3292 12084 3298 12096
rect 3421 12087 3479 12093
rect 3421 12084 3433 12087
rect 3292 12056 3433 12084
rect 3292 12044 3298 12056
rect 3421 12053 3433 12056
rect 3467 12053 3479 12087
rect 3421 12047 3479 12053
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 5828 12084 5856 12124
rect 7006 12112 7012 12164
rect 7064 12152 7070 12164
rect 7668 12152 7696 12183
rect 8294 12180 8300 12232
rect 8352 12220 8358 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 8352 12192 9413 12220
rect 8352 12180 8358 12192
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 10318 12180 10324 12232
rect 10376 12220 10382 12232
rect 10965 12223 11023 12229
rect 10965 12220 10977 12223
rect 10376 12192 10977 12220
rect 10376 12180 10382 12192
rect 10965 12189 10977 12192
rect 11011 12189 11023 12223
rect 11072 12220 11100 12328
rect 11606 12316 11612 12368
rect 11664 12356 11670 12368
rect 11793 12359 11851 12365
rect 11793 12356 11805 12359
rect 11664 12328 11805 12356
rect 11664 12316 11670 12328
rect 11793 12325 11805 12328
rect 11839 12356 11851 12359
rect 16666 12356 16672 12368
rect 11839 12328 14320 12356
rect 11839 12325 11851 12328
rect 11793 12319 11851 12325
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12288 11483 12291
rect 11882 12288 11888 12300
rect 11471 12260 11888 12288
rect 11471 12257 11483 12260
rect 11425 12251 11483 12257
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 12618 12288 12624 12300
rect 12579 12260 12624 12288
rect 12618 12248 12624 12260
rect 12676 12248 12682 12300
rect 12802 12248 12808 12300
rect 12860 12288 12866 12300
rect 12986 12288 12992 12300
rect 12860 12260 12992 12288
rect 12860 12248 12866 12260
rect 12986 12248 12992 12260
rect 13044 12248 13050 12300
rect 11514 12220 11520 12232
rect 11072 12192 11520 12220
rect 10965 12183 11023 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12220 11667 12223
rect 12434 12220 12440 12232
rect 11655 12192 12440 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 12406 12186 12440 12192
rect 12434 12180 12440 12186
rect 12492 12180 12498 12232
rect 14292 12220 14320 12328
rect 14476 12328 16672 12356
rect 14476 12297 14504 12328
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 17604 12356 17632 12396
rect 17681 12393 17693 12427
rect 17727 12424 17739 12427
rect 18322 12424 18328 12436
rect 17727 12396 18328 12424
rect 17727 12393 17739 12396
rect 17681 12387 17739 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19613 12427 19671 12433
rect 19613 12424 19625 12427
rect 19484 12396 19625 12424
rect 19484 12384 19490 12396
rect 19613 12393 19625 12396
rect 19659 12393 19671 12427
rect 19613 12387 19671 12393
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 20220 12396 31754 12424
rect 20220 12384 20226 12396
rect 20346 12356 20352 12368
rect 17604 12328 20352 12356
rect 20346 12316 20352 12328
rect 20404 12316 20410 12368
rect 20622 12316 20628 12368
rect 20680 12316 20686 12368
rect 23474 12356 23480 12368
rect 23387 12328 23480 12356
rect 14461 12291 14519 12297
rect 14461 12257 14473 12291
rect 14507 12257 14519 12291
rect 14461 12251 14519 12257
rect 15105 12291 15163 12297
rect 15105 12257 15117 12291
rect 15151 12288 15163 12291
rect 16298 12288 16304 12300
rect 15151 12260 16304 12288
rect 15151 12257 15163 12260
rect 15105 12251 15163 12257
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 16574 12288 16580 12300
rect 16535 12260 16580 12288
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 18230 12248 18236 12300
rect 18288 12288 18294 12300
rect 18325 12291 18383 12297
rect 18325 12288 18337 12291
rect 18288 12260 18337 12288
rect 18288 12248 18294 12260
rect 18325 12257 18337 12260
rect 18371 12257 18383 12291
rect 18325 12251 18383 12257
rect 20441 12291 20499 12297
rect 20441 12257 20453 12291
rect 20487 12288 20499 12291
rect 20640 12288 20668 12316
rect 23400 12297 23428 12328
rect 23474 12316 23480 12328
rect 23532 12356 23538 12368
rect 24949 12359 25007 12365
rect 24949 12356 24961 12359
rect 23532 12328 24961 12356
rect 23532 12316 23538 12328
rect 24949 12325 24961 12328
rect 24995 12325 25007 12359
rect 24949 12319 25007 12325
rect 20487 12260 20668 12288
rect 23385 12291 23443 12297
rect 20487 12257 20499 12260
rect 20441 12251 20499 12257
rect 23385 12257 23397 12291
rect 23431 12257 23443 12291
rect 24026 12288 24032 12300
rect 23987 12260 24032 12288
rect 23385 12251 23443 12257
rect 24026 12248 24032 12260
rect 24084 12248 24090 12300
rect 14642 12220 14648 12232
rect 14292 12192 14648 12220
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 16114 12220 16120 12232
rect 15335 12192 16120 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12220 17923 12223
rect 18414 12220 18420 12232
rect 17911 12192 18420 12220
rect 17911 12189 17923 12192
rect 17865 12183 17923 12189
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12220 19855 12223
rect 19978 12220 19984 12232
rect 19843 12192 19984 12220
rect 19843 12189 19855 12192
rect 19797 12183 19855 12189
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 20625 12223 20683 12229
rect 20625 12189 20637 12223
rect 20671 12189 20683 12223
rect 21542 12220 21548 12232
rect 21503 12192 21548 12220
rect 20625 12183 20683 12189
rect 9582 12152 9588 12164
rect 7064 12124 7328 12152
rect 7668 12124 9588 12152
rect 7064 12112 7070 12124
rect 7300 12096 7328 12124
rect 9582 12112 9588 12124
rect 9640 12112 9646 12164
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 9732 12124 10088 12152
rect 9732 12112 9738 12124
rect 7190 12084 7196 12096
rect 3568 12056 5856 12084
rect 7151 12056 7196 12084
rect 3568 12044 3574 12056
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7282 12044 7288 12096
rect 7340 12084 7346 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 7340 12056 8309 12084
rect 7340 12044 7346 12056
rect 8297 12053 8309 12056
rect 8343 12053 8355 12087
rect 10060 12084 10088 12124
rect 12250 12112 12256 12164
rect 12308 12152 12314 12164
rect 12713 12155 12771 12161
rect 12308 12124 12572 12152
rect 12308 12112 12314 12124
rect 12434 12084 12440 12096
rect 10060 12056 12440 12084
rect 8297 12047 8355 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12544 12084 12572 12124
rect 12713 12121 12725 12155
rect 12759 12121 12771 12155
rect 13262 12152 13268 12164
rect 13175 12124 13268 12152
rect 12713 12115 12771 12121
rect 12728 12084 12756 12115
rect 13262 12112 13268 12124
rect 13320 12152 13326 12164
rect 13446 12152 13452 12164
rect 13320 12124 13452 12152
rect 13320 12112 13326 12124
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 16393 12155 16451 12161
rect 16393 12152 16405 12155
rect 15252 12124 16405 12152
rect 15252 12112 15258 12124
rect 16393 12121 16405 12124
rect 16439 12121 16451 12155
rect 16393 12115 16451 12121
rect 16574 12112 16580 12164
rect 16632 12152 16638 12164
rect 18506 12152 18512 12164
rect 16632 12124 18512 12152
rect 16632 12112 16638 12124
rect 18506 12112 18512 12124
rect 18564 12112 18570 12164
rect 20640 12152 20668 12183
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 21726 12180 21732 12232
rect 21784 12220 21790 12232
rect 22373 12223 22431 12229
rect 22373 12220 22385 12223
rect 21784 12192 22385 12220
rect 21784 12180 21790 12192
rect 22373 12189 22385 12192
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 24118 12180 24124 12232
rect 24176 12220 24182 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 24176 12192 24593 12220
rect 24176 12180 24182 12192
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 31726 12220 31754 12396
rect 35437 12223 35495 12229
rect 35437 12220 35449 12223
rect 31726 12192 35449 12220
rect 24765 12183 24823 12189
rect 35437 12189 35449 12192
rect 35483 12189 35495 12223
rect 35437 12183 35495 12189
rect 21637 12155 21695 12161
rect 21637 12152 21649 12155
rect 20640 12124 21649 12152
rect 21637 12121 21649 12124
rect 21683 12121 21695 12155
rect 21637 12115 21695 12121
rect 23477 12155 23535 12161
rect 23477 12121 23489 12155
rect 23523 12152 23535 12155
rect 24670 12152 24676 12164
rect 23523 12124 24676 12152
rect 23523 12121 23535 12124
rect 23477 12115 23535 12121
rect 24670 12112 24676 12124
rect 24728 12112 24734 12164
rect 12544 12056 12756 12084
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 14734 12084 14740 12096
rect 14056 12056 14740 12084
rect 14056 12044 14062 12056
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15562 12044 15568 12096
rect 15620 12084 15626 12096
rect 15749 12087 15807 12093
rect 15749 12084 15761 12087
rect 15620 12056 15761 12084
rect 15620 12044 15626 12056
rect 15749 12053 15761 12056
rect 15795 12084 15807 12087
rect 16298 12084 16304 12096
rect 15795 12056 16304 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 20438 12044 20444 12096
rect 20496 12084 20502 12096
rect 21085 12087 21143 12093
rect 21085 12084 21097 12087
rect 20496 12056 21097 12084
rect 20496 12044 20502 12056
rect 21085 12053 21097 12056
rect 21131 12053 21143 12087
rect 21085 12047 21143 12053
rect 21174 12044 21180 12096
rect 21232 12084 21238 12096
rect 22189 12087 22247 12093
rect 22189 12084 22201 12087
rect 21232 12056 22201 12084
rect 21232 12044 21238 12056
rect 22189 12053 22201 12056
rect 22235 12053 22247 12087
rect 22189 12047 22247 12053
rect 23842 12044 23848 12096
rect 23900 12084 23906 12096
rect 24780 12084 24808 12183
rect 23900 12056 24808 12084
rect 35529 12087 35587 12093
rect 23900 12044 23906 12056
rect 35529 12053 35541 12087
rect 35575 12084 35587 12087
rect 36446 12084 36452 12096
rect 35575 12056 36452 12084
rect 35575 12053 35587 12056
rect 35529 12047 35587 12053
rect 36446 12044 36452 12056
rect 36504 12044 36510 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3016 11852 5028 11880
rect 3016 11840 3022 11852
rect 1857 11815 1915 11821
rect 1857 11781 1869 11815
rect 1903 11812 1915 11815
rect 2038 11812 2044 11824
rect 1903 11784 2044 11812
rect 1903 11781 1915 11784
rect 1857 11775 1915 11781
rect 2038 11772 2044 11784
rect 2096 11772 2102 11824
rect 4062 11812 4068 11824
rect 3818 11784 4068 11812
rect 4062 11772 4068 11784
rect 4120 11772 4126 11824
rect 5000 11812 5028 11852
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 5132 11852 5273 11880
rect 5132 11840 5138 11852
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 5810 11880 5816 11892
rect 5408 11852 5816 11880
rect 5408 11840 5414 11852
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 5951 11852 12204 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6270 11812 6276 11824
rect 5000 11784 6276 11812
rect 6270 11772 6276 11784
rect 6328 11772 6334 11824
rect 6914 11812 6920 11824
rect 6564 11784 6920 11812
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11744 1823 11747
rect 1946 11744 1952 11756
rect 1811 11716 1952 11744
rect 1811 11713 1823 11716
rect 1765 11707 1823 11713
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4304 11716 4629 11744
rect 4304 11704 4310 11716
rect 4617 11713 4629 11716
rect 4663 11744 4675 11747
rect 5074 11744 5080 11756
rect 4663 11716 5080 11744
rect 4663 11713 4675 11716
rect 4617 11707 4675 11713
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 5810 11744 5816 11756
rect 5771 11716 5816 11744
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 6564 11753 6592 11784
rect 6914 11772 6920 11784
rect 6972 11772 6978 11824
rect 7193 11815 7251 11821
rect 7193 11781 7205 11815
rect 7239 11812 7251 11815
rect 7282 11812 7288 11824
rect 7239 11784 7288 11812
rect 7239 11781 7251 11784
rect 7193 11775 7251 11781
rect 7282 11772 7288 11784
rect 7340 11772 7346 11824
rect 11149 11815 11207 11821
rect 11149 11812 11161 11815
rect 7392 11784 9062 11812
rect 9876 11784 11161 11812
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11713 6607 11747
rect 6730 11744 6736 11756
rect 6691 11716 6736 11744
rect 6549 11707 6607 11713
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7392 11744 7420 11784
rect 7064 11716 7420 11744
rect 7653 11747 7711 11753
rect 7064 11704 7070 11716
rect 7653 11713 7665 11747
rect 7699 11744 7711 11747
rect 7926 11744 7932 11756
rect 7699 11716 7932 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 1670 11636 1676 11688
rect 1728 11676 1734 11688
rect 2317 11679 2375 11685
rect 2317 11676 2329 11679
rect 1728 11648 2329 11676
rect 1728 11636 1734 11648
rect 2317 11645 2329 11648
rect 2363 11645 2375 11679
rect 2317 11639 2375 11645
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 3050 11676 3056 11688
rect 2639 11648 3056 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 3050 11636 3056 11648
rect 3108 11636 3114 11688
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 4065 11679 4123 11685
rect 4065 11676 4077 11679
rect 3660 11648 4077 11676
rect 3660 11636 3666 11648
rect 4065 11645 4077 11648
rect 4111 11645 4123 11679
rect 4798 11676 4804 11688
rect 4759 11648 4804 11676
rect 4065 11639 4123 11645
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 5718 11636 5724 11688
rect 5776 11676 5782 11688
rect 6086 11676 6092 11688
rect 5776 11648 6092 11676
rect 5776 11636 5782 11648
rect 6086 11636 6092 11648
rect 6144 11676 6150 11688
rect 6454 11676 6460 11688
rect 6144 11648 6460 11676
rect 6144 11636 6150 11648
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 8297 11679 8355 11685
rect 8297 11676 8309 11679
rect 6748 11648 8309 11676
rect 6748 11620 6776 11648
rect 8297 11645 8309 11648
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 8662 11676 8668 11688
rect 8619 11648 8668 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 9582 11636 9588 11688
rect 9640 11676 9646 11688
rect 9876 11676 9904 11784
rect 11149 11781 11161 11784
rect 11195 11781 11207 11815
rect 11149 11775 11207 11781
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11744 10563 11747
rect 12066 11744 12072 11756
rect 10551 11716 12072 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12176 11744 12204 11852
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12492 11852 12572 11880
rect 12492 11840 12498 11852
rect 12544 11812 12572 11852
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 12676 11852 12725 11880
rect 12676 11840 12682 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 12713 11843 12771 11849
rect 13170 11840 13176 11892
rect 13228 11840 13234 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 14240 11852 14289 11880
rect 14240 11840 14246 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 14921 11883 14979 11889
rect 14921 11849 14933 11883
rect 14967 11849 14979 11883
rect 14921 11843 14979 11849
rect 13188 11812 13216 11840
rect 12544 11784 13216 11812
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 14936 11812 14964 11843
rect 15010 11840 15016 11892
rect 15068 11880 15074 11892
rect 16574 11880 16580 11892
rect 15068 11852 16580 11880
rect 15068 11840 15074 11852
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 17037 11883 17095 11889
rect 17037 11849 17049 11883
rect 17083 11880 17095 11883
rect 17218 11880 17224 11892
rect 17083 11852 17224 11880
rect 17083 11849 17095 11852
rect 17037 11843 17095 11849
rect 17218 11840 17224 11852
rect 17276 11840 17282 11892
rect 17589 11883 17647 11889
rect 17589 11849 17601 11883
rect 17635 11880 17647 11883
rect 17954 11880 17960 11892
rect 17635 11852 17960 11880
rect 17635 11849 17647 11852
rect 17589 11843 17647 11849
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 18325 11883 18383 11889
rect 18325 11849 18337 11883
rect 18371 11880 18383 11883
rect 20070 11880 20076 11892
rect 18371 11852 20076 11880
rect 18371 11849 18383 11852
rect 18325 11843 18383 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 21085 11883 21143 11889
rect 21085 11849 21097 11883
rect 21131 11880 21143 11883
rect 21726 11880 21732 11892
rect 21131 11852 21732 11880
rect 21131 11849 21143 11852
rect 21085 11843 21143 11849
rect 21726 11840 21732 11852
rect 21784 11840 21790 11892
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 22152 11852 22197 11880
rect 22152 11840 22158 11852
rect 22554 11840 22560 11892
rect 22612 11880 22618 11892
rect 22741 11883 22799 11889
rect 22741 11880 22753 11883
rect 22612 11852 22753 11880
rect 22612 11840 22618 11852
rect 22741 11849 22753 11852
rect 22787 11849 22799 11883
rect 24670 11880 24676 11892
rect 24631 11852 24676 11880
rect 22741 11843 22799 11849
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 34238 11880 34244 11892
rect 34199 11852 34244 11880
rect 34238 11840 34244 11852
rect 34296 11840 34302 11892
rect 34606 11840 34612 11892
rect 34664 11880 34670 11892
rect 38105 11883 38163 11889
rect 38105 11880 38117 11883
rect 34664 11852 38117 11880
rect 34664 11840 34670 11852
rect 38105 11849 38117 11852
rect 38151 11849 38163 11883
rect 38105 11843 38163 11849
rect 21174 11812 21180 11824
rect 13872 11784 14964 11812
rect 19904 11784 21180 11812
rect 13872 11772 13878 11784
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 12176 11716 13185 11744
rect 13173 11713 13185 11716
rect 13219 11713 13231 11747
rect 14458 11744 14464 11756
rect 14419 11716 14464 11744
rect 13173 11707 13231 11713
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 14792 11716 15117 11744
rect 14792 11704 14798 11716
rect 15105 11713 15117 11716
rect 15151 11713 15163 11747
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 15105 11707 15163 11713
rect 15856 11716 16957 11744
rect 9640 11648 9904 11676
rect 9640 11636 9646 11648
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 10284 11648 10701 11676
rect 10284 11636 10290 11648
rect 10689 11645 10701 11648
rect 10735 11645 10747 11679
rect 10689 11639 10747 11645
rect 10778 11636 10784 11688
rect 10836 11676 10842 11688
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 10836 11648 12265 11676
rect 10836 11636 10842 11648
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 13354 11676 13360 11688
rect 13315 11648 13360 11676
rect 12253 11639 12311 11645
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13504 11648 14320 11676
rect 13504 11636 13510 11648
rect 4338 11608 4344 11620
rect 3620 11580 4344 11608
rect 3620 11552 3648 11580
rect 4338 11568 4344 11580
rect 4396 11568 4402 11620
rect 6730 11568 6736 11620
rect 6788 11568 6794 11620
rect 14182 11608 14188 11620
rect 9968 11580 14188 11608
rect 3602 11500 3608 11552
rect 3660 11500 3666 11552
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 7650 11540 7656 11552
rect 5132 11512 7656 11540
rect 5132 11500 5138 11512
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 7745 11543 7803 11549
rect 7745 11509 7757 11543
rect 7791 11540 7803 11543
rect 9968 11540 9996 11580
rect 14182 11568 14188 11580
rect 14240 11568 14246 11620
rect 7791 11512 9996 11540
rect 10045 11543 10103 11549
rect 7791 11509 7803 11512
rect 7745 11503 7803 11509
rect 10045 11509 10057 11543
rect 10091 11540 10103 11543
rect 10318 11540 10324 11552
rect 10091 11512 10324 11540
rect 10091 11509 10103 11512
rect 10045 11503 10103 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 11974 11540 11980 11552
rect 10468 11512 11980 11540
rect 10468 11500 10474 11512
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 13817 11543 13875 11549
rect 13817 11509 13829 11543
rect 13863 11540 13875 11543
rect 14090 11540 14096 11552
rect 13863 11512 14096 11540
rect 13863 11509 13875 11512
rect 13817 11503 13875 11509
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 14292 11540 14320 11648
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 15565 11679 15623 11685
rect 15565 11676 15577 11679
rect 14608 11648 15577 11676
rect 14608 11636 14614 11648
rect 15565 11645 15577 11648
rect 15611 11645 15623 11679
rect 15746 11676 15752 11688
rect 15707 11648 15752 11676
rect 15565 11639 15623 11645
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 14826 11568 14832 11620
rect 14884 11608 14890 11620
rect 15856 11608 15884 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 17770 11744 17776 11756
rect 17731 11716 17776 11744
rect 16945 11707 17003 11713
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 18233 11747 18291 11753
rect 18233 11713 18245 11747
rect 18279 11744 18291 11747
rect 18690 11744 18696 11756
rect 18279 11716 18696 11744
rect 18279 11713 18291 11716
rect 18233 11707 18291 11713
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11744 18935 11747
rect 19426 11744 19432 11756
rect 18923 11716 19432 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 19061 11679 19119 11685
rect 19061 11645 19073 11679
rect 19107 11676 19119 11679
rect 19904 11676 19932 11784
rect 21174 11772 21180 11784
rect 21232 11772 21238 11824
rect 23661 11815 23719 11821
rect 23661 11781 23673 11815
rect 23707 11812 23719 11815
rect 24578 11812 24584 11824
rect 23707 11784 24584 11812
rect 23707 11781 23719 11784
rect 23661 11775 23719 11781
rect 24578 11772 24584 11784
rect 24636 11772 24642 11824
rect 19981 11747 20039 11753
rect 19981 11713 19993 11747
rect 20027 11744 20039 11747
rect 20530 11744 20536 11756
rect 20027 11716 20536 11744
rect 20027 11713 20039 11716
rect 19981 11707 20039 11713
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 20898 11704 20904 11756
rect 20956 11744 20962 11756
rect 21269 11747 21327 11753
rect 21269 11744 21281 11747
rect 20956 11716 21281 11744
rect 20956 11704 20962 11716
rect 21269 11713 21281 11716
rect 21315 11744 21327 11747
rect 21542 11744 21548 11756
rect 21315 11716 21548 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22649 11747 22707 11753
rect 22649 11713 22661 11747
rect 22695 11744 22707 11747
rect 22830 11744 22836 11756
rect 22695 11716 22836 11744
rect 22695 11713 22707 11716
rect 22649 11707 22707 11713
rect 20162 11676 20168 11688
rect 19107 11648 19932 11676
rect 20123 11648 20168 11676
rect 19107 11645 19119 11648
rect 19061 11639 19119 11645
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 20714 11676 20720 11688
rect 20272 11648 20720 11676
rect 14884 11580 15884 11608
rect 16209 11611 16267 11617
rect 14884 11568 14890 11580
rect 16209 11577 16221 11611
rect 16255 11608 16267 11611
rect 20272 11608 20300 11648
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 16255 11580 20300 11608
rect 16255 11577 16267 11580
rect 16209 11571 16267 11577
rect 20346 11568 20352 11620
rect 20404 11608 20410 11620
rect 22020 11608 22048 11707
rect 22830 11704 22836 11716
rect 22888 11704 22894 11756
rect 24210 11704 24216 11756
rect 24268 11744 24274 11756
rect 24857 11747 24915 11753
rect 24857 11744 24869 11747
rect 24268 11716 24869 11744
rect 24268 11704 24274 11716
rect 24857 11713 24869 11716
rect 24903 11713 24915 11747
rect 24857 11707 24915 11713
rect 30374 11704 30380 11756
rect 30432 11744 30438 11756
rect 34425 11747 34483 11753
rect 34425 11744 34437 11747
rect 30432 11716 34437 11744
rect 30432 11704 30438 11716
rect 34425 11713 34437 11716
rect 34471 11713 34483 11747
rect 38286 11744 38292 11756
rect 38247 11716 38292 11744
rect 34425 11707 34483 11713
rect 38286 11704 38292 11716
rect 38344 11704 38350 11756
rect 23569 11679 23627 11685
rect 23569 11645 23581 11679
rect 23615 11676 23627 11679
rect 25317 11679 25375 11685
rect 25317 11676 25329 11679
rect 23615 11648 25329 11676
rect 23615 11645 23627 11648
rect 23569 11639 23627 11645
rect 25317 11645 25329 11648
rect 25363 11645 25375 11679
rect 25317 11639 25375 11645
rect 23658 11608 23664 11620
rect 20404 11580 23664 11608
rect 20404 11568 20410 11580
rect 23658 11568 23664 11580
rect 23716 11568 23722 11620
rect 23750 11568 23756 11620
rect 23808 11608 23814 11620
rect 24121 11611 24179 11617
rect 24121 11608 24133 11611
rect 23808 11580 24133 11608
rect 23808 11568 23814 11580
rect 24121 11577 24133 11580
rect 24167 11608 24179 11611
rect 24302 11608 24308 11620
rect 24167 11580 24308 11608
rect 24167 11577 24179 11580
rect 24121 11571 24179 11577
rect 24302 11568 24308 11580
rect 24360 11568 24366 11620
rect 17586 11540 17592 11552
rect 14292 11512 17592 11540
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 19518 11540 19524 11552
rect 19479 11512 19524 11540
rect 19518 11500 19524 11512
rect 19576 11540 19582 11552
rect 20438 11540 20444 11552
rect 19576 11512 20444 11540
rect 19576 11500 19582 11512
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 20625 11543 20683 11549
rect 20625 11509 20637 11543
rect 20671 11540 20683 11543
rect 20714 11540 20720 11552
rect 20671 11512 20720 11540
rect 20671 11509 20683 11512
rect 20625 11503 20683 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 7190 11336 7196 11348
rect 6932 11308 7196 11336
rect 3421 11271 3479 11277
rect 3421 11237 3433 11271
rect 3467 11268 3479 11271
rect 3602 11268 3608 11280
rect 3467 11240 3608 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 5905 11271 5963 11277
rect 5905 11237 5917 11271
rect 5951 11268 5963 11271
rect 6932 11268 6960 11308
rect 7190 11296 7196 11308
rect 7248 11336 7254 11348
rect 9122 11336 9128 11348
rect 7248 11308 9128 11336
rect 7248 11296 7254 11308
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 13354 11336 13360 11348
rect 9539 11308 13360 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 14274 11336 14280 11348
rect 13964 11308 14280 11336
rect 13964 11296 13970 11308
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 15102 11296 15108 11348
rect 15160 11336 15166 11348
rect 15841 11339 15899 11345
rect 15841 11336 15853 11339
rect 15160 11308 15853 11336
rect 15160 11296 15166 11308
rect 15841 11305 15853 11308
rect 15887 11305 15899 11339
rect 15841 11299 15899 11305
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 16482 11336 16488 11348
rect 16356 11308 16488 11336
rect 16356 11296 16362 11308
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 18414 11336 18420 11348
rect 18375 11308 18420 11336
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 19521 11339 19579 11345
rect 19521 11336 19533 11339
rect 19392 11308 19533 11336
rect 19392 11296 19398 11308
rect 19521 11305 19533 11308
rect 19567 11305 19579 11339
rect 19521 11299 19579 11305
rect 22649 11339 22707 11345
rect 22649 11305 22661 11339
rect 22695 11336 22707 11339
rect 24210 11336 24216 11348
rect 22695 11308 24216 11336
rect 22695 11305 22707 11308
rect 22649 11299 22707 11305
rect 24210 11296 24216 11308
rect 24268 11296 24274 11348
rect 24578 11336 24584 11348
rect 24539 11308 24584 11336
rect 24578 11296 24584 11308
rect 24636 11296 24642 11348
rect 5951 11240 6960 11268
rect 8128 11240 10272 11268
rect 5951 11237 5963 11240
rect 5905 11231 5963 11237
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 4157 11203 4215 11209
rect 1995 11172 4108 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 1636 11104 1685 11132
rect 1636 11092 1642 11104
rect 1673 11101 1685 11104
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 3602 11064 3608 11076
rect 3174 11036 3608 11064
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 3326 10996 3332 11008
rect 2832 10968 3332 10996
rect 2832 10956 2838 10968
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 4080 11005 4108 11172
rect 4157 11169 4169 11203
rect 4203 11200 4215 11203
rect 4982 11200 4988 11212
rect 4203 11172 4988 11200
rect 4203 11169 4215 11172
rect 4157 11163 4215 11169
rect 4982 11160 4988 11172
rect 5040 11200 5046 11212
rect 6730 11200 6736 11212
rect 5040 11172 6736 11200
rect 5040 11160 5046 11172
rect 6730 11160 6736 11172
rect 6788 11200 6794 11212
rect 6825 11203 6883 11209
rect 6825 11200 6837 11203
rect 6788 11172 6837 11200
rect 6788 11160 6794 11172
rect 6825 11169 6837 11172
rect 6871 11169 6883 11203
rect 6825 11163 6883 11169
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11200 7159 11203
rect 7558 11200 7564 11212
rect 7147 11172 7564 11200
rect 7147 11169 7159 11172
rect 7101 11163 7159 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 8128 11200 8156 11240
rect 8570 11200 8576 11212
rect 7708 11172 8156 11200
rect 8531 11172 8576 11200
rect 7708 11160 7714 11172
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 9030 11160 9036 11212
rect 9088 11200 9094 11212
rect 10137 11203 10195 11209
rect 10137 11200 10149 11203
rect 9088 11172 10149 11200
rect 9088 11160 9094 11172
rect 10137 11169 10149 11172
rect 10183 11169 10195 11203
rect 10244 11200 10272 11240
rect 11514 11228 11520 11280
rect 11572 11268 11578 11280
rect 13078 11268 13084 11280
rect 11572 11240 13084 11268
rect 11572 11228 11578 11240
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 13725 11271 13783 11277
rect 13725 11237 13737 11271
rect 13771 11268 13783 11271
rect 15930 11268 15936 11280
rect 13771 11240 15936 11268
rect 13771 11237 13783 11240
rect 13725 11231 13783 11237
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 10410 11200 10416 11212
rect 10244 11172 10416 11200
rect 10137 11163 10195 11169
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 10962 11160 10968 11212
rect 11020 11200 11026 11212
rect 13906 11200 13912 11212
rect 11020 11172 13912 11200
rect 11020 11160 11026 11172
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11200 14979 11203
rect 15838 11200 15844 11212
rect 14967 11172 15844 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 16500 11200 16528 11296
rect 16500 11172 18736 11200
rect 5534 11092 5540 11144
rect 5592 11092 5598 11144
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9364 11104 9689 11132
rect 9364 11092 9370 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 12526 11132 12532 11144
rect 12487 11104 12532 11132
rect 9677 11095 9735 11101
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11132 12679 11135
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12667 11104 13093 11132
rect 12667 11101 12679 11104
rect 12621 11095 12679 11101
rect 13081 11101 13093 11104
rect 13127 11101 13139 11135
rect 13262 11132 13268 11144
rect 13223 11104 13268 11132
rect 13081 11095 13139 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 14826 11132 14832 11144
rect 14787 11104 14832 11132
rect 14826 11092 14832 11104
rect 14884 11092 14890 11144
rect 16022 11132 16028 11144
rect 15983 11104 16028 11132
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16482 11132 16488 11144
rect 16443 11104 16488 11132
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16666 11132 16672 11144
rect 16627 11104 16672 11132
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 18601 11135 18659 11141
rect 18601 11132 18613 11135
rect 18564 11104 18613 11132
rect 18564 11092 18570 11104
rect 18601 11101 18613 11104
rect 18647 11101 18659 11135
rect 18708 11132 18736 11172
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19518 11200 19524 11212
rect 19392 11172 19524 11200
rect 19392 11160 19398 11172
rect 19518 11160 19524 11172
rect 19576 11160 19582 11212
rect 20165 11203 20223 11209
rect 20165 11169 20177 11203
rect 20211 11200 20223 11203
rect 21269 11203 21327 11209
rect 21269 11200 21281 11203
rect 20211 11172 21281 11200
rect 20211 11169 20223 11172
rect 20165 11163 20223 11169
rect 21269 11169 21281 11172
rect 21315 11169 21327 11203
rect 21269 11163 21327 11169
rect 23293 11203 23351 11209
rect 23293 11169 23305 11203
rect 23339 11200 23351 11203
rect 24118 11200 24124 11212
rect 23339 11172 24124 11200
rect 23339 11169 23351 11172
rect 23293 11163 23351 11169
rect 24118 11160 24124 11172
rect 24176 11160 24182 11212
rect 24302 11160 24308 11212
rect 24360 11200 24366 11212
rect 24360 11172 29776 11200
rect 24360 11160 24366 11172
rect 19429 11135 19487 11141
rect 19429 11132 19441 11135
rect 18708 11104 19441 11132
rect 18601 11095 18659 11101
rect 19429 11101 19441 11104
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 20349 11135 20407 11141
rect 20349 11101 20361 11135
rect 20395 11132 20407 11135
rect 20806 11132 20812 11144
rect 20395 11104 20812 11132
rect 20395 11101 20407 11104
rect 20349 11095 20407 11101
rect 20806 11092 20812 11104
rect 20864 11092 20870 11144
rect 22830 11132 22836 11144
rect 22791 11104 22836 11132
rect 22830 11092 22836 11104
rect 22888 11092 22894 11144
rect 24762 11132 24768 11144
rect 24723 11104 24768 11132
rect 24762 11092 24768 11104
rect 24820 11092 24826 11144
rect 29748 11141 29776 11172
rect 29733 11135 29791 11141
rect 29733 11101 29745 11135
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 4430 11064 4436 11076
rect 4391 11036 4436 11064
rect 4430 11024 4436 11036
rect 4488 11024 4494 11076
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7064 11036 7590 11064
rect 7064 11024 7070 11036
rect 9122 11024 9128 11076
rect 9180 11064 9186 11076
rect 10410 11064 10416 11076
rect 9180 11036 10416 11064
rect 9180 11024 9186 11036
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 11698 11064 11704 11076
rect 11638 11036 11704 11064
rect 11698 11024 11704 11036
rect 11756 11024 11762 11076
rect 17770 11064 17776 11076
rect 17731 11036 17776 11064
rect 17770 11024 17776 11036
rect 17828 11024 17834 11076
rect 29825 11067 29883 11073
rect 29825 11033 29837 11067
rect 29871 11064 29883 11067
rect 30834 11064 30840 11076
rect 29871 11036 30840 11064
rect 29871 11033 29883 11036
rect 29825 11027 29883 11033
rect 30834 11024 30840 11036
rect 30892 11024 30898 11076
rect 4065 10999 4123 11005
rect 4065 10965 4077 10999
rect 4111 10996 4123 10999
rect 9674 10996 9680 11008
rect 4111 10968 9680 10996
rect 4111 10965 4123 10968
rect 4065 10959 4123 10965
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 11885 10999 11943 11005
rect 11885 10996 11897 10999
rect 9824 10968 11897 10996
rect 9824 10956 9830 10968
rect 11885 10965 11897 10968
rect 11931 10965 11943 10999
rect 11885 10959 11943 10965
rect 12158 10956 12164 11008
rect 12216 10996 12222 11008
rect 13170 10996 13176 11008
rect 12216 10968 13176 10996
rect 12216 10956 12222 10968
rect 13170 10956 13176 10968
rect 13228 10956 13234 11008
rect 15562 10956 15568 11008
rect 15620 10996 15626 11008
rect 16758 10996 16764 11008
rect 15620 10968 16764 10996
rect 15620 10956 15626 10968
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 17129 10999 17187 11005
rect 17129 10965 17141 10999
rect 17175 10996 17187 10999
rect 17218 10996 17224 11008
rect 17175 10968 17224 10996
rect 17175 10965 17187 10968
rect 17129 10959 17187 10965
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 20809 10999 20867 11005
rect 20809 10996 20821 10999
rect 20772 10968 20821 10996
rect 20772 10956 20778 10968
rect 20809 10965 20821 10968
rect 20855 10996 20867 10999
rect 21082 10996 21088 11008
rect 20855 10968 21088 10996
rect 20855 10965 20867 10968
rect 20809 10959 20867 10965
rect 21082 10956 21088 10968
rect 21140 10956 21146 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 1762 10792 1768 10804
rect 1719 10764 1768 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 4798 10792 4804 10804
rect 2363 10764 4804 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 8386 10792 8392 10804
rect 5859 10764 8392 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 9122 10792 9128 10804
rect 8527 10764 9128 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 14458 10792 14464 10804
rect 9646 10764 14464 10792
rect 2774 10724 2780 10736
rect 1596 10696 2780 10724
rect 1596 10665 1624 10696
rect 2774 10684 2780 10696
rect 2832 10724 2838 10736
rect 3142 10724 3148 10736
rect 2832 10696 3148 10724
rect 2832 10684 2838 10696
rect 3142 10684 3148 10696
rect 3200 10684 3206 10736
rect 5442 10724 5448 10736
rect 4370 10696 5448 10724
rect 5442 10684 5448 10696
rect 5500 10684 5506 10736
rect 7009 10727 7067 10733
rect 7009 10693 7021 10727
rect 7055 10724 7067 10727
rect 7098 10724 7104 10736
rect 7055 10696 7104 10724
rect 7055 10693 7067 10696
rect 7009 10687 7067 10693
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 9646 10724 9674 10764
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 15565 10795 15623 10801
rect 15565 10761 15577 10795
rect 15611 10792 15623 10795
rect 15746 10792 15752 10804
rect 15611 10764 15752 10792
rect 15611 10761 15623 10764
rect 15565 10755 15623 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 16172 10764 16221 10792
rect 16172 10752 16178 10764
rect 16209 10761 16221 10764
rect 16255 10761 16267 10795
rect 16209 10755 16267 10761
rect 18598 10752 18604 10804
rect 18656 10792 18662 10804
rect 18877 10795 18935 10801
rect 18877 10792 18889 10795
rect 18656 10764 18889 10792
rect 18656 10752 18662 10764
rect 18877 10761 18889 10764
rect 18923 10761 18935 10795
rect 19426 10792 19432 10804
rect 19387 10764 19432 10792
rect 18877 10755 18935 10761
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 20162 10752 20168 10804
rect 20220 10792 20226 10804
rect 20257 10795 20315 10801
rect 20257 10792 20269 10795
rect 20220 10764 20269 10792
rect 20220 10752 20226 10764
rect 20257 10761 20269 10764
rect 20303 10761 20315 10795
rect 20806 10792 20812 10804
rect 20767 10764 20812 10792
rect 20257 10755 20315 10761
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 20990 10752 20996 10804
rect 21048 10792 21054 10804
rect 23198 10792 23204 10804
rect 21048 10764 23204 10792
rect 21048 10752 21054 10764
rect 23198 10752 23204 10764
rect 23256 10752 23262 10804
rect 23385 10795 23443 10801
rect 23385 10761 23397 10795
rect 23431 10792 23443 10795
rect 23842 10792 23848 10804
rect 23431 10764 23848 10792
rect 23431 10761 23443 10764
rect 23385 10755 23443 10761
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 24029 10795 24087 10801
rect 24029 10761 24041 10795
rect 24075 10792 24087 10795
rect 24762 10792 24768 10804
rect 24075 10764 24768 10792
rect 24075 10761 24087 10764
rect 24029 10755 24087 10761
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 27249 10795 27307 10801
rect 27249 10761 27261 10795
rect 27295 10792 27307 10795
rect 30374 10792 30380 10804
rect 27295 10764 30380 10792
rect 27295 10761 27307 10764
rect 27249 10755 27307 10761
rect 30374 10752 30380 10764
rect 30432 10752 30438 10804
rect 8234 10696 9674 10724
rect 10686 10684 10692 10736
rect 10744 10684 10750 10736
rect 12434 10684 12440 10736
rect 12492 10684 12498 10736
rect 13446 10684 13452 10736
rect 13504 10724 13510 10736
rect 16850 10724 16856 10736
rect 13504 10696 16856 10724
rect 13504 10684 13510 10696
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 16942 10684 16948 10736
rect 17000 10724 17006 10736
rect 20438 10724 20444 10736
rect 17000 10696 20444 10724
rect 17000 10684 17006 10696
rect 20438 10684 20444 10696
rect 20496 10684 20502 10736
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 2225 10659 2283 10665
rect 2225 10656 2237 10659
rect 2188 10628 2237 10656
rect 2188 10616 2194 10628
rect 2225 10625 2237 10628
rect 2271 10656 2283 10659
rect 2314 10656 2320 10668
rect 2271 10628 2320 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 5166 10656 5172 10668
rect 5127 10628 5172 10656
rect 5166 10616 5172 10628
rect 5224 10616 5230 10668
rect 5994 10656 6000 10668
rect 5955 10628 6000 10656
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 6730 10656 6736 10668
rect 6691 10628 6736 10656
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 9122 10656 9128 10668
rect 8904 10628 9128 10656
rect 8904 10616 8910 10628
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 14369 10659 14427 10665
rect 14369 10625 14381 10659
rect 14415 10656 14427 10659
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 14415 10628 14841 10656
rect 14415 10625 14427 10628
rect 14369 10619 14427 10625
rect 14829 10625 14841 10628
rect 14875 10625 14887 10659
rect 14829 10619 14887 10625
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2746 10560 2881 10588
rect 1578 10480 1584 10532
rect 1636 10520 1642 10532
rect 2746 10520 2774 10560
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 3142 10588 3148 10600
rect 3103 10560 3148 10588
rect 2869 10551 2927 10557
rect 3142 10548 3148 10560
rect 3200 10548 3206 10600
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10588 5319 10591
rect 8754 10588 8760 10600
rect 5307 10560 8760 10588
rect 5307 10557 5319 10560
rect 5261 10551 5319 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9030 10548 9036 10600
rect 9088 10588 9094 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 9088 10560 9413 10588
rect 9088 10548 9094 10560
rect 9401 10557 9413 10560
rect 9447 10588 9459 10591
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 9447 10560 11713 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 11701 10557 11713 10560
rect 11747 10557 11759 10591
rect 11977 10591 12035 10597
rect 11977 10588 11989 10591
rect 11701 10551 11759 10557
rect 11808 10560 11989 10588
rect 8846 10520 8852 10532
rect 1636 10492 2774 10520
rect 8036 10492 8852 10520
rect 1636 10480 1642 10492
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 4617 10455 4675 10461
rect 4617 10452 4629 10455
rect 4488 10424 4629 10452
rect 4488 10412 4494 10424
rect 4617 10421 4629 10424
rect 4663 10452 4675 10455
rect 4798 10452 4804 10464
rect 4663 10424 4804 10452
rect 4663 10421 4675 10424
rect 4617 10415 4675 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 8036 10452 8064 10492
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 11146 10520 11152 10532
rect 11107 10492 11152 10520
rect 11146 10480 11152 10492
rect 11204 10520 11210 10532
rect 11808 10520 11836 10560
rect 11977 10557 11989 10560
rect 12023 10557 12035 10591
rect 11977 10551 12035 10557
rect 13170 10548 13176 10600
rect 13228 10588 13234 10600
rect 14384 10588 14412 10619
rect 15102 10616 15108 10668
rect 15160 10656 15166 10668
rect 15473 10659 15531 10665
rect 15160 10654 15424 10656
rect 15473 10654 15485 10659
rect 15160 10628 15485 10654
rect 15160 10616 15166 10628
rect 15396 10626 15485 10628
rect 15473 10625 15485 10626
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 16022 10616 16028 10668
rect 16080 10656 16086 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 16080 10628 16129 10656
rect 16080 10616 16086 10628
rect 16117 10625 16129 10628
rect 16163 10656 16175 10659
rect 16390 10656 16396 10668
rect 16163 10628 16396 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 16390 10616 16396 10628
rect 16448 10616 16454 10668
rect 20165 10659 20223 10665
rect 20165 10656 20177 10659
rect 16500 10628 20177 10656
rect 16500 10588 16528 10628
rect 20165 10625 20177 10628
rect 20211 10656 20223 10659
rect 20346 10656 20352 10668
rect 20211 10628 20352 10656
rect 20211 10625 20223 10628
rect 20165 10619 20223 10625
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 20990 10656 20996 10668
rect 20951 10628 20996 10656
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 21082 10616 21088 10668
rect 21140 10656 21146 10668
rect 22649 10659 22707 10665
rect 22649 10656 22661 10659
rect 21140 10628 22661 10656
rect 21140 10616 21146 10628
rect 22649 10625 22661 10628
rect 22695 10625 22707 10659
rect 23566 10656 23572 10668
rect 23527 10628 23572 10656
rect 22649 10619 22707 10625
rect 23566 10616 23572 10628
rect 23624 10616 23630 10668
rect 23658 10616 23664 10668
rect 23716 10656 23722 10668
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23716 10628 24225 10656
rect 23716 10616 23722 10628
rect 24213 10625 24225 10628
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 24912 10628 27169 10656
rect 24912 10616 24918 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 30834 10616 30840 10668
rect 30892 10656 30898 10668
rect 35069 10659 35127 10665
rect 35069 10656 35081 10659
rect 30892 10628 35081 10656
rect 30892 10616 30898 10628
rect 35069 10625 35081 10628
rect 35115 10625 35127 10659
rect 36446 10656 36452 10668
rect 36407 10628 36452 10656
rect 35069 10619 35127 10625
rect 36446 10616 36452 10628
rect 36504 10616 36510 10668
rect 38013 10659 38071 10665
rect 38013 10625 38025 10659
rect 38059 10625 38071 10659
rect 38013 10619 38071 10625
rect 13228 10560 14412 10588
rect 14476 10560 16528 10588
rect 13228 10548 13234 10560
rect 14476 10520 14504 10560
rect 16850 10548 16856 10600
rect 16908 10588 16914 10600
rect 17037 10591 17095 10597
rect 16908 10560 16953 10588
rect 16908 10548 16914 10560
rect 17037 10557 17049 10591
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 18233 10591 18291 10597
rect 18233 10557 18245 10591
rect 18279 10557 18291 10591
rect 18233 10551 18291 10557
rect 18417 10591 18475 10597
rect 18417 10557 18429 10591
rect 18463 10588 18475 10591
rect 18598 10588 18604 10600
rect 18463 10560 18604 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 11204 10492 11836 10520
rect 13004 10492 14504 10520
rect 14921 10523 14979 10529
rect 11204 10480 11210 10492
rect 9674 10461 9680 10464
rect 5132 10424 8064 10452
rect 9658 10455 9680 10461
rect 5132 10412 5138 10424
rect 9658 10421 9670 10455
rect 9658 10415 9680 10421
rect 9674 10412 9680 10415
rect 9732 10412 9738 10464
rect 10410 10412 10416 10464
rect 10468 10452 10474 10464
rect 13004 10452 13032 10492
rect 14921 10489 14933 10523
rect 14967 10520 14979 10523
rect 17052 10520 17080 10551
rect 17218 10520 17224 10532
rect 14967 10492 17080 10520
rect 17179 10492 17224 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 17218 10480 17224 10492
rect 17276 10480 17282 10532
rect 18248 10520 18276 10551
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 38028 10588 38056 10619
rect 35866 10560 38056 10588
rect 19150 10520 19156 10532
rect 18248 10492 19156 10520
rect 19150 10480 19156 10492
rect 19208 10480 19214 10532
rect 22741 10523 22799 10529
rect 22741 10489 22753 10523
rect 22787 10520 22799 10523
rect 24762 10520 24768 10532
rect 22787 10492 24768 10520
rect 22787 10489 22799 10492
rect 22741 10483 22799 10489
rect 24762 10480 24768 10492
rect 24820 10480 24826 10532
rect 34885 10523 34943 10529
rect 34885 10489 34897 10523
rect 34931 10520 34943 10523
rect 35866 10520 35894 10560
rect 34931 10492 35894 10520
rect 34931 10489 34943 10492
rect 34885 10483 34943 10489
rect 10468 10424 13032 10452
rect 13449 10455 13507 10461
rect 10468 10412 10474 10424
rect 13449 10421 13461 10455
rect 13495 10452 13507 10455
rect 13630 10452 13636 10464
rect 13495 10424 13636 10452
rect 13495 10421 13507 10424
rect 13449 10415 13507 10421
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 15838 10452 15844 10464
rect 14231 10424 15844 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 36265 10455 36323 10461
rect 36265 10421 36277 10455
rect 36311 10452 36323 10455
rect 38010 10452 38016 10464
rect 36311 10424 38016 10452
rect 36311 10421 36323 10424
rect 36265 10415 36323 10421
rect 38010 10412 38016 10424
rect 38068 10412 38074 10464
rect 38194 10452 38200 10464
rect 38155 10424 38200 10452
rect 38194 10412 38200 10424
rect 38252 10412 38258 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 5350 10248 5356 10260
rect 4663 10220 5356 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 6546 10248 6552 10260
rect 5460 10220 6552 10248
rect 5074 10180 5080 10192
rect 3804 10152 5080 10180
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 3804 10112 3832 10152
rect 5074 10140 5080 10152
rect 5132 10140 5138 10192
rect 3970 10112 3976 10124
rect 1995 10084 3832 10112
rect 3931 10084 3976 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 3970 10072 3976 10084
rect 4028 10072 4034 10124
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 4157 10115 4215 10121
rect 4157 10112 4169 10115
rect 4120 10084 4169 10112
rect 4120 10072 4126 10084
rect 4157 10081 4169 10084
rect 4203 10081 4215 10115
rect 4157 10075 4215 10081
rect 1578 10004 1584 10056
rect 1636 10044 1642 10056
rect 5460 10053 5488 10220
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7650 10248 7656 10260
rect 7432 10220 7656 10248
rect 7432 10208 7438 10220
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 13078 10248 13084 10260
rect 12124 10220 13084 10248
rect 12124 10208 12130 10220
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 13262 10208 13268 10260
rect 13320 10248 13326 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13320 10220 13553 10248
rect 13320 10208 13326 10220
rect 13541 10217 13553 10220
rect 13587 10217 13599 10251
rect 13541 10211 13599 10217
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14458 10248 14464 10260
rect 13872 10220 14464 10248
rect 13872 10208 13878 10220
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 14642 10248 14648 10260
rect 14603 10220 14648 10248
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 15102 10208 15108 10260
rect 15160 10248 15166 10260
rect 15562 10248 15568 10260
rect 15160 10220 15568 10248
rect 15160 10208 15166 10220
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 16666 10248 16672 10260
rect 15703 10220 16672 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 20165 10251 20223 10257
rect 20165 10217 20177 10251
rect 20211 10248 20223 10251
rect 20990 10248 20996 10260
rect 20211 10220 20996 10248
rect 20211 10217 20223 10220
rect 20165 10211 20223 10217
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 23474 10248 23480 10260
rect 23435 10220 23480 10248
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 8481 10183 8539 10189
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 11882 10180 11888 10192
rect 8527 10152 10272 10180
rect 11795 10152 11888 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 6730 10112 6736 10124
rect 5951 10084 6736 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 9088 10084 10149 10112
rect 9088 10072 9094 10084
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 10244 10112 10272 10152
rect 11882 10140 11888 10152
rect 11940 10180 11946 10192
rect 15930 10180 15936 10192
rect 11940 10152 14596 10180
rect 11940 10140 11946 10152
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 10244 10084 12541 10112
rect 10137 10075 10195 10081
rect 12529 10081 12541 10084
rect 12575 10081 12587 10115
rect 12529 10075 12587 10081
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 13170 10112 13176 10124
rect 12860 10084 13176 10112
rect 12860 10072 12866 10084
rect 13170 10072 13176 10084
rect 13228 10072 13234 10124
rect 1673 10047 1731 10053
rect 1673 10044 1685 10047
rect 1636 10016 1685 10044
rect 1636 10004 1642 10016
rect 1673 10013 1685 10016
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8938 10044 8944 10056
rect 8435 10016 8944 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8938 10004 8944 10016
rect 8996 10044 9002 10056
rect 9306 10044 9312 10056
rect 8996 10016 9312 10044
rect 8996 10004 9002 10016
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9456 10016 9689 10044
rect 9456 10004 9462 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12345 10047 12403 10053
rect 12345 10044 12357 10047
rect 12032 10016 12357 10044
rect 12032 10004 12038 10016
rect 12345 10013 12357 10016
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10044 13507 10047
rect 13814 10044 13820 10056
rect 13495 10016 13820 10044
rect 13495 10013 13507 10016
rect 13449 10007 13507 10013
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 14274 10044 14280 10056
rect 14235 10016 14280 10044
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 5534 9976 5540 9988
rect 3174 9948 5540 9976
rect 5534 9936 5540 9948
rect 5592 9936 5598 9988
rect 6181 9979 6239 9985
rect 6181 9945 6193 9979
rect 6227 9976 6239 9979
rect 6454 9976 6460 9988
rect 6227 9948 6460 9976
rect 6227 9945 6239 9948
rect 6181 9939 6239 9945
rect 6454 9936 6460 9948
rect 6512 9936 6518 9988
rect 6914 9936 6920 9988
rect 6972 9936 6978 9988
rect 8294 9976 8300 9988
rect 7484 9948 8300 9976
rect 2590 9868 2596 9920
rect 2648 9908 2654 9920
rect 3421 9911 3479 9917
rect 3421 9908 3433 9911
rect 2648 9880 3433 9908
rect 2648 9868 2654 9880
rect 3421 9877 3433 9880
rect 3467 9877 3479 9911
rect 3421 9871 3479 9877
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9908 5319 9911
rect 7484 9908 7512 9948
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 10134 9936 10140 9988
rect 10192 9976 10198 9988
rect 10413 9979 10471 9985
rect 10413 9976 10425 9979
rect 10192 9948 10425 9976
rect 10192 9936 10198 9948
rect 10413 9945 10425 9948
rect 10459 9945 10471 9979
rect 11698 9976 11704 9988
rect 11638 9948 11704 9976
rect 10413 9939 10471 9945
rect 11698 9936 11704 9948
rect 11756 9936 11762 9988
rect 14476 9976 14504 10007
rect 11808 9948 14504 9976
rect 14568 9976 14596 10152
rect 15864 10152 15936 10180
rect 15864 10053 15892 10152
rect 15930 10140 15936 10152
rect 15988 10140 15994 10192
rect 16206 10140 16212 10192
rect 16264 10180 16270 10192
rect 17589 10183 17647 10189
rect 17589 10180 17601 10183
rect 16264 10152 17601 10180
rect 16264 10140 16270 10152
rect 17589 10149 17601 10152
rect 17635 10149 17647 10183
rect 17589 10143 17647 10149
rect 18782 10140 18788 10192
rect 18840 10180 18846 10192
rect 19613 10183 19671 10189
rect 18840 10152 19472 10180
rect 18840 10140 18846 10152
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 16482 10112 16488 10124
rect 16347 10084 16488 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 17037 10115 17095 10121
rect 17037 10081 17049 10115
rect 17083 10112 17095 10115
rect 19334 10112 19340 10124
rect 17083 10084 19340 10112
rect 17083 10081 17095 10084
rect 17037 10075 17095 10081
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19444 10112 19472 10152
rect 19613 10149 19625 10183
rect 19659 10180 19671 10183
rect 20254 10180 20260 10192
rect 19659 10152 20260 10180
rect 19659 10149 19671 10152
rect 19613 10143 19671 10149
rect 20254 10140 20260 10152
rect 20312 10140 20318 10192
rect 33965 10115 34023 10121
rect 33965 10112 33977 10115
rect 19444 10084 33977 10112
rect 33965 10081 33977 10084
rect 34011 10081 34023 10115
rect 33965 10075 34023 10081
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 18506 10044 18512 10056
rect 18467 10016 18512 10044
rect 15841 10007 15899 10013
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10044 19579 10047
rect 20254 10044 20260 10056
rect 19567 10016 20260 10044
rect 19567 10013 19579 10016
rect 19521 10007 19579 10013
rect 20254 10004 20260 10016
rect 20312 10004 20318 10056
rect 20346 10004 20352 10056
rect 20404 10044 20410 10056
rect 23109 10047 23167 10053
rect 20404 10016 20449 10044
rect 20404 10004 20410 10016
rect 23109 10013 23121 10047
rect 23155 10013 23167 10047
rect 23290 10044 23296 10056
rect 23251 10016 23296 10044
rect 23109 10007 23167 10013
rect 16758 9976 16764 9988
rect 14568 9948 16764 9976
rect 5307 9880 7512 9908
rect 5307 9877 5319 9880
rect 5261 9871 5319 9877
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 9122 9908 9128 9920
rect 8720 9880 9128 9908
rect 8720 9868 8726 9880
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9493 9911 9551 9917
rect 9493 9877 9505 9911
rect 9539 9908 9551 9911
rect 11808 9908 11836 9948
rect 16758 9936 16764 9948
rect 16816 9936 16822 9988
rect 17126 9936 17132 9988
rect 17184 9976 17190 9988
rect 23124 9976 23152 10007
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 33873 10047 33931 10053
rect 33873 10013 33885 10047
rect 33919 10044 33931 10047
rect 36906 10044 36912 10056
rect 33919 10016 36912 10044
rect 33919 10013 33931 10016
rect 33873 10007 33931 10013
rect 36906 10004 36912 10016
rect 36964 10004 36970 10056
rect 29546 9976 29552 9988
rect 17184 9948 17229 9976
rect 23124 9948 29552 9976
rect 17184 9936 17190 9948
rect 29546 9936 29552 9948
rect 29604 9936 29610 9988
rect 9539 9880 11836 9908
rect 12989 9911 13047 9917
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 12989 9877 13001 9911
rect 13035 9908 13047 9911
rect 14090 9908 14096 9920
rect 13035 9880 14096 9908
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14366 9868 14372 9920
rect 14424 9908 14430 9920
rect 16114 9908 16120 9920
rect 14424 9880 16120 9908
rect 14424 9868 14430 9880
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 7282 9704 7288 9716
rect 4724 9676 5672 9704
rect 3418 9636 3424 9648
rect 3082 9608 3424 9636
rect 3418 9596 3424 9608
rect 3476 9596 3482 9648
rect 4341 9639 4399 9645
rect 4341 9605 4353 9639
rect 4387 9636 4399 9639
rect 4724 9636 4752 9676
rect 4387 9608 4752 9636
rect 4387 9605 4399 9608
rect 4341 9599 4399 9605
rect 4890 9596 4896 9648
rect 4948 9596 4954 9648
rect 5644 9636 5672 9676
rect 6840 9676 7288 9704
rect 6840 9636 6868 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 8904 9676 11652 9704
rect 8904 9664 8910 9676
rect 5644 9608 6868 9636
rect 6917 9639 6975 9645
rect 6917 9605 6929 9639
rect 6963 9636 6975 9639
rect 7190 9636 7196 9648
rect 6963 9608 7196 9636
rect 6963 9605 6975 9608
rect 6917 9599 6975 9605
rect 7190 9596 7196 9608
rect 7248 9596 7254 9648
rect 8202 9636 8208 9648
rect 8142 9608 8208 9636
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 8570 9596 8576 9648
rect 8628 9636 8634 9648
rect 9309 9639 9367 9645
rect 9309 9636 9321 9639
rect 8628 9608 9321 9636
rect 8628 9596 8634 9608
rect 9309 9605 9321 9608
rect 9355 9605 9367 9639
rect 9309 9599 9367 9605
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 11624 9636 11652 9676
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 11756 9676 13584 9704
rect 11756 9664 11762 9676
rect 12066 9636 12072 9648
rect 9640 9608 9798 9636
rect 11624 9608 12072 9636
rect 9640 9596 9646 9608
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 12250 9636 12256 9648
rect 12211 9608 12256 9636
rect 12250 9596 12256 9608
rect 12308 9596 12314 9648
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 13556 9636 13584 9676
rect 14274 9664 14280 9716
rect 14332 9704 14338 9716
rect 18322 9704 18328 9716
rect 14332 9676 18328 9704
rect 14332 9664 14338 9676
rect 18322 9664 18328 9676
rect 18380 9664 18386 9716
rect 19058 9664 19064 9716
rect 19116 9704 19122 9716
rect 21542 9704 21548 9716
rect 19116 9676 21548 9704
rect 19116 9664 19122 9676
rect 21542 9664 21548 9676
rect 21600 9664 21606 9716
rect 23290 9704 23296 9716
rect 23251 9676 23296 9704
rect 23290 9664 23296 9676
rect 23348 9664 23354 9716
rect 14366 9636 14372 9648
rect 12860 9608 13492 9636
rect 13556 9608 14372 9636
rect 12860 9596 12866 9608
rect 6638 9568 6644 9580
rect 6599 9540 6644 9568
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 13464 9577 13492 9608
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 14642 9596 14648 9648
rect 14700 9636 14706 9648
rect 15749 9639 15807 9645
rect 15749 9636 15761 9639
rect 14700 9608 15148 9636
rect 14700 9596 14706 9608
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 10652 9540 12173 9568
rect 10652 9528 10658 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13449 9571 13507 9577
rect 13449 9537 13461 9571
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 14826 9568 14832 9580
rect 14323 9540 14832 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 1854 9500 1860 9512
rect 1815 9472 1860 9500
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9469 3663 9503
rect 3605 9463 3663 9469
rect 3620 9432 3648 9463
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4065 9503 4123 9509
rect 4065 9500 4077 9503
rect 4028 9472 4077 9500
rect 4028 9460 4034 9472
rect 4065 9469 4077 9472
rect 4111 9469 4123 9503
rect 8389 9503 8447 9509
rect 4065 9463 4123 9469
rect 4172 9472 7972 9500
rect 4172 9432 4200 9472
rect 3620 9404 4200 9432
rect 7944 9432 7972 9472
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8478 9500 8484 9512
rect 8435 9472 8484 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 12526 9500 12532 9512
rect 9140 9472 12532 9500
rect 9140 9432 9168 9472
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 13004 9500 13032 9531
rect 13004 9472 14136 9500
rect 7944 9404 9168 9432
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 3620 9364 3648 9404
rect 10410 9392 10416 9444
rect 10468 9432 10474 9444
rect 12342 9432 12348 9444
rect 10468 9404 12348 9432
rect 10468 9392 10474 9404
rect 12342 9392 12348 9404
rect 12400 9432 12406 9444
rect 14108 9441 14136 9472
rect 14093 9435 14151 9441
rect 12400 9404 14044 9432
rect 12400 9392 12406 9404
rect 1912 9336 3648 9364
rect 1912 9324 1918 9336
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 5074 9364 5080 9376
rect 4580 9336 5080 9364
rect 4580 9324 4586 9336
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5810 9364 5816 9376
rect 5771 9336 5816 9364
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 9030 9364 9036 9376
rect 6788 9336 9036 9364
rect 6788 9324 6794 9336
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9306 9324 9312 9376
rect 9364 9364 9370 9376
rect 10781 9367 10839 9373
rect 10781 9364 10793 9367
rect 9364 9336 10793 9364
rect 9364 9324 9370 9336
rect 10781 9333 10793 9336
rect 10827 9333 10839 9367
rect 10781 9327 10839 9333
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 11422 9364 11428 9376
rect 11204 9336 11428 9364
rect 11204 9324 11210 9336
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 13262 9364 13268 9376
rect 12851 9336 13268 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 13504 9336 13553 9364
rect 13504 9324 13510 9336
rect 13541 9333 13553 9336
rect 13587 9333 13599 9367
rect 14016 9364 14044 9404
rect 14093 9401 14105 9435
rect 14139 9401 14151 9435
rect 14093 9395 14151 9401
rect 14292 9364 14320 9531
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 15120 9577 15148 9608
rect 15212 9608 15761 9636
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 15010 9460 15016 9512
rect 15068 9500 15074 9512
rect 15212 9500 15240 9608
rect 15749 9605 15761 9608
rect 15795 9605 15807 9639
rect 15749 9599 15807 9605
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 18046 9636 18052 9648
rect 17083 9608 18052 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18325 9571 18383 9577
rect 18325 9568 18337 9571
rect 17644 9540 18337 9568
rect 17644 9528 17650 9540
rect 18325 9537 18337 9540
rect 18371 9537 18383 9571
rect 23201 9571 23259 9577
rect 23201 9568 23213 9571
rect 18325 9531 18383 9537
rect 22204 9540 23213 9568
rect 22204 9512 22232 9540
rect 23201 9537 23213 9540
rect 23247 9537 23259 9571
rect 23201 9531 23259 9537
rect 15068 9472 15240 9500
rect 15068 9460 15074 9472
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 15657 9503 15715 9509
rect 15657 9500 15669 9503
rect 15344 9472 15669 9500
rect 15344 9460 15350 9472
rect 15657 9469 15669 9472
rect 15703 9469 15715 9503
rect 15657 9463 15715 9469
rect 16945 9503 17003 9509
rect 16945 9469 16957 9503
rect 16991 9500 17003 9503
rect 17034 9500 17040 9512
rect 16991 9472 17040 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 17218 9460 17224 9512
rect 17276 9500 17282 9512
rect 22186 9500 22192 9512
rect 17276 9472 22192 9500
rect 17276 9460 17282 9472
rect 22186 9460 22192 9472
rect 22244 9460 22250 9512
rect 16209 9435 16267 9441
rect 16209 9401 16221 9435
rect 16255 9432 16267 9435
rect 17497 9435 17555 9441
rect 17497 9432 17509 9435
rect 16255 9404 17509 9432
rect 16255 9401 16267 9404
rect 16209 9395 16267 9401
rect 17497 9401 17509 9404
rect 17543 9432 17555 9435
rect 28258 9432 28264 9444
rect 17543 9404 28264 9432
rect 17543 9401 17555 9404
rect 17497 9395 17555 9401
rect 28258 9392 28264 9404
rect 28316 9392 28322 9444
rect 14016 9336 14320 9364
rect 14921 9367 14979 9373
rect 13541 9327 13599 9333
rect 14921 9333 14933 9367
rect 14967 9364 14979 9367
rect 15194 9364 15200 9376
rect 14967 9336 15200 9364
rect 14967 9333 14979 9336
rect 14921 9327 14979 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 18417 9367 18475 9373
rect 18417 9333 18429 9367
rect 18463 9364 18475 9367
rect 18782 9364 18788 9376
rect 18463 9336 18788 9364
rect 18463 9333 18475 9336
rect 18417 9327 18475 9333
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 5718 9160 5724 9172
rect 2004 9132 5580 9160
rect 5679 9132 5724 9160
rect 2004 9120 2010 9132
rect 3326 9092 3332 9104
rect 3287 9064 3332 9092
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 5552 9092 5580 9132
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 9214 9160 9220 9172
rect 5960 9132 9220 9160
rect 5960 9120 5966 9132
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9398 9160 9404 9172
rect 9359 9132 9404 9160
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 11054 9160 11060 9172
rect 9508 9132 11060 9160
rect 5552 9064 6960 9092
rect 3970 9024 3976 9036
rect 1596 8996 3976 9024
rect 1596 8968 1624 8996
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 5258 9024 5264 9036
rect 4295 8996 5264 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 6932 9024 6960 9064
rect 8478 9052 8484 9104
rect 8536 9092 8542 9104
rect 9508 9092 9536 9132
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 12437 9163 12495 9169
rect 12437 9129 12449 9163
rect 12483 9160 12495 9163
rect 14642 9160 14648 9172
rect 12483 9132 14648 9160
rect 12483 9129 12495 9132
rect 12437 9123 12495 9129
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 16669 9163 16727 9169
rect 15804 9132 16620 9160
rect 15804 9120 15810 9132
rect 8536 9064 9536 9092
rect 8536 9052 8542 9064
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 11793 9095 11851 9101
rect 11793 9092 11805 9095
rect 11664 9064 11805 9092
rect 11664 9052 11670 9064
rect 11793 9061 11805 9064
rect 11839 9061 11851 9095
rect 13538 9092 13544 9104
rect 11793 9055 11851 9061
rect 13096 9064 13544 9092
rect 9858 9024 9864 9036
rect 6932 8996 9864 9024
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 10318 9024 10324 9036
rect 10279 8996 10324 9024
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 13096 9033 13124 9064
rect 13538 9052 13544 9064
rect 13596 9052 13602 9104
rect 14829 9095 14887 9101
rect 14829 9061 14841 9095
rect 14875 9092 14887 9095
rect 15470 9092 15476 9104
rect 14875 9064 15476 9092
rect 14875 9061 14887 9064
rect 14829 9055 14887 9061
rect 15470 9052 15476 9064
rect 15528 9092 15534 9104
rect 16592 9092 16620 9132
rect 16669 9129 16681 9163
rect 16715 9160 16727 9163
rect 16850 9160 16856 9172
rect 16715 9132 16856 9160
rect 16715 9129 16727 9132
rect 16669 9123 16727 9129
rect 16850 9120 16856 9132
rect 16908 9160 16914 9172
rect 17402 9160 17408 9172
rect 16908 9132 17408 9160
rect 16908 9120 16914 9132
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 18046 9160 18052 9172
rect 18007 9132 18052 9160
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 21818 9120 21824 9172
rect 21876 9120 21882 9172
rect 21836 9092 21864 9120
rect 22373 9095 22431 9101
rect 22373 9092 22385 9095
rect 15528 9064 16068 9092
rect 16592 9064 22385 9092
rect 15528 9052 15534 9064
rect 13081 9027 13139 9033
rect 13081 9024 13093 9027
rect 12406 8996 13093 9024
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6788 8928 6837 8956
rect 6788 8916 6794 8928
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 8938 8956 8944 8968
rect 8812 8928 8944 8956
rect 8812 8916 8818 8928
rect 8938 8916 8944 8928
rect 8996 8956 9002 8968
rect 9585 8959 9643 8965
rect 9585 8956 9597 8959
rect 8996 8928 9597 8956
rect 8996 8916 9002 8928
rect 9585 8925 9597 8928
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 9824 8928 10057 8956
rect 9824 8916 9830 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 12406 8956 12434 8996
rect 13081 8993 13093 8996
rect 13127 8993 13139 9027
rect 13262 9024 13268 9036
rect 13223 8996 13268 9024
rect 13081 8987 13139 8993
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 16040 9033 16068 9064
rect 22373 9061 22385 9064
rect 22419 9061 22431 9095
rect 22373 9055 22431 9061
rect 16025 9027 16083 9033
rect 13372 8996 15516 9024
rect 11940 8928 12434 8956
rect 12621 8959 12679 8965
rect 11940 8916 11946 8928
rect 12621 8925 12633 8959
rect 12667 8956 12679 8959
rect 13372 8956 13400 8996
rect 15488 8968 15516 8996
rect 16025 8993 16037 9027
rect 16071 8993 16083 9027
rect 16206 9024 16212 9036
rect 16167 8996 16212 9024
rect 16025 8987 16083 8993
rect 16206 8984 16212 8996
rect 16264 8984 16270 9036
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 20070 9024 20076 9036
rect 16356 8996 20076 9024
rect 16356 8984 16362 8996
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 21821 9027 21879 9033
rect 21821 8993 21833 9027
rect 21867 9024 21879 9027
rect 24949 9027 25007 9033
rect 24949 9024 24961 9027
rect 21867 8996 24961 9024
rect 21867 8993 21879 8996
rect 21821 8987 21879 8993
rect 24949 8993 24961 8996
rect 24995 8993 25007 9027
rect 24949 8987 25007 8993
rect 12667 8928 13400 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 14642 8916 14648 8968
rect 14700 8956 14706 8968
rect 14737 8959 14795 8965
rect 14737 8956 14749 8959
rect 14700 8928 14749 8956
rect 14700 8916 14706 8928
rect 14737 8925 14749 8928
rect 14783 8925 14795 8959
rect 15378 8956 15384 8968
rect 15339 8928 15384 8956
rect 14737 8919 14795 8925
rect 15378 8916 15384 8928
rect 15436 8916 15442 8968
rect 15470 8916 15476 8968
rect 15528 8916 15534 8968
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 16408 8928 18245 8956
rect 1854 8888 1860 8900
rect 1815 8860 1860 8888
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 3510 8888 3516 8900
rect 3082 8860 3516 8888
rect 3510 8848 3516 8860
rect 3568 8848 3574 8900
rect 4798 8848 4804 8900
rect 4856 8848 4862 8900
rect 7101 8891 7159 8897
rect 7101 8857 7113 8891
rect 7147 8857 7159 8891
rect 10410 8888 10416 8900
rect 7101 8851 7159 8857
rect 8404 8860 10416 8888
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 6086 8820 6092 8832
rect 3200 8792 6092 8820
rect 3200 8780 3206 8792
rect 6086 8780 6092 8792
rect 6144 8780 6150 8832
rect 7116 8820 7144 8851
rect 8404 8820 8432 8860
rect 10410 8848 10416 8860
rect 10468 8848 10474 8900
rect 11330 8848 11336 8900
rect 11388 8848 11394 8900
rect 14274 8848 14280 8900
rect 14332 8888 14338 8900
rect 16408 8888 16436 8928
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 20990 8916 20996 8968
rect 21048 8956 21054 8968
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 21048 8928 21097 8956
rect 21048 8916 21054 8928
rect 21085 8925 21097 8928
rect 21131 8925 21143 8959
rect 21085 8919 21143 8925
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8956 24915 8959
rect 28442 8956 28448 8968
rect 24903 8928 28448 8956
rect 24903 8925 24915 8928
rect 24857 8919 24915 8925
rect 28442 8916 28448 8928
rect 28500 8916 28506 8968
rect 38010 8956 38016 8968
rect 37971 8928 38016 8956
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 14332 8860 16436 8888
rect 21177 8891 21235 8897
rect 14332 8848 14338 8860
rect 21177 8857 21189 8891
rect 21223 8888 21235 8891
rect 21913 8891 21971 8897
rect 21913 8888 21925 8891
rect 21223 8860 21925 8888
rect 21223 8857 21235 8860
rect 21177 8851 21235 8857
rect 21913 8857 21925 8860
rect 21959 8857 21971 8891
rect 21913 8851 21971 8857
rect 8570 8820 8576 8832
rect 7116 8792 8432 8820
rect 8531 8792 8576 8820
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 9582 8820 9588 8832
rect 8812 8792 9588 8820
rect 8812 8780 8818 8792
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 13538 8820 13544 8832
rect 9916 8792 13544 8820
rect 9916 8780 9922 8792
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 13814 8820 13820 8832
rect 13771 8792 13820 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 15473 8823 15531 8829
rect 15473 8789 15485 8823
rect 15519 8820 15531 8823
rect 16666 8820 16672 8832
rect 15519 8792 16672 8820
rect 15519 8789 15531 8792
rect 15473 8783 15531 8789
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 17405 8823 17463 8829
rect 17405 8820 17417 8823
rect 17368 8792 17417 8820
rect 17368 8780 17374 8792
rect 17405 8789 17417 8792
rect 17451 8789 17463 8823
rect 17405 8783 17463 8789
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 20346 8820 20352 8832
rect 18012 8792 20352 8820
rect 18012 8780 18018 8792
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 2240 8588 3832 8616
rect 2240 8557 2268 8588
rect 2225 8551 2283 8557
rect 2225 8517 2237 8551
rect 2271 8517 2283 8551
rect 2225 8511 2283 8517
rect 3326 8440 3332 8492
rect 3384 8440 3390 8492
rect 3804 8480 3832 8588
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 3936 8588 6040 8616
rect 3936 8576 3942 8588
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 5261 8551 5319 8557
rect 5261 8548 5273 8551
rect 5040 8520 5273 8548
rect 5040 8508 5046 8520
rect 5261 8517 5273 8520
rect 5307 8548 5319 8551
rect 5902 8548 5908 8560
rect 5307 8520 5908 8548
rect 5307 8517 5319 8520
rect 5261 8511 5319 8517
rect 5902 8508 5908 8520
rect 5960 8508 5966 8560
rect 4433 8483 4491 8489
rect 3804 8452 4108 8480
rect 1578 8372 1584 8424
rect 1636 8412 1642 8424
rect 1949 8415 2007 8421
rect 1949 8412 1961 8415
rect 1636 8384 1961 8412
rect 1636 8372 1642 8384
rect 1949 8381 1961 8384
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 2866 8372 2872 8424
rect 2924 8412 2930 8424
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 2924 8384 3985 8412
rect 2924 8372 2930 8384
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 4080 8412 4108 8452
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4614 8480 4620 8492
rect 4479 8452 4620 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 6012 8489 6040 8588
rect 6086 8576 6092 8628
rect 6144 8616 6150 8628
rect 8757 8619 8815 8625
rect 6144 8588 8616 8616
rect 6144 8576 6150 8588
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5997 8483 6055 8489
rect 5215 8452 5856 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 4080 8384 5764 8412
rect 3973 8375 4031 8381
rect 3694 8236 3700 8288
rect 3752 8276 3758 8288
rect 4617 8279 4675 8285
rect 4617 8276 4629 8279
rect 3752 8248 4629 8276
rect 3752 8236 3758 8248
rect 4617 8245 4629 8248
rect 4663 8245 4675 8279
rect 5736 8276 5764 8384
rect 5828 8353 5856 8452
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 6788 8384 7021 8412
rect 6788 8372 6794 8384
rect 7009 8381 7021 8384
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 8588 8412 8616 8588
rect 8757 8585 8769 8619
rect 8803 8616 8815 8619
rect 10134 8616 10140 8628
rect 8803 8588 10140 8616
rect 8803 8585 8815 8588
rect 8757 8579 8815 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10560 8588 10977 8616
rect 10560 8576 10566 8588
rect 10965 8585 10977 8588
rect 11011 8616 11023 8619
rect 15010 8616 15016 8628
rect 11011 8588 14504 8616
rect 14971 8588 15016 8616
rect 11011 8585 11023 8588
rect 10965 8579 11023 8585
rect 9766 8548 9772 8560
rect 9232 8520 9772 8548
rect 9030 8440 9036 8492
rect 9088 8480 9094 8492
rect 9232 8489 9260 8520
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 10042 8508 10048 8560
rect 10100 8508 10106 8560
rect 12250 8548 12256 8560
rect 11723 8520 12256 8548
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 9088 8452 9229 8480
rect 9088 8440 9094 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 11723 8480 11751 8520
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 13722 8548 13728 8560
rect 13202 8520 13728 8548
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 14476 8489 14504 8588
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 18230 8616 18236 8628
rect 15856 8588 18236 8616
rect 15758 8551 15816 8557
rect 15758 8517 15770 8551
rect 15804 8548 15816 8551
rect 15856 8548 15884 8588
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 24854 8616 24860 8628
rect 19306 8588 24860 8616
rect 17310 8548 17316 8560
rect 15804 8520 15884 8548
rect 17271 8520 17316 8548
rect 15804 8517 15816 8520
rect 15758 8511 15816 8517
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 17402 8508 17408 8560
rect 17460 8548 17466 8560
rect 18506 8548 18512 8560
rect 17460 8520 17505 8548
rect 18467 8520 18512 8548
rect 17460 8508 17466 8520
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 9217 8443 9275 8449
rect 10888 8452 11751 8480
rect 14461 8483 14519 8489
rect 10888 8412 10916 8452
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14921 8483 14979 8489
rect 14921 8480 14933 8483
rect 14507 8452 14933 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 14921 8449 14933 8452
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 18414 8440 18420 8492
rect 18472 8480 18478 8492
rect 18472 8452 18517 8480
rect 18472 8440 18478 8452
rect 7331 8384 8524 8412
rect 8588 8384 10916 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 5813 8347 5871 8353
rect 5813 8313 5825 8347
rect 5859 8313 5871 8347
rect 5994 8344 6000 8356
rect 5813 8307 5871 8313
rect 5920 8316 6000 8344
rect 5920 8276 5948 8316
rect 5994 8304 6000 8316
rect 6052 8304 6058 8356
rect 8496 8344 8524 8384
rect 10962 8372 10968 8424
rect 11020 8412 11026 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 11020 8384 11713 8412
rect 11020 8372 11026 8384
rect 11701 8381 11713 8384
rect 11747 8381 11759 8415
rect 11974 8412 11980 8424
rect 11935 8384 11980 8412
rect 11701 8375 11759 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 13446 8412 13452 8424
rect 13407 8384 13452 8412
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 15657 8415 15715 8421
rect 13596 8384 14412 8412
rect 13596 8372 13602 8384
rect 9214 8344 9220 8356
rect 8496 8316 9220 8344
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 14274 8344 14280 8356
rect 14235 8316 14280 8344
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 14384 8344 14412 8384
rect 15657 8381 15669 8415
rect 15703 8412 15715 8415
rect 15746 8412 15752 8424
rect 15703 8384 15752 8412
rect 15703 8381 15715 8384
rect 15657 8375 15715 8381
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8412 15991 8415
rect 16390 8412 16396 8424
rect 15979 8384 16396 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 15948 8344 15976 8375
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 17589 8415 17647 8421
rect 17589 8381 17601 8415
rect 17635 8412 17647 8415
rect 19306 8412 19334 8588
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 20070 8480 20076 8492
rect 20031 8452 20076 8480
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8480 20591 8483
rect 22002 8480 22008 8492
rect 20579 8452 22008 8480
rect 20579 8449 20591 8452
rect 20533 8443 20591 8449
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 28258 8480 28264 8492
rect 28219 8452 28264 8480
rect 28258 8440 28264 8452
rect 28316 8440 28322 8492
rect 20714 8412 20720 8424
rect 17635 8384 19334 8412
rect 20675 8384 20720 8412
rect 17635 8381 17647 8384
rect 17589 8375 17647 8381
rect 14384 8316 15976 8344
rect 16022 8304 16028 8356
rect 16080 8344 16086 8356
rect 17604 8344 17632 8375
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 16080 8316 17632 8344
rect 16080 8304 16086 8316
rect 18046 8304 18052 8356
rect 18104 8344 18110 8356
rect 21082 8344 21088 8356
rect 18104 8316 21088 8344
rect 18104 8304 18110 8316
rect 21082 8304 21088 8316
rect 21140 8304 21146 8356
rect 21177 8347 21235 8353
rect 21177 8313 21189 8347
rect 21223 8344 21235 8347
rect 22094 8344 22100 8356
rect 21223 8316 22100 8344
rect 21223 8313 21235 8316
rect 21177 8307 21235 8313
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 28353 8347 28411 8353
rect 28353 8313 28365 8347
rect 28399 8344 28411 8347
rect 30006 8344 30012 8356
rect 28399 8316 30012 8344
rect 28399 8313 28411 8316
rect 28353 8307 28411 8313
rect 30006 8304 30012 8316
rect 30064 8304 30070 8356
rect 5736 8248 5948 8276
rect 4617 8239 4675 8245
rect 9306 8236 9312 8288
rect 9364 8276 9370 8288
rect 9474 8279 9532 8285
rect 9474 8276 9486 8279
rect 9364 8248 9486 8276
rect 9364 8236 9370 8248
rect 9474 8245 9486 8248
rect 9520 8245 9532 8279
rect 9474 8239 9532 8245
rect 9582 8236 9588 8288
rect 9640 8276 9646 8288
rect 10134 8276 10140 8288
rect 9640 8248 10140 8276
rect 9640 8236 9646 8248
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 12434 8276 12440 8288
rect 11112 8248 12440 8276
rect 11112 8236 11118 8248
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 12526 8236 12532 8288
rect 12584 8276 12590 8288
rect 13998 8276 14004 8288
rect 12584 8248 14004 8276
rect 12584 8236 12590 8248
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 16114 8236 16120 8288
rect 16172 8276 16178 8288
rect 18874 8276 18880 8288
rect 16172 8248 18880 8276
rect 16172 8236 16178 8248
rect 18874 8236 18880 8248
rect 18932 8236 18938 8288
rect 19889 8279 19947 8285
rect 19889 8245 19901 8279
rect 19935 8276 19947 8279
rect 20622 8276 20628 8288
rect 19935 8248 20628 8276
rect 19935 8245 19947 8248
rect 19889 8239 19947 8245
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 2590 8072 2596 8084
rect 1912 8044 2596 8072
rect 1912 8032 1918 8044
rect 2590 8032 2596 8044
rect 2648 8072 2654 8084
rect 4617 8075 4675 8081
rect 2648 8044 4568 8072
rect 2648 8032 2654 8044
rect 3786 7964 3792 8016
rect 3844 8004 3850 8016
rect 4065 8007 4123 8013
rect 4065 8004 4077 8007
rect 3844 7976 4077 8004
rect 3844 7964 3850 7976
rect 4065 7973 4077 7976
rect 4111 7973 4123 8007
rect 4540 8004 4568 8044
rect 4617 8041 4629 8075
rect 4663 8072 4675 8075
rect 5166 8072 5172 8084
rect 4663 8044 5172 8072
rect 4663 8041 4675 8044
rect 4617 8035 4675 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 11054 8072 11060 8084
rect 5276 8044 11060 8072
rect 5276 8004 5304 8044
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 12437 8075 12495 8081
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 12710 8072 12716 8084
rect 12483 8044 12716 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 17126 8072 17132 8084
rect 15703 8044 17132 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 17402 8072 17408 8084
rect 17363 8044 17408 8072
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 19426 8072 19432 8084
rect 17552 8044 19432 8072
rect 17552 8032 17558 8044
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 20441 8075 20499 8081
rect 20441 8041 20453 8075
rect 20487 8072 20499 8075
rect 20714 8072 20720 8084
rect 20487 8044 20720 8072
rect 20487 8041 20499 8044
rect 20441 8035 20499 8041
rect 20714 8032 20720 8044
rect 20772 8032 20778 8084
rect 7282 8004 7288 8016
rect 4540 7976 5304 8004
rect 7243 7976 7288 8004
rect 4065 7967 4123 7973
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 9493 8007 9551 8013
rect 8220 7976 9444 8004
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 1903 7908 3556 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 3528 7868 3556 7908
rect 3602 7896 3608 7948
rect 3660 7936 3666 7948
rect 3660 7908 4844 7936
rect 3660 7896 3666 7908
rect 3878 7868 3884 7880
rect 3528 7840 3884 7868
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 4816 7877 4844 7908
rect 6454 7896 6460 7948
rect 6512 7936 6518 7948
rect 8220 7936 8248 7976
rect 6512 7908 8248 7936
rect 6512 7896 6518 7908
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 9306 7936 9312 7948
rect 8352 7908 9312 7936
rect 8352 7896 8358 7908
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 9416 7936 9444 7976
rect 9493 7973 9505 8007
rect 9539 8004 9551 8007
rect 9539 7976 10180 8004
rect 9539 7973 9551 7976
rect 9493 7967 9551 7973
rect 9416 7908 9720 7936
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4801 7871 4859 7877
rect 4019 7840 4752 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4062 7800 4068 7812
rect 3082 7772 4068 7800
rect 4062 7760 4068 7772
rect 4120 7760 4126 7812
rect 4724 7800 4752 7840
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5040 7840 5549 7868
rect 5040 7828 5046 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 8312 7868 8340 7896
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8312 7840 8401 7868
rect 5537 7831 5595 7837
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9272 7840 9413 7868
rect 9272 7828 9278 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9692 7868 9720 7908
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 9824 7908 10057 7936
rect 9824 7896 9830 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 10152 7936 10180 7976
rect 11422 7964 11428 8016
rect 11480 8004 11486 8016
rect 11480 7976 18276 8004
rect 11480 7964 11486 7976
rect 12066 7936 12072 7948
rect 10152 7908 12072 7936
rect 10045 7899 10103 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 12768 7908 14473 7936
rect 12768 7896 12774 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 16298 7936 16304 7948
rect 16259 7908 16304 7936
rect 14461 7899 14519 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 16448 7908 17632 7936
rect 16448 7896 16454 7908
rect 9950 7868 9956 7880
rect 9692 7840 9956 7868
rect 9401 7831 9459 7837
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 11422 7828 11428 7880
rect 11480 7828 11486 7880
rect 11698 7828 11704 7880
rect 11756 7868 11762 7880
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 11756 7840 12357 7868
rect 11756 7828 11762 7840
rect 12345 7837 12357 7840
rect 12391 7837 12403 7871
rect 12345 7831 12403 7837
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 13081 7871 13139 7877
rect 12492 7840 13032 7868
rect 12492 7828 12498 7840
rect 5350 7800 5356 7812
rect 4724 7772 5356 7800
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 5718 7760 5724 7812
rect 5776 7800 5782 7812
rect 5813 7803 5871 7809
rect 5813 7800 5825 7803
rect 5776 7772 5825 7800
rect 5776 7760 5782 7772
rect 5813 7769 5825 7772
rect 5859 7769 5871 7803
rect 8294 7800 8300 7812
rect 7038 7772 8300 7800
rect 5813 7763 5871 7769
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 8481 7803 8539 7809
rect 8481 7769 8493 7803
rect 8527 7800 8539 7803
rect 10226 7800 10232 7812
rect 8527 7772 10232 7800
rect 8527 7769 8539 7772
rect 8481 7763 8539 7769
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 10318 7760 10324 7812
rect 10376 7800 10382 7812
rect 12710 7800 12716 7812
rect 10376 7772 10421 7800
rect 11723 7772 12716 7800
rect 10376 7760 10382 7772
rect 3326 7732 3332 7744
rect 3239 7704 3332 7732
rect 3326 7692 3332 7704
rect 3384 7732 3390 7744
rect 8202 7732 8208 7744
rect 3384 7704 8208 7732
rect 3384 7692 3390 7704
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8570 7692 8576 7744
rect 8628 7732 8634 7744
rect 9030 7732 9036 7744
rect 8628 7704 9036 7732
rect 8628 7692 8634 7704
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 11723 7732 11751 7772
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 9364 7704 11751 7732
rect 11793 7735 11851 7741
rect 9364 7692 9370 7704
rect 11793 7701 11805 7735
rect 11839 7732 11851 7735
rect 12066 7732 12072 7744
rect 11839 7704 12072 7732
rect 11839 7701 11851 7704
rect 11793 7695 11851 7701
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 13004 7732 13032 7840
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13096 7800 13124 7831
rect 13170 7828 13176 7880
rect 13228 7868 13234 7880
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 13228 7840 13277 7868
rect 13228 7828 13234 7840
rect 13265 7837 13277 7840
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13872 7840 14289 7868
rect 13872 7828 13878 7840
rect 14277 7837 14289 7840
rect 14323 7868 14335 7871
rect 15010 7868 15016 7880
rect 14323 7840 15016 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7868 16543 7871
rect 16942 7868 16948 7880
rect 16531 7840 16948 7868
rect 16531 7837 16543 7840
rect 16485 7831 16543 7837
rect 15654 7800 15660 7812
rect 13096 7772 15660 7800
rect 15654 7760 15660 7772
rect 15712 7760 15718 7812
rect 15856 7800 15884 7831
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17604 7877 17632 7908
rect 18248 7877 18276 7976
rect 18322 7964 18328 8016
rect 18380 8004 18386 8016
rect 27801 8007 27859 8013
rect 27801 8004 27813 8007
rect 18380 7976 27813 8004
rect 18380 7964 18386 7976
rect 27801 7973 27813 7976
rect 27847 7973 27859 8007
rect 27801 7967 27859 7973
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7837 17647 7871
rect 17589 7831 17647 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 20622 7868 20628 7880
rect 20583 7840 20628 7868
rect 18693 7831 18751 7837
rect 17494 7800 17500 7812
rect 15856 7772 17500 7800
rect 17494 7760 17500 7772
rect 17552 7760 17558 7812
rect 17678 7760 17684 7812
rect 17736 7800 17742 7812
rect 18708 7800 18736 7831
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 21913 7871 21971 7877
rect 21913 7868 21925 7871
rect 20864 7840 21925 7868
rect 20864 7828 20870 7840
rect 21913 7837 21925 7840
rect 21959 7868 21971 7871
rect 22741 7871 22799 7877
rect 22741 7868 22753 7871
rect 21959 7840 22753 7868
rect 21959 7837 21971 7840
rect 21913 7831 21971 7837
rect 22741 7837 22753 7840
rect 22787 7837 22799 7871
rect 22741 7831 22799 7837
rect 27709 7871 27767 7877
rect 27709 7837 27721 7871
rect 27755 7868 27767 7871
rect 30190 7868 30196 7880
rect 27755 7840 30196 7868
rect 27755 7837 27767 7840
rect 27709 7831 27767 7837
rect 30190 7828 30196 7840
rect 30248 7828 30254 7880
rect 17736 7772 18736 7800
rect 17736 7760 17742 7772
rect 20530 7760 20536 7812
rect 20588 7800 20594 7812
rect 22462 7800 22468 7812
rect 20588 7772 22468 7800
rect 20588 7760 20594 7772
rect 22462 7760 22468 7772
rect 22520 7760 22526 7812
rect 13630 7732 13636 7744
rect 13004 7704 13636 7732
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7732 13783 7735
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 13771 7704 14933 7732
rect 13771 7701 13783 7704
rect 13725 7695 13783 7701
rect 14921 7701 14933 7704
rect 14967 7732 14979 7735
rect 16574 7732 16580 7744
rect 14967 7704 16580 7732
rect 14967 7701 14979 7704
rect 14921 7695 14979 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 16945 7735 17003 7741
rect 16945 7732 16957 7735
rect 16908 7704 16957 7732
rect 16908 7692 16914 7704
rect 16945 7701 16957 7704
rect 16991 7701 17003 7735
rect 16945 7695 17003 7701
rect 17586 7692 17592 7744
rect 17644 7732 17650 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 17644 7704 18061 7732
rect 17644 7692 17650 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 18049 7695 18107 7701
rect 18322 7692 18328 7744
rect 18380 7732 18386 7744
rect 18785 7735 18843 7741
rect 18785 7732 18797 7735
rect 18380 7704 18797 7732
rect 18380 7692 18386 7704
rect 18785 7701 18797 7704
rect 18831 7701 18843 7735
rect 18785 7695 18843 7701
rect 22005 7735 22063 7741
rect 22005 7701 22017 7735
rect 22051 7732 22063 7735
rect 22186 7732 22192 7744
rect 22051 7704 22192 7732
rect 22051 7701 22063 7704
rect 22005 7695 22063 7701
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 22557 7735 22615 7741
rect 22557 7701 22569 7735
rect 22603 7732 22615 7735
rect 22646 7732 22652 7744
rect 22603 7704 22652 7732
rect 22603 7701 22615 7704
rect 22557 7695 22615 7701
rect 22646 7692 22652 7704
rect 22704 7692 22710 7744
rect 23201 7735 23259 7741
rect 23201 7701 23213 7735
rect 23247 7732 23259 7735
rect 23290 7732 23296 7744
rect 23247 7704 23296 7732
rect 23247 7701 23259 7704
rect 23201 7695 23259 7701
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 6546 7528 6552 7540
rect 4632 7500 6552 7528
rect 1854 7460 1860 7472
rect 1815 7432 1860 7460
rect 1854 7420 1860 7432
rect 1912 7420 1918 7472
rect 4632 7460 4660 7500
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6914 7528 6920 7540
rect 6687 7500 6920 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 8846 7528 8852 7540
rect 7852 7500 8852 7528
rect 3082 7432 4660 7460
rect 5997 7463 6055 7469
rect 5997 7429 6009 7463
rect 6043 7460 6055 7463
rect 7742 7460 7748 7472
rect 6043 7432 7748 7460
rect 6043 7429 6055 7432
rect 5997 7423 6055 7429
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 5350 7352 5356 7404
rect 5408 7352 5414 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5460 7364 6561 7392
rect 5460 7336 5488 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 7469 7395 7527 7401
rect 7469 7361 7481 7395
rect 7515 7392 7527 7395
rect 7852 7392 7880 7500
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9030 7488 9036 7540
rect 9088 7528 9094 7540
rect 10594 7528 10600 7540
rect 9088 7500 10600 7528
rect 9088 7488 9094 7500
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 11149 7531 11207 7537
rect 11149 7497 11161 7531
rect 11195 7528 11207 7531
rect 12986 7528 12992 7540
rect 11195 7500 12992 7528
rect 11195 7497 11207 7500
rect 11149 7491 11207 7497
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 16025 7531 16083 7537
rect 13504 7500 15332 7528
rect 13504 7488 13510 7500
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 8205 7463 8263 7469
rect 8205 7460 8217 7463
rect 8168 7432 8217 7460
rect 8168 7420 8174 7432
rect 8205 7429 8217 7432
rect 8251 7429 8263 7463
rect 11054 7460 11060 7472
rect 9430 7432 11060 7460
rect 8205 7423 8263 7429
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 11974 7460 11980 7472
rect 11935 7432 11980 7460
rect 11974 7420 11980 7432
rect 12032 7420 12038 7472
rect 13998 7460 14004 7472
rect 13202 7432 14004 7460
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 14093 7463 14151 7469
rect 14093 7429 14105 7463
rect 14139 7460 14151 7463
rect 15194 7460 15200 7472
rect 14139 7432 15200 7460
rect 14139 7429 14151 7432
rect 14093 7423 14151 7429
rect 15194 7420 15200 7432
rect 15252 7420 15258 7472
rect 15304 7460 15332 7500
rect 16025 7497 16037 7531
rect 16071 7528 16083 7531
rect 16206 7528 16212 7540
rect 16071 7500 16212 7528
rect 16071 7497 16083 7500
rect 16025 7491 16083 7497
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 16942 7528 16948 7540
rect 16903 7500 16948 7528
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17034 7488 17040 7540
rect 17092 7528 17098 7540
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 17092 7500 17509 7528
rect 17092 7488 17098 7500
rect 17497 7497 17509 7500
rect 17543 7497 17555 7531
rect 18230 7528 18236 7540
rect 18191 7500 18236 7528
rect 17497 7491 17555 7497
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 18874 7528 18880 7540
rect 18835 7500 18880 7528
rect 18874 7488 18880 7500
rect 18932 7488 18938 7540
rect 29546 7528 29552 7540
rect 29507 7500 29552 7528
rect 29546 7488 29552 7500
rect 29604 7488 29610 7540
rect 33870 7528 33876 7540
rect 33831 7500 33876 7528
rect 33870 7488 33876 7500
rect 33928 7488 33934 7540
rect 36906 7488 36912 7540
rect 36964 7528 36970 7540
rect 38105 7531 38163 7537
rect 38105 7528 38117 7531
rect 36964 7500 38117 7528
rect 36964 7488 36970 7500
rect 38105 7497 38117 7500
rect 38151 7497 38163 7531
rect 38105 7491 38163 7497
rect 18322 7460 18328 7472
rect 15304 7432 18328 7460
rect 18322 7420 18328 7432
rect 18380 7420 18386 7472
rect 18598 7420 18604 7472
rect 18656 7460 18662 7472
rect 20990 7460 20996 7472
rect 18656 7432 20996 7460
rect 18656 7420 18662 7432
rect 20990 7420 20996 7432
rect 21048 7420 21054 7472
rect 22186 7460 22192 7472
rect 22147 7432 22192 7460
rect 22186 7420 22192 7432
rect 22244 7420 22250 7472
rect 23290 7460 23296 7472
rect 23251 7432 23296 7460
rect 23290 7420 23296 7432
rect 23348 7420 23354 7472
rect 23382 7420 23388 7472
rect 23440 7460 23446 7472
rect 23440 7432 23485 7460
rect 23440 7420 23446 7432
rect 9950 7392 9956 7404
rect 7515 7364 7880 7392
rect 9911 7364 9956 7392
rect 7515 7361 7527 7364
rect 7469 7355 7527 7361
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 10962 7392 10968 7404
rect 10376 7364 10968 7392
rect 10376 7352 10382 7364
rect 10962 7352 10968 7364
rect 11020 7392 11026 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11020 7364 11713 7392
rect 11020 7352 11026 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7392 14703 7395
rect 14918 7392 14924 7404
rect 14691 7364 14924 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7392 15347 7395
rect 15838 7392 15844 7404
rect 15335 7364 15844 7392
rect 15335 7361 15347 7364
rect 15289 7355 15347 7361
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7361 16267 7395
rect 16209 7355 16267 7361
rect 1578 7324 1584 7336
rect 1539 7296 1584 7324
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 3878 7284 3884 7336
rect 3936 7324 3942 7336
rect 3973 7327 4031 7333
rect 3973 7324 3985 7327
rect 3936 7296 3985 7324
rect 3936 7284 3942 7296
rect 3973 7293 3985 7296
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 4614 7324 4620 7336
rect 4295 7296 4620 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 5442 7284 5448 7336
rect 5500 7284 5506 7336
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 7929 7327 7987 7333
rect 7929 7324 7941 7327
rect 6788 7296 7941 7324
rect 6788 7284 6794 7296
rect 7929 7293 7941 7296
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 10502 7324 10508 7336
rect 8260 7296 9260 7324
rect 10463 7296 10508 7324
rect 8260 7284 8266 7296
rect 7282 7256 7288 7268
rect 7243 7228 7288 7256
rect 7282 7216 7288 7228
rect 7340 7216 7346 7268
rect 9232 7256 9260 7296
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7324 10747 7327
rect 13446 7324 13452 7336
rect 10735 7296 11836 7324
rect 10735 7293 10747 7296
rect 10689 7287 10747 7293
rect 11146 7256 11152 7268
rect 9232 7228 11152 7256
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 8938 7188 8944 7200
rect 3375 7160 8944 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 8938 7148 8944 7160
rect 8996 7188 9002 7200
rect 11698 7188 11704 7200
rect 8996 7160 11704 7188
rect 8996 7148 9002 7160
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 11808 7188 11836 7296
rect 13096 7296 13452 7324
rect 13096 7188 13124 7296
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 16224 7324 16252 7355
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16816 7364 16865 7392
rect 16816 7352 16822 7364
rect 16853 7361 16865 7364
rect 16899 7392 16911 7395
rect 17681 7395 17739 7401
rect 17681 7392 17693 7395
rect 16899 7364 17693 7392
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 17681 7361 17693 7364
rect 17727 7361 17739 7395
rect 17681 7355 17739 7361
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 17920 7364 18153 7392
rect 17920 7352 17926 7364
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7361 18843 7395
rect 18785 7355 18843 7361
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7392 19487 7395
rect 19886 7392 19892 7404
rect 19475 7364 19892 7392
rect 19475 7361 19487 7364
rect 19429 7355 19487 7361
rect 17034 7324 17040 7336
rect 14047 7296 15148 7324
rect 16224 7296 17040 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 15120 7265 15148 7296
rect 17034 7284 17040 7296
rect 17092 7284 17098 7336
rect 18800 7324 18828 7355
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 20070 7352 20076 7404
rect 20128 7392 20134 7404
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 20128 7364 20545 7392
rect 20128 7352 20134 7364
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 29457 7395 29515 7401
rect 29457 7361 29469 7395
rect 29503 7392 29515 7395
rect 33781 7395 33839 7401
rect 29503 7364 31754 7392
rect 29503 7361 29515 7364
rect 29457 7355 29515 7361
rect 19334 7324 19340 7336
rect 18800 7296 19340 7324
rect 19334 7284 19340 7296
rect 19392 7284 19398 7336
rect 22094 7284 22100 7336
rect 22152 7324 22158 7336
rect 22741 7327 22799 7333
rect 22152 7296 22197 7324
rect 22152 7284 22158 7296
rect 22741 7293 22753 7327
rect 22787 7324 22799 7327
rect 23937 7327 23995 7333
rect 23937 7324 23949 7327
rect 22787 7296 23949 7324
rect 22787 7293 22799 7296
rect 22741 7287 22799 7293
rect 23937 7293 23949 7296
rect 23983 7324 23995 7327
rect 29546 7324 29552 7336
rect 23983 7296 29552 7324
rect 23983 7293 23995 7296
rect 23937 7287 23995 7293
rect 29546 7284 29552 7296
rect 29604 7284 29610 7336
rect 31726 7324 31754 7364
rect 33781 7361 33793 7395
rect 33827 7392 33839 7395
rect 35710 7392 35716 7404
rect 33827 7364 35716 7392
rect 33827 7361 33839 7364
rect 33781 7355 33839 7361
rect 35710 7352 35716 7364
rect 35768 7352 35774 7404
rect 38286 7392 38292 7404
rect 38247 7364 38292 7392
rect 38286 7352 38292 7364
rect 38344 7352 38350 7404
rect 34698 7324 34704 7336
rect 31726 7296 34704 7324
rect 34698 7284 34704 7296
rect 34756 7284 34762 7336
rect 15105 7259 15163 7265
rect 15105 7225 15117 7259
rect 15151 7225 15163 7259
rect 15105 7219 15163 7225
rect 16482 7216 16488 7268
rect 16540 7256 16546 7268
rect 16942 7256 16948 7268
rect 16540 7228 16948 7256
rect 16540 7216 16546 7228
rect 16942 7216 16948 7228
rect 17000 7216 17006 7268
rect 17586 7216 17592 7268
rect 17644 7256 17650 7268
rect 19521 7259 19579 7265
rect 19521 7256 19533 7259
rect 17644 7228 19533 7256
rect 17644 7216 17650 7228
rect 19521 7225 19533 7228
rect 19567 7225 19579 7259
rect 19521 7219 19579 7225
rect 13446 7188 13452 7200
rect 11808 7160 13124 7188
rect 13407 7160 13452 7188
rect 13446 7148 13452 7160
rect 13504 7188 13510 7200
rect 17862 7188 17868 7200
rect 13504 7160 17868 7188
rect 13504 7148 13510 7160
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 20625 7191 20683 7197
rect 20625 7157 20637 7191
rect 20671 7188 20683 7191
rect 20990 7188 20996 7200
rect 20671 7160 20996 7188
rect 20671 7157 20683 7160
rect 20625 7151 20683 7157
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1936 6987 1994 6993
rect 1936 6953 1948 6987
rect 1982 6984 1994 6987
rect 3326 6984 3332 6996
rect 1982 6956 3332 6984
rect 1982 6953 1994 6956
rect 1936 6947 1994 6953
rect 3326 6944 3332 6956
rect 3384 6944 3390 6996
rect 4236 6987 4294 6993
rect 4236 6953 4248 6987
rect 4282 6984 4294 6987
rect 4614 6984 4620 6996
rect 4282 6956 4620 6984
rect 4282 6953 4294 6956
rect 4236 6947 4294 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 7088 6987 7146 6993
rect 7088 6953 7100 6987
rect 7134 6984 7146 6987
rect 7742 6984 7748 6996
rect 7134 6956 7748 6984
rect 7134 6953 7146 6956
rect 7088 6947 7146 6953
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 13446 6984 13452 6996
rect 10100 6956 13452 6984
rect 10100 6944 10106 6956
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 13630 6944 13636 6996
rect 13688 6984 13694 6996
rect 16206 6984 16212 6996
rect 13688 6956 16212 6984
rect 13688 6944 13694 6956
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 17494 6944 17500 6996
rect 17552 6984 17558 6996
rect 17589 6987 17647 6993
rect 17589 6984 17601 6987
rect 17552 6956 17601 6984
rect 17552 6944 17558 6956
rect 17589 6953 17601 6956
rect 17635 6953 17647 6987
rect 17589 6947 17647 6953
rect 22465 6987 22523 6993
rect 22465 6953 22477 6987
rect 22511 6984 22523 6987
rect 23382 6984 23388 6996
rect 22511 6956 23388 6984
rect 22511 6953 22523 6956
rect 22465 6947 22523 6953
rect 23382 6944 23388 6956
rect 23440 6944 23446 6996
rect 9692 6888 10456 6916
rect 3878 6848 3884 6860
rect 1688 6820 3884 6848
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 1688 6789 1716 6820
rect 3878 6808 3884 6820
rect 3936 6848 3942 6860
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3936 6820 3985 6848
rect 3936 6808 3942 6820
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 6730 6848 6736 6860
rect 5040 6820 6736 6848
rect 5040 6808 5046 6820
rect 6730 6808 6736 6820
rect 6788 6848 6794 6860
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6788 6820 6837 6848
rect 6788 6808 6794 6820
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 9692 6848 9720 6888
rect 7156 6820 9720 6848
rect 7156 6808 7162 6820
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 10318 6848 10324 6860
rect 9824 6820 10324 6848
rect 9824 6808 9830 6820
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10428 6848 10456 6888
rect 12066 6876 12072 6928
rect 12124 6916 12130 6928
rect 14550 6916 14556 6928
rect 12124 6888 14556 6916
rect 12124 6876 12130 6888
rect 14550 6876 14556 6888
rect 14608 6876 14614 6928
rect 15856 6888 19334 6916
rect 11330 6848 11336 6860
rect 10428 6820 11336 6848
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 13170 6848 13176 6860
rect 11900 6820 13176 6848
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 1636 6752 1685 6780
rect 1636 6740 1642 6752
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 5718 6780 5724 6792
rect 5592 6752 5724 6780
rect 5592 6740 5598 6752
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 5994 6780 6000 6792
rect 5955 6752 6000 6780
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 9858 6780 9864 6792
rect 9819 6752 9864 6780
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 2222 6672 2228 6724
rect 2280 6712 2286 6724
rect 2280 6684 2438 6712
rect 2280 6672 2286 6684
rect 5258 6672 5264 6724
rect 5316 6672 5322 6724
rect 5552 6684 7420 6712
rect 2314 6604 2320 6656
rect 2372 6644 2378 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 2372 6616 3433 6644
rect 2372 6604 2378 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 5552 6644 5580 6684
rect 4212 6616 5580 6644
rect 4212 6604 4218 6616
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 7282 6644 7288 6656
rect 5776 6616 7288 6644
rect 5776 6604 5782 6616
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7392 6644 7420 6684
rect 7558 6672 7564 6724
rect 7616 6672 7622 6724
rect 10226 6712 10232 6724
rect 8404 6684 10232 6712
rect 7834 6644 7840 6656
rect 7392 6616 7840 6644
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 8404 6644 8432 6684
rect 10226 6672 10232 6684
rect 10284 6672 10290 6724
rect 10502 6672 10508 6724
rect 10560 6712 10566 6724
rect 10597 6715 10655 6721
rect 10597 6712 10609 6715
rect 10560 6684 10609 6712
rect 10560 6672 10566 6684
rect 10597 6681 10609 6684
rect 10643 6681 10655 6715
rect 10597 6675 10655 6681
rect 11146 6672 11152 6724
rect 11204 6672 11210 6724
rect 8570 6644 8576 6656
rect 8168 6616 8432 6644
rect 8531 6616 8576 6644
rect 8168 6604 8174 6616
rect 8570 6604 8576 6616
rect 8628 6644 8634 6656
rect 9490 6644 9496 6656
rect 8628 6616 9496 6644
rect 8628 6604 8634 6616
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 11900 6644 11928 6820
rect 13170 6808 13176 6820
rect 13228 6808 13234 6860
rect 13265 6851 13323 6857
rect 13265 6817 13277 6851
rect 13311 6848 13323 6851
rect 15378 6848 15384 6860
rect 13311 6820 15384 6848
rect 13311 6817 13323 6820
rect 13265 6811 13323 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 15856 6857 15884 6888
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6817 15899 6851
rect 15841 6811 15899 6817
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 17037 6851 17095 6857
rect 17037 6848 17049 6851
rect 16071 6820 17049 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 17037 6817 17049 6820
rect 17083 6817 17095 6851
rect 19306 6848 19334 6888
rect 19426 6876 19432 6928
rect 19484 6916 19490 6928
rect 20438 6916 20444 6928
rect 19484 6888 20444 6916
rect 19484 6876 19490 6888
rect 20438 6876 20444 6888
rect 20496 6876 20502 6928
rect 20824 6888 21128 6916
rect 20257 6851 20315 6857
rect 20257 6848 20269 6851
rect 19306 6820 20269 6848
rect 17037 6811 17095 6817
rect 20257 6817 20269 6820
rect 20303 6817 20315 6851
rect 20824 6848 20852 6888
rect 20990 6848 20996 6860
rect 20257 6811 20315 6817
rect 20732 6820 20852 6848
rect 20951 6820 20996 6848
rect 13078 6780 13084 6792
rect 13039 6752 13084 6780
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 14274 6740 14280 6792
rect 14332 6780 14338 6792
rect 14461 6783 14519 6789
rect 14332 6752 14377 6780
rect 14332 6740 14338 6752
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 16850 6780 16856 6792
rect 14507 6752 16856 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 17773 6783 17831 6789
rect 17000 6752 17045 6780
rect 17000 6740 17006 6752
rect 17773 6749 17785 6783
rect 17819 6780 17831 6783
rect 17862 6780 17868 6792
rect 17819 6752 17868 6780
rect 17819 6749 17831 6752
rect 17773 6743 17831 6749
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 18417 6783 18475 6789
rect 18417 6780 18429 6783
rect 18104 6752 18429 6780
rect 18104 6740 18110 6752
rect 18417 6749 18429 6752
rect 18463 6749 18475 6783
rect 18417 6743 18475 6749
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 18656 6752 19441 6780
rect 18656 6740 18662 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 19521 6783 19579 6789
rect 19521 6749 19533 6783
rect 19567 6780 19579 6783
rect 19978 6780 19984 6792
rect 19567 6752 19984 6780
rect 19567 6749 19579 6752
rect 19521 6743 19579 6749
rect 11974 6672 11980 6724
rect 12032 6712 12038 6724
rect 14366 6712 14372 6724
rect 12032 6684 14372 6712
rect 12032 6672 12038 6684
rect 14366 6672 14372 6684
rect 14424 6672 14430 6724
rect 19444 6712 19472 6743
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 20165 6783 20223 6789
rect 20165 6749 20177 6783
rect 20211 6780 20223 6783
rect 20732 6780 20760 6820
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 20211 6752 20760 6780
rect 20809 6783 20867 6789
rect 20211 6749 20223 6752
rect 20165 6743 20223 6749
rect 20809 6749 20821 6783
rect 20855 6749 20867 6783
rect 21100 6780 21128 6888
rect 21453 6851 21511 6857
rect 21453 6817 21465 6851
rect 21499 6848 21511 6851
rect 22094 6848 22100 6860
rect 21499 6820 22100 6848
rect 21499 6817 21511 6820
rect 21453 6811 21511 6817
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 24578 6848 24584 6860
rect 22480 6820 24584 6848
rect 22480 6780 22508 6820
rect 24578 6808 24584 6820
rect 24636 6808 24642 6860
rect 31941 6851 31999 6857
rect 31941 6848 31953 6851
rect 31726 6820 31953 6848
rect 22646 6780 22652 6792
rect 21100 6752 22508 6780
rect 22607 6752 22652 6780
rect 20809 6743 20867 6749
rect 20714 6712 20720 6724
rect 19444 6684 20720 6712
rect 20714 6672 20720 6684
rect 20772 6672 20778 6724
rect 20824 6712 20852 6743
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 31202 6712 31208 6724
rect 20824 6684 31208 6712
rect 31202 6672 31208 6684
rect 31260 6672 31266 6724
rect 12066 6644 12072 6656
rect 9723 6616 11928 6644
rect 12027 6616 12072 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 13078 6604 13084 6656
rect 13136 6644 13142 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 13136 6616 13737 6644
rect 13136 6604 13142 6616
rect 13725 6613 13737 6616
rect 13771 6644 13783 6647
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 13771 6616 14933 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 14921 6613 14933 6616
rect 14967 6613 14979 6647
rect 14921 6607 14979 6613
rect 15010 6604 15016 6656
rect 15068 6644 15074 6656
rect 16485 6647 16543 6653
rect 16485 6644 16497 6647
rect 15068 6616 16497 6644
rect 15068 6604 15074 6616
rect 16485 6613 16497 6616
rect 16531 6613 16543 6647
rect 16485 6607 16543 6613
rect 17034 6604 17040 6656
rect 17092 6644 17098 6656
rect 18233 6647 18291 6653
rect 18233 6644 18245 6647
rect 17092 6616 18245 6644
rect 17092 6604 17098 6616
rect 18233 6613 18245 6616
rect 18279 6613 18291 6647
rect 18233 6607 18291 6613
rect 21450 6604 21456 6656
rect 21508 6644 21514 6656
rect 31726 6644 31754 6820
rect 31941 6817 31953 6820
rect 31987 6817 31999 6851
rect 31941 6811 31999 6817
rect 31849 6783 31907 6789
rect 31849 6749 31861 6783
rect 31895 6780 31907 6783
rect 33870 6780 33876 6792
rect 31895 6752 33876 6780
rect 31895 6749 31907 6752
rect 31849 6743 31907 6749
rect 33870 6740 33876 6752
rect 33928 6740 33934 6792
rect 21508 6616 31754 6644
rect 21508 6604 21514 6616
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 2498 6400 2504 6452
rect 2556 6400 2562 6452
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 2740 6412 9720 6440
rect 2740 6400 2746 6412
rect 2516 6372 2544 6400
rect 4065 6375 4123 6381
rect 2516 6344 2806 6372
rect 4065 6341 4077 6375
rect 4111 6372 4123 6375
rect 4154 6372 4160 6384
rect 4111 6344 4160 6372
rect 4111 6341 4123 6344
rect 4065 6335 4123 6341
rect 4154 6332 4160 6344
rect 4212 6332 4218 6384
rect 4617 6375 4675 6381
rect 4617 6372 4629 6375
rect 4448 6344 4629 6372
rect 1578 6196 1584 6248
rect 1636 6236 1642 6248
rect 2041 6239 2099 6245
rect 2041 6236 2053 6239
rect 1636 6208 2053 6236
rect 1636 6196 1642 6208
rect 2041 6205 2053 6208
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 2774 6236 2780 6248
rect 2363 6208 2780 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 4448 6236 4476 6344
rect 4617 6341 4629 6344
rect 4663 6341 4675 6375
rect 7098 6372 7104 6384
rect 4617 6335 4675 6341
rect 5644 6344 7104 6372
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6304 4583 6307
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 4571 6276 5181 6304
rect 4571 6273 4583 6276
rect 4525 6267 4583 6273
rect 4632 6248 4660 6276
rect 5169 6273 5181 6276
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 5644 6304 5672 6344
rect 7098 6332 7104 6344
rect 7156 6332 7162 6384
rect 7282 6372 7288 6384
rect 7243 6344 7288 6372
rect 7282 6332 7288 6344
rect 7340 6332 7346 6384
rect 9692 6372 9720 6412
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 11974 6440 11980 6452
rect 9916 6412 11980 6440
rect 9916 6400 9922 6412
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 15657 6443 15715 6449
rect 15657 6440 15669 6443
rect 12768 6412 15669 6440
rect 12768 6400 12774 6412
rect 15657 6409 15669 6412
rect 15703 6409 15715 6443
rect 15657 6403 15715 6409
rect 16117 6443 16175 6449
rect 16117 6409 16129 6443
rect 16163 6440 16175 6443
rect 16390 6440 16396 6452
rect 16163 6412 16396 6440
rect 16163 6409 16175 6412
rect 16117 6403 16175 6409
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 18690 6400 18696 6452
rect 18748 6440 18754 6452
rect 18785 6443 18843 6449
rect 18785 6440 18797 6443
rect 18748 6412 18797 6440
rect 18748 6400 18754 6412
rect 18785 6409 18797 6412
rect 18831 6409 18843 6443
rect 18785 6403 18843 6409
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 19300 6412 19441 6440
rect 19300 6400 19306 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 20717 6443 20775 6449
rect 20717 6409 20729 6443
rect 20763 6440 20775 6443
rect 21634 6440 21640 6452
rect 20763 6412 21640 6440
rect 20763 6409 20775 6412
rect 20717 6403 20775 6409
rect 21634 6400 21640 6412
rect 21692 6400 21698 6452
rect 9692 6344 12466 6372
rect 13906 6332 13912 6384
rect 13964 6372 13970 6384
rect 14185 6375 14243 6381
rect 14185 6372 14197 6375
rect 13964 6344 14197 6372
rect 13964 6332 13970 6344
rect 14185 6341 14197 6344
rect 14231 6372 14243 6375
rect 14274 6372 14280 6384
rect 14231 6344 14280 6372
rect 14231 6341 14243 6344
rect 14185 6335 14243 6341
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 17034 6372 17040 6384
rect 16995 6344 17040 6372
rect 17034 6332 17040 6344
rect 17092 6332 17098 6384
rect 20070 6372 20076 6384
rect 20031 6344 20076 6372
rect 20070 6332 20076 6344
rect 20128 6332 20134 6384
rect 20456 6344 21312 6372
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5307 6276 5672 6304
rect 5736 6276 5825 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 4448 6208 4568 6236
rect 4540 6168 4568 6208
rect 4614 6196 4620 6248
rect 4672 6196 4678 6248
rect 5184 6236 5212 6267
rect 5442 6236 5448 6248
rect 5184 6208 5448 6236
rect 5442 6196 5448 6208
rect 5500 6236 5506 6248
rect 5736 6236 5764 6276
rect 5813 6273 5825 6276
rect 5859 6304 5871 6307
rect 6454 6304 6460 6316
rect 5859 6276 6460 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6454 6264 6460 6276
rect 6512 6304 6518 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6512 6276 6561 6304
rect 6512 6264 6518 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6549 6267 6607 6273
rect 6656 6276 7205 6304
rect 6656 6236 6684 6276
rect 7193 6273 7205 6276
rect 7239 6304 7251 6307
rect 8018 6304 8024 6316
rect 7239 6276 8024 6304
rect 7239 6273 7251 6276
rect 7193 6267 7251 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 11054 6304 11060 6316
rect 9522 6276 11060 6304
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 11422 6304 11428 6316
rect 11195 6276 11428 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11422 6264 11428 6276
rect 11480 6264 11486 6316
rect 15286 6264 15292 6316
rect 15344 6264 15350 6316
rect 16298 6304 16304 6316
rect 16259 6276 16304 6304
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 17678 6264 17684 6316
rect 17736 6304 17742 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 17736 6276 18245 6304
rect 17736 6264 17742 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 19334 6304 19340 6316
rect 18739 6276 19340 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 19334 6264 19340 6276
rect 19392 6264 19398 6316
rect 19978 6304 19984 6316
rect 19939 6276 19984 6304
rect 19978 6264 19984 6276
rect 20036 6304 20042 6316
rect 20456 6304 20484 6344
rect 20622 6304 20628 6316
rect 20036 6276 20484 6304
rect 20583 6276 20628 6304
rect 20036 6264 20042 6276
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 21284 6313 21312 6344
rect 21269 6307 21327 6313
rect 21269 6273 21281 6307
rect 21315 6273 21327 6307
rect 21269 6267 21327 6273
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6304 22339 6307
rect 24210 6304 24216 6316
rect 22327 6276 24216 6304
rect 22327 6273 22339 6276
rect 22281 6267 22339 6273
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 29546 6304 29552 6316
rect 29507 6276 29552 6304
rect 29546 6264 29552 6276
rect 29604 6264 29610 6316
rect 5500 6208 5764 6236
rect 5828 6208 6684 6236
rect 5500 6196 5506 6208
rect 5626 6168 5632 6180
rect 4540 6140 5632 6168
rect 5626 6128 5632 6140
rect 5684 6128 5690 6180
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 5828 6100 5856 6208
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 6788 6208 8125 6236
rect 6788 6196 6794 6208
rect 8113 6205 8125 6208
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 10042 6236 10048 6248
rect 8435 6208 10048 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 10137 6239 10195 6245
rect 10137 6205 10149 6239
rect 10183 6205 10195 6239
rect 10137 6199 10195 6205
rect 5905 6171 5963 6177
rect 5905 6137 5917 6171
rect 5951 6168 5963 6171
rect 10152 6168 10180 6199
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 10376 6208 11713 6236
rect 10376 6196 10382 6208
rect 11701 6205 11713 6208
rect 11747 6236 11759 6239
rect 11974 6236 11980 6248
rect 11747 6208 11836 6236
rect 11935 6208 11980 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 10870 6168 10876 6180
rect 5951 6140 8156 6168
rect 10152 6140 10876 6168
rect 5951 6137 5963 6140
rect 5905 6131 5963 6137
rect 2464 6072 5856 6100
rect 6641 6103 6699 6109
rect 2464 6060 2470 6072
rect 6641 6069 6653 6103
rect 6687 6100 6699 6103
rect 6822 6100 6828 6112
rect 6687 6072 6828 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 8128 6100 8156 6140
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 10965 6171 11023 6177
rect 10965 6137 10977 6171
rect 11011 6168 11023 6171
rect 11606 6168 11612 6180
rect 11011 6140 11612 6168
rect 11011 6137 11023 6140
rect 10965 6131 11023 6137
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 8754 6100 8760 6112
rect 8128 6072 8760 6100
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 11698 6100 11704 6112
rect 9456 6072 11704 6100
rect 9456 6060 9462 6072
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 11808 6100 11836 6208
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 13906 6236 13912 6248
rect 13004 6208 13912 6236
rect 13004 6100 13032 6208
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 16945 6239 17003 6245
rect 16945 6236 16957 6239
rect 16540 6208 16957 6236
rect 16540 6196 16546 6208
rect 16945 6205 16957 6208
rect 16991 6205 17003 6239
rect 17218 6236 17224 6248
rect 17179 6208 17224 6236
rect 16945 6199 17003 6205
rect 17218 6196 17224 6208
rect 17276 6196 17282 6248
rect 19150 6196 19156 6248
rect 19208 6236 19214 6248
rect 21450 6236 21456 6248
rect 19208 6208 21456 6236
rect 19208 6196 19214 6208
rect 21450 6196 21456 6208
rect 21508 6196 21514 6248
rect 13446 6168 13452 6180
rect 13407 6140 13452 6168
rect 13446 6128 13452 6140
rect 13504 6128 13510 6180
rect 15286 6128 15292 6180
rect 15344 6168 15350 6180
rect 21358 6168 21364 6180
rect 15344 6140 18184 6168
rect 21319 6140 21364 6168
rect 15344 6128 15350 6140
rect 11808 6072 13032 6100
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 16022 6100 16028 6112
rect 13872 6072 16028 6100
rect 13872 6060 13878 6072
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 18156 6100 18184 6140
rect 21358 6128 21364 6140
rect 21416 6128 21422 6180
rect 22373 6103 22431 6109
rect 22373 6100 22385 6103
rect 18156 6072 22385 6100
rect 22373 6069 22385 6072
rect 22419 6069 22431 6103
rect 29638 6100 29644 6112
rect 29599 6072 29644 6100
rect 22373 6063 22431 6069
rect 29638 6060 29644 6072
rect 29696 6060 29702 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1844 5899 1902 5905
rect 1844 5865 1856 5899
rect 1890 5896 1902 5899
rect 4062 5896 4068 5908
rect 1890 5868 4068 5896
rect 1890 5865 1902 5868
rect 1844 5859 1902 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 7653 5899 7711 5905
rect 7653 5896 7665 5899
rect 6604 5868 7665 5896
rect 6604 5856 6610 5868
rect 7653 5865 7665 5868
rect 7699 5865 7711 5899
rect 8570 5896 8576 5908
rect 7653 5859 7711 5865
rect 8128 5868 8576 5896
rect 2958 5788 2964 5840
rect 3016 5828 3022 5840
rect 3329 5831 3387 5837
rect 3329 5828 3341 5831
rect 3016 5800 3341 5828
rect 3016 5788 3022 5800
rect 3329 5797 3341 5800
rect 3375 5797 3387 5831
rect 8128 5828 8156 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9306 5896 9312 5908
rect 9267 5868 9312 5896
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 9953 5899 10011 5905
rect 9953 5896 9965 5899
rect 9640 5868 9965 5896
rect 9640 5856 9646 5868
rect 9953 5865 9965 5868
rect 9999 5865 10011 5899
rect 9953 5859 10011 5865
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 10962 5896 10968 5908
rect 10836 5868 10968 5896
rect 10836 5856 10842 5868
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 11882 5896 11888 5908
rect 11296 5868 11888 5896
rect 11296 5856 11302 5868
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 18509 5899 18567 5905
rect 18509 5896 18521 5899
rect 12124 5868 18521 5896
rect 12124 5856 12130 5868
rect 18509 5865 18521 5868
rect 18555 5865 18567 5899
rect 18509 5859 18567 5865
rect 19426 5856 19432 5908
rect 19484 5896 19490 5908
rect 19521 5899 19579 5905
rect 19521 5896 19533 5899
rect 19484 5868 19533 5896
rect 19484 5856 19490 5868
rect 19521 5865 19533 5868
rect 19567 5865 19579 5899
rect 19521 5859 19579 5865
rect 20809 5899 20867 5905
rect 20809 5865 20821 5899
rect 20855 5896 20867 5899
rect 20898 5896 20904 5908
rect 20855 5868 20904 5896
rect 20855 5865 20867 5868
rect 20809 5859 20867 5865
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 21266 5856 21272 5908
rect 21324 5896 21330 5908
rect 21453 5899 21511 5905
rect 21453 5896 21465 5899
rect 21324 5868 21465 5896
rect 21324 5856 21330 5868
rect 21453 5865 21465 5868
rect 21499 5865 21511 5899
rect 21453 5859 21511 5865
rect 22094 5856 22100 5908
rect 22152 5896 22158 5908
rect 22152 5868 22197 5896
rect 22152 5856 22158 5868
rect 18598 5828 18604 5840
rect 3329 5791 3387 5797
rect 6472 5800 8156 5828
rect 8220 5800 10640 5828
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5760 5411 5763
rect 6472 5760 6500 5800
rect 5399 5732 6500 5760
rect 5399 5729 5411 5732
rect 5353 5723 5411 5729
rect 6546 5720 6552 5772
rect 6604 5720 6610 5772
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 4062 5692 4068 5704
rect 2990 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4212 5664 4257 5692
rect 4212 5652 4218 5664
rect 4982 5652 4988 5704
rect 5040 5692 5046 5704
rect 5077 5695 5135 5701
rect 5077 5692 5089 5695
rect 5040 5664 5089 5692
rect 5040 5652 5046 5664
rect 5077 5661 5089 5664
rect 5123 5661 5135 5695
rect 6564 5692 6592 5720
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 6564 5664 7573 5692
rect 5077 5655 5135 5661
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8220 5701 8248 5800
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 8343 5732 9996 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 8076 5664 8217 5692
rect 8076 5652 8082 5664
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8478 5692 8484 5704
rect 8205 5655 8263 5661
rect 8312 5664 8484 5692
rect 6730 5624 6736 5636
rect 4264 5596 5580 5624
rect 6578 5596 6736 5624
rect 4062 5556 4068 5568
rect 3975 5528 4068 5556
rect 4062 5516 4068 5528
rect 4120 5556 4126 5568
rect 4264 5556 4292 5596
rect 5552 5568 5580 5596
rect 6730 5584 6736 5596
rect 6788 5584 6794 5636
rect 7101 5627 7159 5633
rect 7101 5593 7113 5627
rect 7147 5624 7159 5627
rect 7282 5624 7288 5636
rect 7147 5596 7288 5624
rect 7147 5593 7159 5596
rect 7101 5587 7159 5593
rect 7282 5584 7288 5596
rect 7340 5624 7346 5636
rect 8312 5624 8340 5664
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 9180 5664 9229 5692
rect 9180 5652 9186 5664
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 7340 5596 8340 5624
rect 7340 5584 7346 5596
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 9876 5624 9904 5655
rect 8444 5596 9904 5624
rect 9968 5624 9996 5732
rect 10318 5720 10324 5772
rect 10376 5760 10382 5772
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 10376 5732 10517 5760
rect 10376 5720 10382 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10612 5760 10640 5800
rect 11808 5800 14412 5828
rect 11808 5760 11836 5800
rect 10612 5732 11836 5760
rect 10505 5723 10563 5729
rect 12066 5720 12072 5772
rect 12124 5720 12130 5772
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 12400 5732 12541 5760
rect 12400 5720 12406 5732
rect 12529 5729 12541 5732
rect 12575 5729 12587 5763
rect 13078 5760 13084 5772
rect 13039 5732 13084 5760
rect 12529 5723 12587 5729
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 13725 5763 13783 5769
rect 13725 5729 13737 5763
rect 13771 5760 13783 5763
rect 13814 5760 13820 5772
rect 13771 5732 13820 5760
rect 13771 5729 13783 5732
rect 13725 5723 13783 5729
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 13906 5720 13912 5772
rect 13964 5760 13970 5772
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 13964 5732 14289 5760
rect 13964 5720 13970 5732
rect 14277 5729 14289 5732
rect 14323 5729 14335 5763
rect 14384 5760 14412 5800
rect 15580 5800 18604 5828
rect 15580 5760 15608 5800
rect 18598 5788 18604 5800
rect 18656 5788 18662 5840
rect 16022 5760 16028 5772
rect 14384 5732 15608 5760
rect 15983 5732 16028 5760
rect 14277 5723 14335 5729
rect 16022 5720 16028 5732
rect 16080 5720 16086 5772
rect 16482 5760 16488 5772
rect 16443 5732 16488 5760
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 17218 5720 17224 5772
rect 17276 5760 17282 5772
rect 23382 5760 23388 5772
rect 17276 5732 23388 5760
rect 17276 5720 17282 5732
rect 23382 5720 23388 5732
rect 23440 5720 23446 5772
rect 12084 5692 12112 5720
rect 11914 5664 12112 5692
rect 16298 5652 16304 5704
rect 16356 5692 16362 5704
rect 17129 5695 17187 5701
rect 17129 5692 17141 5695
rect 16356 5664 17141 5692
rect 16356 5652 16362 5664
rect 17129 5661 17141 5664
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5692 17831 5695
rect 17954 5692 17960 5704
rect 17819 5664 17960 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 17954 5652 17960 5664
rect 18012 5692 18018 5704
rect 18414 5692 18420 5704
rect 18012 5664 18420 5692
rect 18012 5652 18018 5664
rect 18414 5652 18420 5664
rect 18472 5652 18478 5704
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 19392 5664 19441 5692
rect 19392 5652 19398 5664
rect 19429 5661 19441 5664
rect 19475 5692 19487 5695
rect 19518 5692 19524 5704
rect 19475 5664 19524 5692
rect 19475 5661 19487 5664
rect 19429 5655 19487 5661
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 19978 5652 19984 5704
rect 20036 5692 20042 5704
rect 20073 5695 20131 5701
rect 20073 5692 20085 5695
rect 20036 5664 20085 5692
rect 20036 5652 20042 5664
rect 20073 5661 20085 5664
rect 20119 5661 20131 5695
rect 20073 5655 20131 5661
rect 20162 5652 20168 5704
rect 20220 5692 20226 5704
rect 20622 5692 20628 5704
rect 20220 5664 20628 5692
rect 20220 5652 20226 5664
rect 20622 5652 20628 5664
rect 20680 5692 20686 5704
rect 20717 5695 20775 5701
rect 20717 5692 20729 5695
rect 20680 5664 20729 5692
rect 20680 5652 20686 5664
rect 20717 5661 20729 5664
rect 20763 5692 20775 5695
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 20763 5664 21373 5692
rect 20763 5661 20775 5664
rect 20717 5655 20775 5661
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 22005 5695 22063 5701
rect 22005 5661 22017 5695
rect 22051 5661 22063 5695
rect 24762 5692 24768 5704
rect 24723 5664 24768 5692
rect 22005 5655 22063 5661
rect 10686 5624 10692 5636
rect 9968 5596 10692 5624
rect 8444 5584 8450 5596
rect 10686 5584 10692 5596
rect 10744 5584 10750 5636
rect 10778 5584 10784 5636
rect 10836 5624 10842 5636
rect 13173 5627 13231 5633
rect 10836 5596 10881 5624
rect 12084 5596 13124 5624
rect 10836 5584 10842 5596
rect 4120 5528 4292 5556
rect 4341 5559 4399 5565
rect 4120 5516 4126 5528
rect 4341 5525 4353 5559
rect 4387 5556 4399 5559
rect 4706 5556 4712 5568
rect 4387 5528 4712 5556
rect 4387 5525 4399 5528
rect 4341 5519 4399 5525
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 5534 5516 5540 5568
rect 5592 5516 5598 5568
rect 8662 5516 8668 5568
rect 8720 5556 8726 5568
rect 9582 5556 9588 5568
rect 8720 5528 9588 5556
rect 8720 5516 8726 5528
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 10502 5556 10508 5568
rect 9732 5528 10508 5556
rect 9732 5516 9738 5528
rect 10502 5516 10508 5528
rect 10560 5516 10566 5568
rect 11422 5516 11428 5568
rect 11480 5556 11486 5568
rect 12084 5556 12112 5596
rect 11480 5528 12112 5556
rect 13096 5556 13124 5596
rect 13173 5593 13185 5627
rect 13219 5624 13231 5627
rect 14550 5624 14556 5636
rect 13219 5596 14412 5624
rect 14511 5596 14556 5624
rect 13219 5593 13231 5596
rect 13173 5587 13231 5593
rect 13906 5556 13912 5568
rect 13096 5528 13912 5556
rect 11480 5516 11486 5528
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 14384 5556 14412 5596
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 17865 5627 17923 5633
rect 17865 5624 17877 5627
rect 15778 5596 17877 5624
rect 17865 5593 17877 5596
rect 17911 5593 17923 5627
rect 22020 5624 22048 5655
rect 24762 5652 24768 5664
rect 24820 5652 24826 5704
rect 29638 5652 29644 5704
rect 29696 5692 29702 5704
rect 35161 5695 35219 5701
rect 35161 5692 35173 5695
rect 29696 5664 35173 5692
rect 29696 5652 29702 5664
rect 35161 5661 35173 5664
rect 35207 5661 35219 5695
rect 38013 5695 38071 5701
rect 38013 5692 38025 5695
rect 35161 5655 35219 5661
rect 35866 5664 38025 5692
rect 22186 5624 22192 5636
rect 17865 5587 17923 5593
rect 19444 5596 22192 5624
rect 19444 5568 19472 5596
rect 22186 5584 22192 5596
rect 22244 5584 22250 5636
rect 17221 5559 17279 5565
rect 17221 5556 17233 5559
rect 14384 5528 17233 5556
rect 17221 5525 17233 5528
rect 17267 5525 17279 5559
rect 17221 5519 17279 5525
rect 19426 5516 19432 5568
rect 19484 5516 19490 5568
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 20165 5559 20223 5565
rect 20165 5556 20177 5559
rect 20036 5528 20177 5556
rect 20036 5516 20042 5528
rect 20165 5525 20177 5528
rect 20211 5525 20223 5559
rect 20165 5519 20223 5525
rect 24581 5559 24639 5565
rect 24581 5525 24593 5559
rect 24627 5556 24639 5559
rect 25682 5556 25688 5568
rect 24627 5528 25688 5556
rect 24627 5525 24639 5528
rect 24581 5519 24639 5525
rect 25682 5516 25688 5528
rect 25740 5516 25746 5568
rect 34977 5559 35035 5565
rect 34977 5525 34989 5559
rect 35023 5556 35035 5559
rect 35866 5556 35894 5664
rect 38013 5661 38025 5664
rect 38059 5661 38071 5695
rect 38013 5655 38071 5661
rect 38194 5556 38200 5568
rect 35023 5528 35894 5556
rect 38155 5528 38200 5556
rect 35023 5525 35035 5528
rect 34977 5519 35035 5525
rect 38194 5516 38200 5528
rect 38252 5516 38258 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 4801 5355 4859 5361
rect 4801 5352 4813 5355
rect 4028 5324 4813 5352
rect 4028 5312 4034 5324
rect 4801 5321 4813 5324
rect 4847 5321 4859 5355
rect 4801 5315 4859 5321
rect 5445 5355 5503 5361
rect 5445 5321 5457 5355
rect 5491 5352 5503 5355
rect 7006 5352 7012 5364
rect 5491 5324 7012 5352
rect 5491 5321 5503 5324
rect 5445 5315 5503 5321
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 10318 5352 10324 5364
rect 9140 5324 10324 5352
rect 6914 5284 6920 5296
rect 4172 5256 6920 5284
rect 1486 5176 1492 5228
rect 1544 5216 1550 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1544 5188 1593 5216
rect 1544 5176 1550 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 3786 5176 3792 5228
rect 3844 5176 3850 5228
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5117 2467 5151
rect 2682 5148 2688 5160
rect 2643 5120 2688 5148
rect 2409 5111 2467 5117
rect 1578 5040 1584 5092
rect 1636 5080 1642 5092
rect 2424 5080 2452 5111
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 4172 5157 4200 5256
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 8202 5284 8208 5296
rect 8142 5256 8208 5284
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 8665 5287 8723 5293
rect 8665 5253 8677 5287
rect 8711 5284 8723 5287
rect 9030 5284 9036 5296
rect 8711 5256 9036 5284
rect 8711 5253 8723 5256
rect 8665 5247 8723 5253
rect 9030 5244 9036 5256
rect 9088 5244 9094 5296
rect 4614 5176 4620 5228
rect 4672 5216 4678 5228
rect 9140 5225 9168 5324
rect 10318 5312 10324 5324
rect 10376 5352 10382 5364
rect 11698 5352 11704 5364
rect 10376 5324 11704 5352
rect 10376 5312 10382 5324
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 11808 5324 15148 5352
rect 11808 5284 11836 5324
rect 10626 5256 11836 5284
rect 11974 5244 11980 5296
rect 12032 5284 12038 5296
rect 12250 5284 12256 5296
rect 12032 5256 12256 5284
rect 12032 5244 12038 5256
rect 12250 5244 12256 5256
rect 12308 5244 12314 5296
rect 13446 5284 13452 5296
rect 13202 5256 13452 5284
rect 13446 5244 13452 5256
rect 13504 5244 13510 5296
rect 13630 5284 13636 5296
rect 13556 5256 13636 5284
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4672 5188 4721 5216
rect 4672 5176 4678 5188
rect 4709 5185 4721 5188
rect 4755 5216 4767 5219
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 4755 5188 5365 5216
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 5353 5185 5365 5188
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 11698 5216 11704 5228
rect 11659 5188 11704 5216
rect 9125 5179 9183 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 13556 5216 13584 5256
rect 13630 5244 13636 5256
rect 13688 5244 13694 5296
rect 14185 5287 14243 5293
rect 14185 5284 14197 5287
rect 13740 5256 14197 5284
rect 13372 5188 13584 5216
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5117 4215 5151
rect 6641 5151 6699 5157
rect 6641 5148 6653 5151
rect 4157 5111 4215 5117
rect 6012 5120 6653 5148
rect 1636 5052 2452 5080
rect 1636 5040 1642 5052
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 2424 5012 2452 5052
rect 6012 5024 6040 5120
rect 6641 5117 6653 5120
rect 6687 5117 6699 5151
rect 6914 5148 6920 5160
rect 6827 5120 6920 5148
rect 6641 5111 6699 5117
rect 6914 5108 6920 5120
rect 6972 5148 6978 5160
rect 7466 5148 7472 5160
rect 6972 5120 7472 5148
rect 6972 5108 6978 5120
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5148 9459 5151
rect 13372 5148 13400 5188
rect 9447 5120 13400 5148
rect 13449 5151 13507 5157
rect 9447 5117 9459 5120
rect 9401 5111 9459 5117
rect 13449 5117 13461 5151
rect 13495 5148 13507 5151
rect 13538 5148 13544 5160
rect 13495 5120 13544 5148
rect 13495 5117 13507 5120
rect 13449 5111 13507 5117
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 11606 5080 11612 5092
rect 10428 5052 11612 5080
rect 4062 5012 4068 5024
rect 2424 4984 4068 5012
rect 4062 4972 4068 4984
rect 4120 5012 4126 5024
rect 4982 5012 4988 5024
rect 4120 4984 4988 5012
rect 4120 4972 4126 4984
rect 4982 4972 4988 4984
rect 5040 5012 5046 5024
rect 5994 5012 6000 5024
rect 5040 4984 6000 5012
rect 5040 4972 5046 4984
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 10428 5012 10456 5052
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 13740 5080 13768 5256
rect 14185 5253 14197 5256
rect 14231 5253 14243 5287
rect 15120 5284 15148 5324
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 15252 5324 15301 5352
rect 15252 5312 15258 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 15289 5315 15347 5321
rect 15841 5355 15899 5361
rect 15841 5321 15853 5355
rect 15887 5352 15899 5355
rect 17034 5352 17040 5364
rect 15887 5324 17040 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 17310 5312 17316 5364
rect 17368 5352 17374 5364
rect 18877 5355 18935 5361
rect 18877 5352 18889 5355
rect 17368 5324 18889 5352
rect 17368 5312 17374 5324
rect 18877 5321 18889 5324
rect 18923 5321 18935 5355
rect 20070 5352 20076 5364
rect 18877 5315 18935 5321
rect 19628 5324 20076 5352
rect 17862 5284 17868 5296
rect 15120 5256 17868 5284
rect 14185 5247 14243 5253
rect 17862 5244 17868 5256
rect 17920 5244 17926 5296
rect 19518 5284 19524 5296
rect 19479 5256 19524 5284
rect 19518 5244 19524 5256
rect 19576 5244 19582 5296
rect 19628 5228 19656 5324
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 20809 5355 20867 5361
rect 20809 5321 20821 5355
rect 20855 5352 20867 5355
rect 21174 5352 21180 5364
rect 20855 5324 21180 5352
rect 20855 5321 20867 5324
rect 20809 5315 20867 5321
rect 21174 5312 21180 5324
rect 21232 5312 21238 5364
rect 31312 5324 31754 5352
rect 23382 5244 23388 5296
rect 23440 5284 23446 5296
rect 31312 5284 31340 5324
rect 23440 5256 31340 5284
rect 31726 5284 31754 5324
rect 31726 5256 35894 5284
rect 23440 5244 23446 5256
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5216 15255 5219
rect 15470 5216 15476 5228
rect 15243 5188 15476 5216
rect 15243 5185 15255 5188
rect 15197 5179 15255 5185
rect 15470 5176 15476 5188
rect 15528 5216 15534 5228
rect 15654 5216 15660 5228
rect 15528 5188 15660 5216
rect 15528 5176 15534 5188
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5216 16083 5219
rect 16114 5216 16120 5228
rect 16071 5188 16120 5216
rect 16071 5185 16083 5188
rect 16025 5179 16083 5185
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 16632 5188 16865 5216
rect 16632 5176 16638 5188
rect 16853 5185 16865 5188
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17681 5219 17739 5225
rect 17681 5216 17693 5219
rect 16991 5188 17693 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17681 5185 17693 5188
rect 17727 5185 17739 5219
rect 18138 5216 18144 5228
rect 18099 5188 18144 5216
rect 17681 5179 17739 5185
rect 18138 5176 18144 5188
rect 18196 5176 18202 5228
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5216 18843 5219
rect 19058 5216 19064 5228
rect 18831 5188 19064 5216
rect 18831 5185 18843 5188
rect 18785 5179 18843 5185
rect 19058 5176 19064 5188
rect 19116 5176 19122 5228
rect 19429 5219 19487 5225
rect 19429 5185 19441 5219
rect 19475 5216 19487 5219
rect 19610 5216 19616 5228
rect 19475 5188 19616 5216
rect 19475 5185 19487 5188
rect 19429 5179 19487 5185
rect 19610 5176 19616 5188
rect 19668 5176 19674 5228
rect 20070 5216 20076 5228
rect 19983 5188 20076 5216
rect 14090 5148 14096 5160
rect 14051 5120 14096 5148
rect 14090 5108 14096 5120
rect 14148 5108 14154 5160
rect 18046 5148 18052 5160
rect 14200 5120 18052 5148
rect 13004 5052 13768 5080
rect 6604 4984 10456 5012
rect 6604 4972 6610 4984
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 10873 5015 10931 5021
rect 10873 5012 10885 5015
rect 10560 4984 10885 5012
rect 10560 4972 10566 4984
rect 10873 4981 10885 4984
rect 10919 4981 10931 5015
rect 10873 4975 10931 4981
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 13004 5012 13032 5052
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 14200 5080 14228 5120
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 19334 5108 19340 5160
rect 19392 5148 19398 5160
rect 19996 5148 20024 5188
rect 20070 5176 20076 5188
rect 20128 5176 20134 5228
rect 20714 5216 20720 5228
rect 20675 5188 20720 5216
rect 20714 5176 20720 5188
rect 20772 5216 20778 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 20772 5188 22017 5216
rect 20772 5176 20778 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22646 5216 22652 5228
rect 22607 5188 22652 5216
rect 22005 5179 22063 5185
rect 22646 5176 22652 5188
rect 22704 5176 22710 5228
rect 31110 5216 31116 5228
rect 31071 5188 31116 5216
rect 31110 5176 31116 5188
rect 31168 5176 31174 5228
rect 31202 5176 31208 5228
rect 31260 5216 31266 5228
rect 32469 5219 32527 5225
rect 32469 5216 32481 5219
rect 31260 5188 31305 5216
rect 31726 5188 32481 5216
rect 31260 5176 31266 5188
rect 19392 5120 20024 5148
rect 19392 5108 19398 5120
rect 30006 5108 30012 5160
rect 30064 5148 30070 5160
rect 31726 5148 31754 5188
rect 32469 5185 32481 5188
rect 32515 5185 32527 5219
rect 35866 5216 35894 5256
rect 37461 5219 37519 5225
rect 37461 5216 37473 5219
rect 35866 5188 37473 5216
rect 32469 5179 32527 5185
rect 37461 5185 37473 5188
rect 37507 5185 37519 5219
rect 37461 5179 37519 5185
rect 37553 5219 37611 5225
rect 37553 5185 37565 5219
rect 37599 5216 37611 5219
rect 38289 5219 38347 5225
rect 38289 5216 38301 5219
rect 37599 5188 38301 5216
rect 37599 5185 37611 5188
rect 37553 5179 37611 5185
rect 38289 5185 38301 5188
rect 38335 5185 38347 5219
rect 38289 5179 38347 5185
rect 30064 5120 31754 5148
rect 30064 5108 30070 5120
rect 13872 5052 14228 5080
rect 13872 5040 13878 5052
rect 14458 5040 14464 5092
rect 14516 5080 14522 5092
rect 14645 5083 14703 5089
rect 14645 5080 14657 5083
rect 14516 5052 14657 5080
rect 14516 5040 14522 5052
rect 14645 5049 14657 5052
rect 14691 5049 14703 5083
rect 14645 5043 14703 5049
rect 14734 5040 14740 5092
rect 14792 5080 14798 5092
rect 18233 5083 18291 5089
rect 18233 5080 18245 5083
rect 14792 5052 18245 5080
rect 14792 5040 14798 5052
rect 18233 5049 18245 5052
rect 18279 5049 18291 5083
rect 18233 5043 18291 5049
rect 22094 5040 22100 5092
rect 22152 5080 22158 5092
rect 22152 5052 22197 5080
rect 22152 5040 22158 5052
rect 31110 5040 31116 5092
rect 31168 5080 31174 5092
rect 34422 5080 34428 5092
rect 31168 5052 34428 5080
rect 31168 5040 31174 5052
rect 34422 5040 34428 5052
rect 34480 5040 34486 5092
rect 11112 4984 13032 5012
rect 11112 4972 11118 4984
rect 13630 4972 13636 5024
rect 13688 5012 13694 5024
rect 15470 5012 15476 5024
rect 13688 4984 15476 5012
rect 13688 4972 13694 4984
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 15930 4972 15936 5024
rect 15988 5012 15994 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 15988 4984 17509 5012
rect 15988 4972 15994 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 20165 5015 20223 5021
rect 20165 4981 20177 5015
rect 20211 5012 20223 5015
rect 20622 5012 20628 5024
rect 20211 4984 20628 5012
rect 20211 4981 20223 4984
rect 20165 4975 20223 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 22370 4972 22376 5024
rect 22428 5012 22434 5024
rect 22741 5015 22799 5021
rect 22741 5012 22753 5015
rect 22428 4984 22753 5012
rect 22428 4972 22434 4984
rect 22741 4981 22753 4984
rect 22787 4981 22799 5015
rect 22741 4975 22799 4981
rect 32309 5015 32367 5021
rect 32309 4981 32321 5015
rect 32355 5012 32367 5015
rect 35802 5012 35808 5024
rect 32355 4984 35808 5012
rect 32355 4981 32367 4984
rect 32309 4975 32367 4981
rect 35802 4972 35808 4984
rect 35860 4972 35866 5024
rect 38010 4972 38016 5024
rect 38068 5012 38074 5024
rect 38105 5015 38163 5021
rect 38105 5012 38117 5015
rect 38068 4984 38117 5012
rect 38068 4972 38074 4984
rect 38105 4981 38117 4984
rect 38151 4981 38163 5015
rect 38105 4975 38163 4981
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 6546 4808 6552 4820
rect 2746 4780 6552 4808
rect 2746 4684 2774 4780
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 8386 4808 8392 4820
rect 7791 4780 8392 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9140 4780 9352 4808
rect 7101 4743 7159 4749
rect 7101 4709 7113 4743
rect 7147 4740 7159 4743
rect 9140 4740 9168 4780
rect 7147 4712 9168 4740
rect 9324 4740 9352 4780
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 15930 4808 15936 4820
rect 9456 4780 15936 4808
rect 9456 4768 9462 4780
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 16114 4808 16120 4820
rect 16075 4780 16120 4808
rect 16114 4768 16120 4780
rect 16172 4768 16178 4820
rect 17494 4808 17500 4820
rect 17455 4780 17500 4808
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 19521 4811 19579 4817
rect 19521 4777 19533 4811
rect 19567 4808 19579 4811
rect 20346 4808 20352 4820
rect 19567 4780 20352 4808
rect 19567 4777 19579 4780
rect 19521 4771 19579 4777
rect 20346 4768 20352 4780
rect 20404 4768 20410 4820
rect 20809 4811 20867 4817
rect 20809 4777 20821 4811
rect 20855 4808 20867 4811
rect 21082 4808 21088 4820
rect 20855 4780 21088 4808
rect 20855 4777 20867 4780
rect 20809 4771 20867 4777
rect 21082 4768 21088 4780
rect 21140 4768 21146 4820
rect 21453 4811 21511 4817
rect 21453 4777 21465 4811
rect 21499 4808 21511 4811
rect 21542 4808 21548 4820
rect 21499 4780 21548 4808
rect 21499 4777 21511 4780
rect 21453 4771 21511 4777
rect 21542 4768 21548 4780
rect 21600 4768 21606 4820
rect 12342 4740 12348 4752
rect 9324 4712 10732 4740
rect 7147 4709 7159 4712
rect 7101 4703 7159 4709
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4672 2191 4675
rect 2314 4672 2320 4684
rect 2179 4644 2320 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 2682 4632 2688 4684
rect 2740 4644 2774 4684
rect 6546 4672 6552 4684
rect 6507 4644 6552 4672
rect 2740 4632 2746 4644
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 8996 4644 9168 4672
rect 8996 4632 9002 4644
rect 1854 4604 1860 4616
rect 1815 4576 1860 4604
rect 1854 4564 1860 4576
rect 1912 4564 1918 4616
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 2958 4604 2964 4616
rect 2915 4576 2964 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 4120 4576 4537 4604
rect 4120 4564 4126 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4604 7343 4607
rect 7742 4604 7748 4616
rect 7331 4576 7748 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4604 7987 4607
rect 8294 4604 8300 4616
rect 7975 4576 8300 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 9030 4604 9036 4616
rect 8435 4576 9036 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 3142 4536 3148 4548
rect 3103 4508 3148 4536
rect 3142 4496 3148 4508
rect 3200 4496 3206 4548
rect 4801 4539 4859 4545
rect 4801 4505 4813 4539
rect 4847 4505 4859 4539
rect 6454 4536 6460 4548
rect 6026 4508 6460 4536
rect 4801 4499 4859 4505
rect 4816 4468 4844 4499
rect 6454 4496 6460 4508
rect 6512 4496 6518 4548
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 8404 4536 8432 4567
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 9140 4613 9168 4644
rect 9398 4632 9404 4684
rect 9456 4672 9462 4684
rect 10134 4672 10140 4684
rect 9456 4644 10140 4672
rect 9456 4632 9462 4644
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10318 4632 10324 4684
rect 10376 4672 10382 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 10376 4644 10609 4672
rect 10376 4632 10382 4644
rect 10597 4641 10609 4644
rect 10643 4641 10655 4675
rect 10704 4672 10732 4712
rect 11900 4712 12348 4740
rect 11900 4672 11928 4712
rect 12342 4700 12348 4712
rect 12400 4700 12406 4752
rect 13814 4740 13820 4752
rect 13372 4712 13820 4740
rect 10704 4644 11928 4672
rect 10597 4635 10655 4641
rect 12986 4632 12992 4684
rect 13044 4672 13050 4684
rect 13265 4675 13323 4681
rect 13044 4644 13216 4672
rect 13044 4632 13050 4644
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 9950 4604 9956 4616
rect 9364 4576 9956 4604
rect 9364 4564 9370 4576
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 12250 4564 12256 4616
rect 12308 4604 12314 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 12308 4576 12633 4604
rect 12308 4564 12314 4576
rect 12621 4573 12633 4576
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4573 13139 4607
rect 13188 4604 13216 4644
rect 13265 4641 13277 4675
rect 13311 4672 13323 4675
rect 13372 4672 13400 4712
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 15378 4700 15384 4752
rect 15436 4740 15442 4752
rect 15565 4743 15623 4749
rect 15565 4740 15577 4743
rect 15436 4712 15577 4740
rect 15436 4700 15442 4712
rect 15565 4709 15577 4712
rect 15611 4709 15623 4743
rect 15565 4703 15623 4709
rect 18601 4743 18659 4749
rect 18601 4709 18613 4743
rect 18647 4740 18659 4743
rect 21910 4740 21916 4752
rect 18647 4712 21916 4740
rect 18647 4709 18659 4712
rect 18601 4703 18659 4709
rect 21910 4700 21916 4712
rect 21968 4700 21974 4752
rect 13311 4644 13400 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 13906 4632 13912 4684
rect 13964 4672 13970 4684
rect 18138 4672 18144 4684
rect 13964 4644 15516 4672
rect 13964 4632 13970 4644
rect 13725 4607 13783 4613
rect 13725 4604 13737 4607
rect 13188 4576 13737 4604
rect 13081 4567 13139 4573
rect 13725 4573 13737 4576
rect 13771 4604 13783 4607
rect 13771 4576 14228 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 7156 4508 8432 4536
rect 8481 4539 8539 4545
rect 7156 4496 7162 4508
rect 8481 4505 8493 4539
rect 8527 4536 8539 4539
rect 10873 4539 10931 4545
rect 8527 4508 10824 4536
rect 8527 4505 8539 4508
rect 8481 4499 8539 4505
rect 6362 4468 6368 4480
rect 4816 4440 6368 4468
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 9030 4428 9036 4480
rect 9088 4468 9094 4480
rect 9309 4471 9367 4477
rect 9309 4468 9321 4471
rect 9088 4440 9321 4468
rect 9088 4428 9094 4440
rect 9309 4437 9321 4440
rect 9355 4437 9367 4471
rect 10042 4468 10048 4480
rect 10003 4440 10048 4468
rect 9309 4431 9367 4437
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 10796 4468 10824 4508
rect 10873 4505 10885 4539
rect 10919 4536 10931 4539
rect 10962 4536 10968 4548
rect 10919 4508 10968 4536
rect 10919 4505 10931 4508
rect 10873 4499 10931 4505
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 12710 4536 12716 4548
rect 12098 4508 12716 4536
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 13096 4536 13124 4567
rect 14200 4536 14228 4576
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 15488 4613 15516 4644
rect 16316 4644 18144 4672
rect 15473 4607 15531 4613
rect 15068 4576 15113 4604
rect 15068 4564 15074 4576
rect 15473 4573 15485 4607
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 16206 4564 16212 4616
rect 16264 4604 16270 4616
rect 16316 4613 16344 4644
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 20165 4675 20223 4681
rect 20165 4641 20177 4675
rect 20211 4672 20223 4675
rect 20438 4672 20444 4684
rect 20211 4644 20444 4672
rect 20211 4641 20223 4644
rect 20165 4635 20223 4641
rect 20438 4632 20444 4644
rect 20496 4632 20502 4684
rect 16301 4607 16359 4613
rect 16301 4604 16313 4607
rect 16264 4576 16313 4604
rect 16264 4564 16270 4576
rect 16301 4573 16313 4576
rect 16347 4573 16359 4607
rect 16758 4604 16764 4616
rect 16719 4576 16764 4604
rect 16301 4567 16359 4573
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 16942 4564 16948 4616
rect 17000 4604 17006 4616
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 17000 4576 17417 4604
rect 17000 4564 17006 4576
rect 17405 4573 17417 4576
rect 17451 4604 17463 4607
rect 17954 4604 17960 4616
rect 17451 4576 17960 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 17954 4564 17960 4576
rect 18012 4604 18018 4616
rect 18414 4604 18420 4616
rect 18012 4576 18420 4604
rect 18012 4564 18018 4576
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 18782 4604 18788 4616
rect 18743 4576 18788 4604
rect 18782 4564 18788 4576
rect 18840 4564 18846 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19076 4576 19441 4604
rect 14369 4539 14427 4545
rect 14369 4536 14381 4539
rect 13096 4508 13860 4536
rect 14200 4508 14381 4536
rect 13630 4468 13636 4480
rect 10796 4440 13636 4468
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 13832 4468 13860 4508
rect 14369 4505 14381 4508
rect 14415 4505 14427 4539
rect 14369 4499 14427 4505
rect 14461 4539 14519 4545
rect 14461 4505 14473 4539
rect 14507 4536 14519 4539
rect 14734 4536 14740 4548
rect 14507 4508 14740 4536
rect 14507 4505 14519 4508
rect 14461 4499 14519 4505
rect 14734 4496 14740 4508
rect 14792 4496 14798 4548
rect 16853 4539 16911 4545
rect 16853 4536 16865 4539
rect 15120 4508 16865 4536
rect 15120 4468 15148 4508
rect 16853 4505 16865 4508
rect 16899 4505 16911 4539
rect 18432 4536 18460 4564
rect 19076 4548 19104 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 20070 4604 20076 4616
rect 20031 4576 20076 4604
rect 19429 4567 19487 4573
rect 20070 4564 20076 4576
rect 20128 4604 20134 4616
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 20128 4576 20729 4604
rect 20128 4564 20134 4576
rect 20717 4573 20729 4576
rect 20763 4604 20775 4607
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 20763 4576 21373 4604
rect 20763 4573 20775 4576
rect 20717 4567 20775 4573
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21997 4607 22055 4613
rect 21997 4604 22009 4607
rect 21361 4567 21419 4573
rect 21928 4576 22009 4604
rect 19058 4536 19064 4548
rect 18432 4508 19064 4536
rect 16853 4499 16911 4505
rect 19058 4496 19064 4508
rect 19116 4496 19122 4548
rect 13832 4440 15148 4468
rect 15470 4428 15476 4480
rect 15528 4468 15534 4480
rect 19426 4468 19432 4480
rect 15528 4440 19432 4468
rect 15528 4428 15534 4440
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 20070 4468 20076 4480
rect 19668 4440 20076 4468
rect 19668 4428 19674 4440
rect 20070 4428 20076 4440
rect 20128 4468 20134 4480
rect 21928 4468 21956 4576
rect 21997 4573 22009 4576
rect 22043 4573 22055 4607
rect 21997 4567 22055 4573
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 22244 4576 22661 4604
rect 22244 4564 22250 4576
rect 22649 4573 22661 4576
rect 22695 4604 22707 4607
rect 23106 4604 23112 4616
rect 22695 4576 23112 4604
rect 22695 4573 22707 4576
rect 22649 4567 22707 4573
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 22094 4496 22100 4548
rect 22152 4536 22158 4548
rect 22152 4508 22197 4536
rect 22152 4496 22158 4508
rect 22002 4468 22008 4480
rect 20128 4440 22008 4468
rect 20128 4428 20134 4440
rect 22002 4428 22008 4440
rect 22060 4428 22066 4480
rect 22738 4468 22744 4480
rect 22699 4440 22744 4468
rect 22738 4428 22744 4440
rect 22796 4428 22802 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 3142 4224 3148 4276
rect 3200 4264 3206 4276
rect 5905 4267 5963 4273
rect 3200 4236 5764 4264
rect 3200 4224 3206 4236
rect 5166 4156 5172 4208
rect 5224 4156 5230 4208
rect 5736 4196 5764 4236
rect 5905 4233 5917 4267
rect 5951 4264 5963 4267
rect 6362 4264 6368 4276
rect 5951 4236 6368 4264
rect 5951 4233 5963 4236
rect 5905 4227 5963 4233
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 8018 4224 8024 4276
rect 8076 4264 8082 4276
rect 11974 4264 11980 4276
rect 8076 4236 11980 4264
rect 8076 4224 8082 4236
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12066 4224 12072 4276
rect 12124 4264 12130 4276
rect 13446 4264 13452 4276
rect 12124 4236 13452 4264
rect 12124 4224 12130 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 22738 4264 22744 4276
rect 13556 4236 22744 4264
rect 7650 4196 7656 4208
rect 5736 4168 7656 4196
rect 7650 4156 7656 4168
rect 7708 4156 7714 4208
rect 9582 4196 9588 4208
rect 9246 4168 9588 4196
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 12250 4196 12256 4208
rect 9824 4168 12256 4196
rect 9824 4156 9830 4168
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 13556 4196 13584 4236
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 13202 4168 13584 4196
rect 13630 4156 13636 4208
rect 13688 4196 13694 4208
rect 13688 4168 14766 4196
rect 13688 4156 13694 4168
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 17865 4199 17923 4205
rect 17865 4196 17877 4199
rect 17184 4168 17877 4196
rect 17184 4156 17190 4168
rect 17865 4165 17877 4168
rect 17911 4165 17923 4199
rect 17865 4159 17923 4165
rect 18340 4168 18644 4196
rect 1854 4128 1860 4140
rect 1815 4100 1860 4128
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2958 4128 2964 4140
rect 2919 4100 2964 4128
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 7098 4128 7104 4140
rect 5776 4100 7104 4128
rect 5776 4088 5782 4100
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 9306 4088 9312 4140
rect 9364 4128 9370 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 9364 4100 10517 4128
rect 9364 4088 9370 4100
rect 10505 4097 10517 4100
rect 10551 4128 10563 4131
rect 10965 4131 11023 4137
rect 10965 4128 10977 4131
rect 10551 4100 10977 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 10965 4097 10977 4100
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11698 4128 11704 4140
rect 11112 4100 11157 4128
rect 11659 4100 11704 4128
rect 11112 4088 11118 4100
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4128 17371 4131
rect 17678 4128 17684 4140
rect 17359 4100 17684 4128
rect 17359 4097 17371 4100
rect 17313 4091 17371 4097
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 17773 4131 17831 4137
rect 17773 4097 17785 4131
rect 17819 4128 17831 4131
rect 18340 4128 18368 4168
rect 17819 4100 18368 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 3234 4060 3240 4072
rect 2179 4032 2774 4060
rect 3195 4032 3240 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 2746 3924 2774 4032
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4157 4063 4215 4069
rect 4157 4060 4169 4063
rect 4120 4032 4169 4060
rect 4120 4020 4126 4032
rect 4157 4029 4169 4032
rect 4203 4029 4215 4063
rect 4157 4023 4215 4029
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 4479 4032 5948 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 5920 3992 5948 4032
rect 5994 4020 6000 4072
rect 6052 4060 6058 4072
rect 7466 4060 7472 4072
rect 6052 4032 7472 4060
rect 6052 4020 6058 4032
rect 7466 4020 7472 4032
rect 7524 4060 7530 4072
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7524 4032 7757 4060
rect 7524 4020 7530 4032
rect 7745 4029 7757 4032
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 9674 4060 9680 4072
rect 8067 4032 9680 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 9824 4032 9869 4060
rect 9824 4020 9830 4032
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 11422 4060 11428 4072
rect 10008 4032 11428 4060
rect 10008 4020 10014 4032
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11974 4060 11980 4072
rect 11935 4032 11980 4060
rect 11974 4020 11980 4032
rect 12032 4060 12038 4072
rect 13722 4060 13728 4072
rect 12032 4032 13728 4060
rect 12032 4020 12038 4032
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 13998 4060 14004 4072
rect 13959 4032 14004 4060
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 14108 4032 14289 4060
rect 7282 3992 7288 4004
rect 5920 3964 7288 3992
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 10226 3952 10232 4004
rect 10284 3992 10290 4004
rect 14108 3992 14136 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 17586 4020 17592 4072
rect 17644 4060 17650 4072
rect 17788 4060 17816 4091
rect 18414 4088 18420 4140
rect 18472 4128 18478 4140
rect 18472 4100 18517 4128
rect 18472 4088 18478 4100
rect 17644 4032 17816 4060
rect 17644 4020 17650 4032
rect 17862 4020 17868 4072
rect 17920 4060 17926 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 17920 4032 18521 4060
rect 17920 4020 17926 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18616 4060 18644 4168
rect 19426 4156 19432 4208
rect 19484 4196 19490 4208
rect 19484 4168 20392 4196
rect 19484 4156 19490 4168
rect 19058 4088 19064 4140
rect 19116 4128 19122 4140
rect 20364 4137 20392 4168
rect 19705 4131 19763 4137
rect 19116 4100 19161 4128
rect 19116 4088 19122 4100
rect 19705 4097 19717 4131
rect 19751 4097 19763 4131
rect 19705 4091 19763 4097
rect 20349 4131 20407 4137
rect 20349 4097 20361 4131
rect 20395 4097 20407 4131
rect 20349 4091 20407 4097
rect 19334 4060 19340 4072
rect 18616 4032 19340 4060
rect 18509 4023 18567 4029
rect 19334 4020 19340 4032
rect 19392 4060 19398 4072
rect 19720 4060 19748 4091
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20772 4100 21005 4128
rect 20772 4088 20778 4100
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 22002 4128 22008 4140
rect 21963 4100 22008 4128
rect 20993 4091 21051 4097
rect 22002 4088 22008 4100
rect 22060 4128 22066 4140
rect 22646 4128 22652 4140
rect 22060 4100 22652 4128
rect 22060 4088 22066 4100
rect 22646 4088 22652 4100
rect 22704 4088 22710 4140
rect 26694 4088 26700 4140
rect 26752 4128 26758 4140
rect 27341 4131 27399 4137
rect 27341 4128 27353 4131
rect 26752 4100 27353 4128
rect 26752 4088 26758 4100
rect 27341 4097 27353 4100
rect 27387 4097 27399 4131
rect 27341 4091 27399 4097
rect 19392 4032 19748 4060
rect 19392 4020 19398 4032
rect 19794 4020 19800 4072
rect 19852 4060 19858 4072
rect 26602 4060 26608 4072
rect 19852 4032 26608 4060
rect 19852 4020 19858 4032
rect 26602 4020 26608 4032
rect 26660 4020 26666 4072
rect 16850 3992 16856 4004
rect 10284 3964 11192 3992
rect 10284 3952 10290 3964
rect 4614 3924 4620 3936
rect 2746 3896 4620 3924
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5442 3884 5448 3936
rect 5500 3924 5506 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 5500 3896 7205 3924
rect 5500 3884 5506 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 7193 3887 7251 3893
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 10410 3884 10416 3936
rect 10468 3924 10474 3936
rect 11054 3924 11060 3936
rect 10468 3896 11060 3924
rect 10468 3884 10474 3896
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11164 3924 11192 3964
rect 13004 3964 14136 3992
rect 15580 3964 16856 3992
rect 12434 3924 12440 3936
rect 11164 3896 12440 3924
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 13004 3924 13032 3964
rect 12584 3896 13032 3924
rect 13449 3927 13507 3933
rect 12584 3884 12590 3896
rect 13449 3893 13461 3927
rect 13495 3924 13507 3927
rect 14366 3924 14372 3936
rect 13495 3896 14372 3924
rect 13495 3893 13507 3896
rect 13449 3887 13507 3893
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 14458 3884 14464 3936
rect 14516 3924 14522 3936
rect 15580 3924 15608 3964
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 17129 3995 17187 4001
rect 17129 3961 17141 3995
rect 17175 3992 17187 3995
rect 19426 3992 19432 4004
rect 17175 3964 19432 3992
rect 17175 3961 17187 3964
rect 17129 3955 17187 3961
rect 19426 3952 19432 3964
rect 19484 3952 19490 4004
rect 20806 3952 20812 4004
rect 20864 3992 20870 4004
rect 22741 3995 22799 4001
rect 22741 3992 22753 3995
rect 20864 3964 22753 3992
rect 20864 3952 20870 3964
rect 22741 3961 22753 3964
rect 22787 3961 22799 3995
rect 22741 3955 22799 3961
rect 14516 3896 15608 3924
rect 14516 3884 14522 3896
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 15749 3927 15807 3933
rect 15749 3924 15761 3927
rect 15712 3896 15761 3924
rect 15712 3884 15718 3896
rect 15749 3893 15761 3896
rect 15795 3893 15807 3927
rect 19150 3924 19156 3936
rect 19111 3896 19156 3924
rect 15749 3887 15807 3893
rect 19150 3884 19156 3896
rect 19208 3884 19214 3936
rect 19242 3884 19248 3936
rect 19300 3924 19306 3936
rect 19797 3927 19855 3933
rect 19797 3924 19809 3927
rect 19300 3896 19809 3924
rect 19300 3884 19306 3896
rect 19797 3893 19809 3896
rect 19843 3893 19855 3927
rect 19797 3887 19855 3893
rect 20441 3927 20499 3933
rect 20441 3893 20453 3927
rect 20487 3924 20499 3927
rect 20530 3924 20536 3936
rect 20487 3896 20536 3924
rect 20487 3893 20499 3896
rect 20441 3887 20499 3893
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 20898 3884 20904 3936
rect 20956 3924 20962 3936
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20956 3896 21097 3924
rect 20956 3884 20962 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 22097 3927 22155 3933
rect 22097 3893 22109 3927
rect 22143 3924 22155 3927
rect 22278 3924 22284 3936
rect 22143 3896 22284 3924
rect 22143 3893 22155 3896
rect 22097 3887 22155 3893
rect 22278 3884 22284 3896
rect 22336 3884 22342 3936
rect 27157 3927 27215 3933
rect 27157 3893 27169 3927
rect 27203 3924 27215 3927
rect 28902 3924 28908 3936
rect 27203 3896 28908 3924
rect 27203 3893 27215 3896
rect 27157 3887 27215 3893
rect 28902 3884 28908 3896
rect 28960 3884 28966 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 10226 3720 10232 3732
rect 2884 3692 10232 3720
rect 2884 3593 2912 3692
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 10318 3680 10324 3732
rect 10376 3720 10382 3732
rect 10376 3692 16804 3720
rect 10376 3680 10382 3692
rect 3234 3612 3240 3664
rect 3292 3652 3298 3664
rect 13722 3652 13728 3664
rect 3292 3624 6132 3652
rect 3292 3612 3298 3624
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 5626 3584 5632 3596
rect 4295 3556 5632 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 5994 3584 6000 3596
rect 5955 3556 6000 3584
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 6104 3584 6132 3624
rect 10980 3624 12112 3652
rect 13683 3624 13728 3652
rect 9766 3584 9772 3596
rect 6104 3556 9772 3584
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 2590 3516 2596 3528
rect 2551 3488 2596 3516
rect 1673 3479 1731 3485
rect 1688 3380 1716 3479
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3016 3488 3985 3516
rect 3016 3476 3022 3488
rect 3973 3485 3985 3488
rect 4019 3516 4031 3519
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4019 3488 4905 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4893 3485 4905 3488
rect 4939 3516 4951 3519
rect 5718 3516 5724 3528
rect 4939 3488 5724 3516
rect 4939 3485 4951 3488
rect 4893 3479 4951 3485
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 8018 3516 8024 3528
rect 7979 3488 8024 3516
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9364 3488 9505 3516
rect 9364 3476 9370 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 10980 3516 11008 3624
rect 11514 3584 11520 3596
rect 11475 3556 11520 3584
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 11698 3544 11704 3596
rect 11756 3584 11762 3596
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 11756 3556 11989 3584
rect 11756 3544 11762 3556
rect 11977 3553 11989 3556
rect 12023 3553 12035 3587
rect 12084 3584 12112 3624
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 16022 3652 16028 3664
rect 15983 3624 16028 3652
rect 16022 3612 16028 3624
rect 16080 3612 16086 3664
rect 16577 3655 16635 3661
rect 16577 3621 16589 3655
rect 16623 3621 16635 3655
rect 16577 3615 16635 3621
rect 13446 3584 13452 3596
rect 12084 3556 13452 3584
rect 11977 3547 12035 3553
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 16592 3584 16620 3615
rect 13648 3556 16620 3584
rect 10902 3488 11008 3516
rect 9493 3479 9551 3485
rect 1949 3451 2007 3457
rect 1949 3417 1961 3451
rect 1995 3448 2007 3451
rect 5074 3448 5080 3460
rect 1995 3420 5080 3448
rect 1995 3417 2007 3420
rect 1949 3411 2007 3417
rect 5074 3408 5080 3420
rect 5132 3408 5138 3460
rect 5169 3451 5227 3457
rect 5169 3417 5181 3451
rect 5215 3417 5227 3451
rect 5169 3411 5227 3417
rect 1854 3380 1860 3392
rect 1688 3352 1860 3380
rect 1854 3340 1860 3352
rect 1912 3380 1918 3392
rect 3510 3380 3516 3392
rect 1912 3352 3516 3380
rect 1912 3340 1918 3352
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 5184 3380 5212 3411
rect 5810 3408 5816 3460
rect 5868 3448 5874 3460
rect 6273 3451 6331 3457
rect 6273 3448 6285 3451
rect 5868 3420 6285 3448
rect 5868 3408 5874 3420
rect 6273 3417 6285 3420
rect 6319 3417 6331 3451
rect 7834 3448 7840 3460
rect 7498 3420 7840 3448
rect 6273 3411 6331 3417
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 9766 3448 9772 3460
rect 9727 3420 9772 3448
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 12158 3448 12164 3460
rect 11480 3420 12164 3448
rect 11480 3408 11486 3420
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 12250 3408 12256 3460
rect 12308 3448 12314 3460
rect 13538 3448 13544 3460
rect 12308 3420 12353 3448
rect 13478 3420 13544 3448
rect 12308 3408 12314 3420
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 10410 3380 10416 3392
rect 5184 3352 10416 3380
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 10686 3340 10692 3392
rect 10744 3380 10750 3392
rect 13648 3380 13676 3556
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14274 3516 14280 3528
rect 14056 3488 14280 3516
rect 14056 3476 14062 3488
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 16776 3525 16804 3692
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 19242 3720 19248 3732
rect 17460 3692 19248 3720
rect 17460 3680 17466 3692
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 19518 3720 19524 3732
rect 19479 3692 19524 3720
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 21450 3720 21456 3732
rect 21411 3692 21456 3720
rect 21450 3680 21456 3692
rect 21508 3680 21514 3732
rect 22462 3720 22468 3732
rect 22423 3692 22468 3720
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 23198 3680 23204 3732
rect 23256 3720 23262 3732
rect 23293 3723 23351 3729
rect 23293 3720 23305 3723
rect 23256 3692 23305 3720
rect 23256 3680 23262 3692
rect 23293 3689 23305 3692
rect 23339 3689 23351 3723
rect 26694 3720 26700 3732
rect 26655 3692 26700 3720
rect 23293 3683 23351 3689
rect 26694 3680 26700 3692
rect 26752 3680 26758 3732
rect 31386 3680 31392 3732
rect 31444 3720 31450 3732
rect 38105 3723 38163 3729
rect 38105 3720 38117 3723
rect 31444 3692 38117 3720
rect 31444 3680 31450 3692
rect 38105 3689 38117 3692
rect 38151 3689 38163 3723
rect 38105 3683 38163 3689
rect 16850 3612 16856 3664
rect 16908 3652 16914 3664
rect 19794 3652 19800 3664
rect 16908 3624 19800 3652
rect 16908 3612 16914 3624
rect 19794 3612 19800 3624
rect 19852 3612 19858 3664
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 18601 3587 18659 3593
rect 18601 3584 18613 3587
rect 18288 3556 18613 3584
rect 18288 3544 18294 3556
rect 18601 3553 18613 3556
rect 18647 3553 18659 3587
rect 18601 3547 18659 3553
rect 19444 3556 20760 3584
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 16908 3488 17233 3516
rect 16908 3476 16914 3488
rect 17221 3485 17233 3488
rect 17267 3516 17279 3519
rect 17862 3516 17868 3528
rect 17267 3488 17868 3516
rect 17267 3485 17279 3488
rect 17221 3479 17279 3485
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 18472 3488 18521 3516
rect 18472 3476 18478 3488
rect 18509 3485 18521 3488
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 13722 3408 13728 3460
rect 13780 3448 13786 3460
rect 14458 3448 14464 3460
rect 13780 3420 14464 3448
rect 13780 3408 13786 3420
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 14553 3451 14611 3457
rect 14553 3417 14565 3451
rect 14599 3448 14611 3451
rect 14826 3448 14832 3460
rect 14599 3420 14832 3448
rect 14599 3417 14611 3420
rect 14553 3411 14611 3417
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 17313 3451 17371 3457
rect 17313 3448 17325 3451
rect 15778 3420 17325 3448
rect 17313 3417 17325 3420
rect 17359 3417 17371 3451
rect 18524 3448 18552 3479
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19444 3525 19472 3556
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 19392 3488 19441 3516
rect 19392 3476 19398 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 20070 3516 20076 3528
rect 20031 3488 20076 3516
rect 19429 3479 19487 3485
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 20732 3525 20760 3556
rect 22094 3544 22100 3596
rect 22152 3584 22158 3596
rect 22152 3556 22692 3584
rect 22152 3544 22158 3556
rect 22664 3525 22692 3556
rect 20717 3519 20775 3525
rect 20717 3485 20729 3519
rect 20763 3516 20775 3519
rect 21361 3519 21419 3525
rect 21361 3516 21373 3519
rect 20763 3488 21373 3516
rect 20763 3485 20775 3488
rect 20717 3479 20775 3485
rect 21361 3485 21373 3488
rect 21407 3485 21419 3519
rect 21361 3479 21419 3485
rect 22649 3519 22707 3525
rect 22649 3485 22661 3519
rect 22695 3485 22707 3519
rect 22649 3479 22707 3485
rect 22741 3519 22799 3525
rect 22741 3485 22753 3519
rect 22787 3485 22799 3519
rect 23474 3516 23480 3528
rect 23435 3488 23480 3516
rect 22741 3479 22799 3485
rect 22756 3448 22784 3479
rect 23474 3476 23480 3488
rect 23532 3516 23538 3528
rect 23753 3519 23811 3525
rect 23753 3516 23765 3519
rect 23532 3488 23765 3516
rect 23532 3476 23538 3488
rect 23753 3485 23765 3488
rect 23799 3485 23811 3519
rect 26602 3516 26608 3528
rect 26563 3488 26608 3516
rect 23753 3479 23811 3485
rect 26602 3476 26608 3488
rect 26660 3476 26666 3528
rect 38286 3516 38292 3528
rect 38247 3488 38292 3516
rect 38286 3476 38292 3488
rect 38344 3476 38350 3528
rect 18524 3420 22784 3448
rect 17313 3411 17371 3417
rect 17954 3380 17960 3392
rect 10744 3352 13676 3380
rect 17915 3352 17960 3380
rect 10744 3340 10750 3352
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 20070 3340 20076 3392
rect 20128 3380 20134 3392
rect 20165 3383 20223 3389
rect 20165 3380 20177 3383
rect 20128 3352 20177 3380
rect 20128 3340 20134 3352
rect 20165 3349 20177 3352
rect 20211 3349 20223 3383
rect 20165 3343 20223 3349
rect 20346 3340 20352 3392
rect 20404 3380 20410 3392
rect 20809 3383 20867 3389
rect 20809 3380 20821 3383
rect 20404 3352 20821 3380
rect 20404 3340 20410 3352
rect 20809 3349 20821 3352
rect 20855 3349 20867 3383
rect 22830 3380 22836 3392
rect 22791 3352 22836 3380
rect 20809 3343 20867 3349
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 6917 3179 6975 3185
rect 6917 3145 6929 3179
rect 6963 3176 6975 3179
rect 7098 3176 7104 3188
rect 6963 3148 7104 3176
rect 6963 3145 6975 3148
rect 6917 3139 6975 3145
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 12158 3176 12164 3188
rect 8220 3148 12164 3176
rect 3878 3108 3884 3120
rect 3082 3080 3884 3108
rect 3878 3068 3884 3080
rect 3936 3068 3942 3120
rect 8110 3108 8116 3120
rect 5658 3080 8116 3108
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 8220 3117 8248 3148
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 12986 3176 12992 3188
rect 12400 3148 12992 3176
rect 12400 3136 12406 3148
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 13449 3179 13507 3185
rect 13449 3176 13461 3179
rect 13412 3148 13461 3176
rect 13412 3136 13418 3148
rect 13449 3145 13461 3148
rect 13495 3145 13507 3179
rect 13449 3139 13507 3145
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 18141 3179 18199 3185
rect 18141 3176 18153 3179
rect 13688 3148 18153 3176
rect 13688 3136 13694 3148
rect 18141 3145 18153 3148
rect 18187 3145 18199 3179
rect 18141 3139 18199 3145
rect 18322 3136 18328 3188
rect 18380 3176 18386 3188
rect 23201 3179 23259 3185
rect 23201 3176 23213 3179
rect 18380 3148 23213 3176
rect 18380 3136 18386 3148
rect 23201 3145 23213 3148
rect 23247 3145 23259 3179
rect 23934 3176 23940 3188
rect 23895 3148 23940 3176
rect 23201 3139 23259 3145
rect 23934 3136 23940 3148
rect 23992 3136 23998 3188
rect 35710 3136 35716 3188
rect 35768 3176 35774 3188
rect 36725 3179 36783 3185
rect 36725 3176 36737 3179
rect 35768 3148 36737 3176
rect 35768 3136 35774 3148
rect 36725 3145 36737 3148
rect 36771 3145 36783 3179
rect 36725 3139 36783 3145
rect 8212 3111 8270 3117
rect 8212 3077 8224 3111
rect 8258 3077 8270 3111
rect 10226 3108 10232 3120
rect 9430 3080 10232 3108
rect 8212 3071 8270 3077
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 10505 3111 10563 3117
rect 10505 3108 10517 3111
rect 10336 3080 10517 3108
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 4120 3012 4169 3040
rect 4120 3000 4126 3012
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 4157 3003 4215 3009
rect 5644 3012 6653 3040
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 1360 2944 1593 2972
rect 1360 2932 1366 2944
rect 1581 2941 1593 2944
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 3418 2972 3424 2984
rect 1903 2944 3424 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 5644 2972 5672 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 5902 2972 5908 2984
rect 3568 2944 5672 2972
rect 5863 2944 5908 2972
rect 3568 2932 3574 2944
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 6656 2972 6684 3003
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 7929 3043 7987 3049
rect 7929 3040 7941 3043
rect 7524 3012 7941 3040
rect 7524 3000 7530 3012
rect 7929 3009 7941 3012
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 10336 3040 10364 3080
rect 10505 3077 10517 3080
rect 10551 3077 10563 3111
rect 10505 3071 10563 3077
rect 10597 3111 10655 3117
rect 10597 3077 10609 3111
rect 10643 3108 10655 3111
rect 10686 3108 10692 3120
rect 10643 3080 10692 3108
rect 10643 3077 10655 3080
rect 10597 3071 10655 3077
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 11514 3068 11520 3120
rect 11572 3108 11578 3120
rect 11977 3111 12035 3117
rect 11977 3108 11989 3111
rect 11572 3080 11989 3108
rect 11572 3068 11578 3080
rect 11977 3077 11989 3080
rect 12023 3077 12035 3111
rect 11977 3071 12035 3077
rect 13262 3068 13268 3120
rect 13320 3108 13326 3120
rect 14366 3108 14372 3120
rect 13320 3080 14372 3108
rect 13320 3068 13326 3080
rect 14366 3068 14372 3080
rect 14424 3068 14430 3120
rect 17954 3108 17960 3120
rect 15502 3080 17960 3108
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 11698 3040 11704 3052
rect 10192 3012 10364 3040
rect 11659 3012 11704 3040
rect 10192 3000 10198 3012
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 13078 3000 13084 3052
rect 13136 3000 13142 3052
rect 16666 3000 16672 3052
rect 16724 3040 16730 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16724 3012 17049 3040
rect 16724 3000 16730 3012
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 9950 2972 9956 2984
rect 6656 2944 9260 2972
rect 9863 2944 9956 2972
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2904 3387 2907
rect 4154 2904 4160 2916
rect 3375 2876 4160 2904
rect 3375 2873 3387 2876
rect 3329 2867 3387 2873
rect 4154 2864 4160 2876
rect 4212 2864 4218 2916
rect 9232 2904 9260 2944
rect 9950 2932 9956 2944
rect 10008 2972 10014 2984
rect 10502 2972 10508 2984
rect 10008 2944 10508 2972
rect 10008 2932 10014 2944
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 13722 2972 13728 2984
rect 11195 2944 13728 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 13998 2981 14004 2984
rect 13990 2975 14004 2981
rect 13990 2941 14002 2975
rect 14056 2972 14062 2984
rect 14056 2944 14090 2972
rect 13990 2935 14004 2941
rect 13998 2932 14004 2935
rect 14056 2932 14062 2944
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 17696 2972 17724 3003
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18785 3043 18843 3049
rect 18785 3040 18797 3043
rect 17920 3012 18797 3040
rect 17920 3000 17926 3012
rect 18785 3009 18797 3012
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 19392 3012 19441 3040
rect 19392 3000 19398 3012
rect 19429 3009 19441 3012
rect 19475 3040 19487 3043
rect 20073 3043 20131 3049
rect 20073 3040 20085 3043
rect 19475 3012 20085 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 20073 3009 20085 3012
rect 20119 3040 20131 3043
rect 20717 3043 20775 3049
rect 20717 3040 20729 3043
rect 20119 3012 20729 3040
rect 20119 3009 20131 3012
rect 20073 3003 20131 3009
rect 20717 3009 20729 3012
rect 20763 3040 20775 3043
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 20763 3012 22017 3040
rect 20763 3009 20775 3012
rect 20717 3003 20775 3009
rect 22005 3009 22017 3012
rect 22051 3040 22063 3043
rect 22649 3043 22707 3049
rect 22649 3040 22661 3043
rect 22051 3012 22661 3040
rect 22051 3009 22063 3012
rect 22005 3003 22063 3009
rect 22649 3009 22661 3012
rect 22695 3009 22707 3043
rect 23106 3040 23112 3052
rect 23067 3012 23112 3040
rect 22649 3003 22707 3009
rect 23106 3000 23112 3012
rect 23164 3000 23170 3052
rect 23566 3000 23572 3052
rect 23624 3040 23630 3052
rect 23661 3043 23719 3049
rect 23661 3040 23673 3043
rect 23624 3012 23673 3040
rect 23624 3000 23630 3012
rect 23661 3009 23673 3012
rect 23707 3040 23719 3043
rect 24121 3043 24179 3049
rect 24121 3040 24133 3043
rect 23707 3012 24133 3040
rect 23707 3009 23719 3012
rect 23661 3003 23719 3009
rect 24121 3009 24133 3012
rect 24167 3009 24179 3043
rect 24121 3003 24179 3009
rect 36909 3043 36967 3049
rect 36909 3009 36921 3043
rect 36955 3040 36967 3043
rect 37274 3040 37280 3052
rect 36955 3012 37280 3040
rect 36955 3009 36967 3012
rect 36909 3003 36967 3009
rect 37274 3000 37280 3012
rect 37332 3000 37338 3052
rect 38010 3040 38016 3052
rect 37971 3012 38016 3040
rect 38010 3000 38016 3012
rect 38068 3000 38074 3052
rect 14424 2944 17724 2972
rect 14424 2932 14430 2944
rect 11606 2904 11612 2916
rect 9232 2876 11612 2904
rect 11606 2864 11612 2876
rect 11664 2864 11670 2916
rect 15746 2904 15752 2916
rect 15707 2876 15752 2904
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 15838 2864 15844 2916
rect 15896 2864 15902 2916
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 18598 2904 18604 2916
rect 16899 2876 18604 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 22186 2864 22192 2916
rect 22244 2904 22250 2916
rect 22741 2907 22799 2913
rect 22741 2904 22753 2907
rect 22244 2876 22753 2904
rect 22244 2864 22250 2876
rect 22741 2873 22753 2876
rect 22787 2873 22799 2907
rect 22741 2867 22799 2873
rect 4420 2839 4478 2845
rect 4420 2805 4432 2839
rect 4466 2836 4478 2839
rect 7650 2836 7656 2848
rect 4466 2808 7656 2836
rect 4466 2805 4478 2808
rect 4420 2799 4478 2805
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 13630 2836 13636 2848
rect 10192 2808 13636 2836
rect 10192 2796 10198 2808
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 13814 2796 13820 2848
rect 13872 2836 13878 2848
rect 14258 2839 14316 2845
rect 14258 2836 14270 2839
rect 13872 2808 14270 2836
rect 13872 2796 13878 2808
rect 14258 2805 14270 2808
rect 14304 2805 14316 2839
rect 15856 2836 15884 2864
rect 17497 2839 17555 2845
rect 17497 2836 17509 2839
rect 15856 2808 17509 2836
rect 14258 2799 14316 2805
rect 17497 2805 17509 2808
rect 17543 2805 17555 2839
rect 18874 2836 18880 2848
rect 18835 2808 18880 2836
rect 17497 2799 17555 2805
rect 18874 2796 18880 2808
rect 18932 2796 18938 2848
rect 18966 2796 18972 2848
rect 19024 2836 19030 2848
rect 19521 2839 19579 2845
rect 19521 2836 19533 2839
rect 19024 2808 19533 2836
rect 19024 2796 19030 2808
rect 19521 2805 19533 2808
rect 19567 2805 19579 2839
rect 20162 2836 20168 2848
rect 20123 2808 20168 2836
rect 19521 2799 19579 2805
rect 20162 2796 20168 2808
rect 20220 2796 20226 2848
rect 20714 2796 20720 2848
rect 20772 2836 20778 2848
rect 20809 2839 20867 2845
rect 20809 2836 20821 2839
rect 20772 2808 20821 2836
rect 20772 2796 20778 2808
rect 20809 2805 20821 2808
rect 20855 2805 20867 2839
rect 20809 2799 20867 2805
rect 22094 2796 22100 2848
rect 22152 2836 22158 2848
rect 38194 2836 38200 2848
rect 22152 2808 22197 2836
rect 38155 2808 38200 2836
rect 22152 2796 22158 2808
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 3418 2632 3424 2644
rect 3331 2604 3424 2632
rect 3418 2592 3424 2604
rect 3476 2632 3482 2644
rect 4982 2632 4988 2644
rect 3476 2604 4988 2632
rect 3476 2592 3482 2604
rect 4982 2592 4988 2604
rect 5040 2592 5046 2644
rect 9766 2592 9772 2644
rect 9824 2632 9830 2644
rect 11057 2635 11115 2641
rect 9824 2604 10640 2632
rect 9824 2592 9830 2604
rect 4062 2564 4068 2576
rect 2976 2536 4068 2564
rect 2976 2496 3004 2536
rect 4062 2524 4068 2536
rect 4120 2564 4126 2576
rect 4120 2536 4200 2564
rect 4120 2524 4126 2536
rect 4172 2505 4200 2536
rect 5902 2524 5908 2576
rect 5960 2564 5966 2576
rect 10612 2564 10640 2604
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 11146 2632 11152 2644
rect 11103 2604 11152 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11256 2604 14412 2632
rect 11256 2564 11284 2604
rect 5960 2536 6684 2564
rect 10612 2536 11284 2564
rect 5960 2524 5966 2536
rect 1688 2468 3004 2496
rect 4157 2499 4215 2505
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1688 2437 1716 2468
rect 4157 2465 4169 2499
rect 4203 2465 4215 2499
rect 4157 2459 4215 2465
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6549 2499 6607 2505
rect 6549 2496 6561 2499
rect 6052 2468 6561 2496
rect 6052 2456 6058 2468
rect 6549 2465 6561 2468
rect 6595 2465 6607 2499
rect 6656 2496 6684 2536
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 6656 2468 6837 2496
rect 6549 2459 6607 2465
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 9306 2496 9312 2508
rect 7524 2468 9312 2496
rect 7524 2456 7530 2468
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 11698 2496 11704 2508
rect 11659 2468 11704 2496
rect 11698 2456 11704 2468
rect 11756 2496 11762 2508
rect 14274 2496 14280 2508
rect 11756 2468 14280 2496
rect 11756 2456 11762 2468
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 14384 2496 14412 2604
rect 14642 2592 14648 2644
rect 14700 2632 14706 2644
rect 14700 2604 15792 2632
rect 14700 2592 14706 2604
rect 15764 2564 15792 2604
rect 16758 2592 16764 2644
rect 16816 2632 16822 2644
rect 17497 2635 17555 2641
rect 17497 2632 17509 2635
rect 16816 2604 17509 2632
rect 16816 2592 16822 2604
rect 17497 2601 17509 2604
rect 17543 2601 17555 2635
rect 17497 2595 17555 2601
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 20162 2632 20168 2644
rect 19392 2604 20168 2632
rect 19392 2592 19398 2604
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 20254 2592 20260 2644
rect 20312 2632 20318 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 20312 2604 22017 2632
rect 20312 2592 20318 2604
rect 22005 2601 22017 2604
rect 22051 2601 22063 2635
rect 22005 2595 22063 2601
rect 24210 2592 24216 2644
rect 24268 2632 24274 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 24268 2604 27169 2632
rect 24268 2592 24274 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27157 2595 27215 2601
rect 28442 2592 28448 2644
rect 28500 2632 28506 2644
rect 29733 2635 29791 2641
rect 29733 2632 29745 2635
rect 28500 2604 29745 2632
rect 28500 2592 28506 2604
rect 29733 2601 29745 2604
rect 29779 2601 29791 2635
rect 29733 2595 29791 2601
rect 30190 2592 30196 2644
rect 30248 2632 30254 2644
rect 32309 2635 32367 2641
rect 32309 2632 32321 2635
rect 30248 2604 32321 2632
rect 30248 2592 30254 2604
rect 32309 2601 32321 2604
rect 32355 2601 32367 2635
rect 32309 2595 32367 2601
rect 34698 2592 34704 2644
rect 34756 2632 34762 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 34756 2604 34897 2632
rect 34756 2592 34762 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 34885 2595 34943 2601
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 15764 2536 16865 2564
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 16853 2527 16911 2533
rect 17218 2524 17224 2576
rect 17276 2564 17282 2576
rect 22830 2564 22836 2576
rect 17276 2536 22836 2564
rect 17276 2524 17282 2536
rect 22830 2524 22836 2536
rect 22888 2524 22894 2576
rect 24578 2564 24584 2576
rect 24539 2536 24584 2564
rect 24578 2524 24584 2536
rect 24636 2524 24642 2576
rect 34422 2524 34428 2576
rect 34480 2564 34486 2576
rect 35529 2567 35587 2573
rect 35529 2564 35541 2567
rect 34480 2536 35541 2564
rect 34480 2524 34486 2536
rect 35529 2533 35541 2536
rect 35575 2533 35587 2567
rect 35529 2527 35587 2533
rect 35618 2524 35624 2576
rect 35676 2564 35682 2576
rect 36725 2567 36783 2573
rect 36725 2564 36737 2567
rect 35676 2536 36737 2564
rect 35676 2524 35682 2536
rect 36725 2533 36737 2536
rect 36771 2533 36783 2567
rect 36725 2527 36783 2533
rect 15562 2496 15568 2508
rect 14384 2468 15568 2496
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 18966 2496 18972 2508
rect 15856 2468 18972 2496
rect 1673 2431 1731 2437
rect 1673 2428 1685 2431
rect 1360 2400 1685 2428
rect 1360 2388 1366 2400
rect 1673 2397 1685 2400
rect 1719 2397 1731 2431
rect 15856 2428 15884 2468
rect 18966 2456 18972 2468
rect 19024 2456 19030 2508
rect 19426 2456 19432 2508
rect 19484 2496 19490 2508
rect 22738 2496 22744 2508
rect 19484 2468 19932 2496
rect 22699 2468 22744 2496
rect 19484 2456 19490 2468
rect 15686 2400 15884 2428
rect 1673 2391 1731 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16816 2400 17049 2428
rect 16816 2388 16822 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 18598 2428 18604 2440
rect 18559 2400 18604 2428
rect 17681 2391 17739 2397
rect 1946 2360 1952 2372
rect 1907 2332 1952 2360
rect 1946 2320 1952 2332
rect 2004 2320 2010 2372
rect 4430 2360 4436 2372
rect 3174 2332 4292 2360
rect 4391 2332 4436 2360
rect 4264 2292 4292 2332
rect 4430 2320 4436 2332
rect 4488 2320 4494 2372
rect 6822 2360 6828 2372
rect 5658 2332 6828 2360
rect 6822 2320 6828 2332
rect 6880 2320 6886 2372
rect 8478 2360 8484 2372
rect 8050 2332 8484 2360
rect 8478 2320 8484 2332
rect 8536 2320 8542 2372
rect 8570 2320 8576 2372
rect 8628 2360 8634 2372
rect 9582 2360 9588 2372
rect 8628 2332 8673 2360
rect 9543 2332 9588 2360
rect 8628 2320 8634 2332
rect 9582 2320 9588 2332
rect 9640 2320 9646 2372
rect 10042 2320 10048 2372
rect 10100 2320 10106 2372
rect 10870 2320 10876 2372
rect 10928 2360 10934 2372
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 10928 2332 11989 2360
rect 10928 2320 10934 2332
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 14458 2360 14464 2372
rect 13202 2332 14464 2360
rect 11977 2323 12035 2329
rect 14458 2320 14464 2332
rect 14516 2320 14522 2372
rect 14550 2320 14556 2372
rect 14608 2360 14614 2372
rect 14608 2332 14653 2360
rect 14608 2320 14614 2332
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17696 2360 17724 2391
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 18782 2388 18788 2440
rect 18840 2428 18846 2440
rect 19904 2437 19932 2468
rect 22738 2456 22744 2468
rect 22796 2456 22802 2508
rect 25682 2456 25688 2508
rect 25740 2496 25746 2508
rect 25740 2468 27844 2496
rect 25740 2456 25746 2468
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 18840 2400 19625 2428
rect 18840 2388 18846 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 19889 2431 19947 2437
rect 19889 2397 19901 2431
rect 19935 2397 19947 2431
rect 20993 2431 21051 2437
rect 20993 2428 21005 2431
rect 19889 2391 19947 2397
rect 20456 2400 21005 2428
rect 16172 2332 17724 2360
rect 16172 2320 16178 2332
rect 5442 2292 5448 2304
rect 4264 2264 5448 2292
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 5905 2295 5963 2301
rect 5905 2261 5917 2295
rect 5951 2292 5963 2295
rect 6914 2292 6920 2304
rect 5951 2264 6920 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 13449 2295 13507 2301
rect 13449 2292 13461 2295
rect 11020 2264 13461 2292
rect 11020 2252 11026 2264
rect 13449 2261 13461 2264
rect 13495 2261 13507 2295
rect 14568 2292 14596 2320
rect 20456 2304 20484 2400
rect 20993 2397 21005 2400
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21324 2400 22201 2428
rect 21324 2388 21330 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2428 22707 2431
rect 23106 2428 23112 2440
rect 22695 2400 23112 2428
rect 22695 2397 22707 2400
rect 22649 2391 22707 2397
rect 23106 2388 23112 2400
rect 23164 2388 23170 2440
rect 23293 2431 23351 2437
rect 23293 2397 23305 2431
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 21910 2320 21916 2372
rect 21968 2360 21974 2372
rect 23308 2360 23336 2391
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24544 2400 24777 2428
rect 24544 2388 24550 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 27816 2437 27844 2468
rect 28902 2456 28908 2508
rect 28960 2496 28966 2508
rect 28960 2468 31064 2496
rect 28960 2456 28966 2468
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 26476 2400 27353 2428
rect 26476 2388 26482 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 27801 2431 27859 2437
rect 27801 2397 27813 2431
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 31036 2437 31064 2468
rect 35802 2456 35808 2508
rect 35860 2496 35866 2508
rect 35860 2468 37504 2496
rect 35860 2456 35866 2468
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 31021 2431 31079 2437
rect 31021 2397 31033 2431
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 32272 2400 32505 2428
rect 32272 2388 32278 2400
rect 32493 2397 32505 2400
rect 32539 2397 32551 2431
rect 32493 2391 32551 2397
rect 34146 2388 34152 2440
rect 34204 2428 34210 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34204 2400 35081 2428
rect 34204 2388 34210 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35069 2391 35127 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 37476 2437 37504 2468
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 36909 2431 36967 2437
rect 36909 2397 36921 2431
rect 36955 2397 36967 2431
rect 36909 2391 36967 2397
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 21968 2332 23336 2360
rect 21968 2320 21974 2332
rect 33870 2320 33876 2372
rect 33928 2360 33934 2372
rect 35618 2360 35624 2372
rect 33928 2332 35624 2360
rect 33928 2320 33934 2332
rect 35618 2320 35624 2332
rect 35676 2320 35682 2372
rect 36924 2360 36952 2391
rect 38654 2360 38660 2372
rect 36924 2332 38660 2360
rect 38654 2320 38660 2332
rect 38712 2320 38718 2372
rect 15286 2292 15292 2304
rect 14568 2264 15292 2292
rect 13449 2255 13507 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 16025 2295 16083 2301
rect 16025 2292 16037 2295
rect 15620 2264 16037 2292
rect 15620 2252 15626 2264
rect 16025 2261 16037 2264
rect 16071 2292 16083 2295
rect 18506 2292 18512 2304
rect 16071 2264 18512 2292
rect 16071 2261 16083 2264
rect 16025 2255 16083 2261
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18748 2264 18797 2292
rect 18748 2252 18754 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 19426 2292 19432 2304
rect 19387 2264 19432 2292
rect 18785 2255 18843 2261
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 20036 2264 20085 2292
rect 20036 2252 20042 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20438 2292 20444 2304
rect 20399 2264 20444 2292
rect 20073 2255 20131 2261
rect 20438 2252 20444 2264
rect 20496 2252 20502 2304
rect 20806 2292 20812 2304
rect 20767 2264 20812 2292
rect 20806 2252 20812 2264
rect 20864 2252 20870 2304
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23256 2264 23489 2292
rect 23256 2252 23262 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 27985 2295 28043 2301
rect 27985 2292 27997 2295
rect 27764 2264 27997 2292
rect 27764 2252 27770 2264
rect 27985 2261 27997 2264
rect 28031 2261 28043 2295
rect 27985 2255 28043 2261
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 30984 2264 31217 2292
rect 30984 2252 30990 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 37366 2252 37372 2304
rect 37424 2292 37430 2304
rect 37645 2295 37703 2301
rect 37645 2292 37657 2295
rect 37424 2264 37657 2292
rect 37424 2252 37430 2264
rect 37645 2261 37657 2264
rect 37691 2261 37703 2295
rect 37645 2255 37703 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 4430 2048 4436 2100
rect 4488 2088 4494 2100
rect 9950 2088 9956 2100
rect 4488 2060 9956 2088
rect 4488 2048 4494 2060
rect 9950 2048 9956 2060
rect 10008 2048 10014 2100
rect 14458 2048 14464 2100
rect 14516 2088 14522 2100
rect 17218 2088 17224 2100
rect 14516 2060 17224 2088
rect 14516 2048 14522 2060
rect 17218 2048 17224 2060
rect 17276 2048 17282 2100
rect 8478 1980 8484 2032
rect 8536 2020 8542 2032
rect 13262 2020 13268 2032
rect 8536 1992 13268 2020
rect 8536 1980 8542 1992
rect 13262 1980 13268 1992
rect 13320 1980 13326 2032
rect 13446 1980 13452 2032
rect 13504 2020 13510 2032
rect 20346 2020 20352 2032
rect 13504 1992 20352 2020
rect 13504 1980 13510 1992
rect 20346 1980 20352 1992
rect 20404 1980 20410 2032
rect 5810 1912 5816 1964
rect 5868 1952 5874 1964
rect 20438 1952 20444 1964
rect 5868 1924 20444 1952
rect 5868 1912 5874 1924
rect 20438 1912 20444 1924
rect 20496 1912 20502 1964
rect 11606 1844 11612 1896
rect 11664 1884 11670 1896
rect 20806 1884 20812 1896
rect 11664 1856 20812 1884
rect 11664 1844 11670 1856
rect 20806 1844 20812 1856
rect 20864 1844 20870 1896
rect 8294 1776 8300 1828
rect 8352 1816 8358 1828
rect 19334 1816 19340 1828
rect 8352 1788 19340 1816
rect 8352 1776 8358 1788
rect 19334 1776 19340 1788
rect 19392 1776 19398 1828
rect 12250 1708 12256 1760
rect 12308 1748 12314 1760
rect 18782 1748 18788 1760
rect 12308 1720 18788 1748
rect 12308 1708 12314 1720
rect 18782 1708 18788 1720
rect 18840 1708 18846 1760
rect 9582 1640 9588 1692
rect 9640 1680 9646 1692
rect 15654 1680 15660 1692
rect 9640 1652 15660 1680
rect 9640 1640 9646 1652
rect 15654 1640 15660 1652
rect 15712 1640 15718 1692
rect 5534 1572 5540 1624
rect 5592 1612 5598 1624
rect 5592 1584 13124 1612
rect 5592 1572 5598 1584
rect 13096 1476 13124 1584
rect 13262 1572 13268 1624
rect 13320 1612 13326 1624
rect 20714 1612 20720 1624
rect 13320 1584 20720 1612
rect 13320 1572 13326 1584
rect 20714 1572 20720 1584
rect 20772 1572 20778 1624
rect 20530 1476 20536 1488
rect 13096 1448 20536 1476
rect 20530 1436 20536 1448
rect 20588 1436 20594 1488
rect 8570 1368 8576 1420
rect 8628 1408 8634 1420
rect 14550 1408 14556 1420
rect 8628 1380 14556 1408
rect 8628 1368 8634 1380
rect 14550 1368 14556 1380
rect 14608 1368 14614 1420
rect 15470 1368 15476 1420
rect 15528 1408 15534 1420
rect 16114 1408 16120 1420
rect 15528 1380 16120 1408
rect 15528 1368 15534 1380
rect 16114 1368 16120 1380
rect 16172 1368 16178 1420
rect 14 1300 20 1352
rect 72 1340 78 1352
rect 4706 1340 4712 1352
rect 72 1312 4712 1340
rect 72 1300 78 1312
rect 4706 1300 4712 1312
rect 4764 1300 4770 1352
rect 20070 1340 20076 1352
rect 4816 1312 20076 1340
rect 3786 1232 3792 1284
rect 3844 1272 3850 1284
rect 4816 1272 4844 1312
rect 20070 1300 20076 1312
rect 20128 1300 20134 1352
rect 18874 1272 18880 1284
rect 3844 1244 4844 1272
rect 4908 1244 18880 1272
rect 3844 1232 3850 1244
rect 3970 1096 3976 1148
rect 4028 1136 4034 1148
rect 4908 1136 4936 1244
rect 18874 1232 18880 1244
rect 18932 1232 18938 1284
rect 4982 1164 4988 1216
rect 5040 1204 5046 1216
rect 20622 1204 20628 1216
rect 5040 1176 20628 1204
rect 5040 1164 5046 1176
rect 20622 1164 20628 1176
rect 20680 1164 20686 1216
rect 4028 1108 4936 1136
rect 4028 1096 4034 1108
rect 7558 1096 7564 1148
rect 7616 1136 7622 1148
rect 22370 1136 22376 1148
rect 7616 1108 22376 1136
rect 7616 1096 7622 1108
rect 22370 1096 22376 1108
rect 22428 1096 22434 1148
rect 5258 1028 5264 1080
rect 5316 1068 5322 1080
rect 19150 1068 19156 1080
rect 5316 1040 19156 1068
rect 5316 1028 5322 1040
rect 19150 1028 19156 1040
rect 19208 1028 19214 1080
rect 6638 960 6644 1012
rect 6696 1000 6702 1012
rect 20254 1000 20260 1012
rect 6696 972 20260 1000
rect 6696 960 6702 972
rect 20254 960 20260 972
rect 20312 960 20318 1012
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 7104 37272 7156 37324
rect 1860 37204 1912 37256
rect 1952 37204 2004 37256
rect 3148 37247 3200 37256
rect 3148 37213 3157 37247
rect 3157 37213 3191 37247
rect 3191 37213 3200 37247
rect 3148 37204 3200 37213
rect 3976 37247 4028 37256
rect 3976 37213 3985 37247
rect 3985 37213 4019 37247
rect 4019 37213 4028 37247
rect 3976 37204 4028 37213
rect 6736 37204 6788 37256
rect 7472 37247 7524 37256
rect 7472 37213 7481 37247
rect 7481 37213 7515 37247
rect 7515 37213 7524 37247
rect 7472 37204 7524 37213
rect 8392 37204 8444 37256
rect 10324 37204 10376 37256
rect 11612 37204 11664 37256
rect 12900 37204 12952 37256
rect 14924 37247 14976 37256
rect 14924 37213 14933 37247
rect 14933 37213 14967 37247
rect 14967 37213 14976 37247
rect 14924 37204 14976 37213
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 18144 37247 18196 37256
rect 18144 37213 18153 37247
rect 18153 37213 18187 37247
rect 18187 37213 18196 37247
rect 18144 37204 18196 37213
rect 19432 37247 19484 37256
rect 19432 37213 19441 37247
rect 19441 37213 19475 37247
rect 19475 37213 19484 37247
rect 19432 37204 19484 37213
rect 20720 37204 20772 37256
rect 22560 37204 22612 37256
rect 22928 37204 22980 37256
rect 24676 37204 24728 37256
rect 27068 37204 27120 37256
rect 27804 37204 27856 37256
rect 30380 37204 30432 37256
rect 31760 37204 31812 37256
rect 33508 37204 33560 37256
rect 34796 37204 34848 37256
rect 36728 37204 36780 37256
rect 2780 37136 2832 37188
rect 2872 37068 2924 37120
rect 6552 37136 6604 37188
rect 3884 37068 3936 37120
rect 5172 37068 5224 37120
rect 9128 37111 9180 37120
rect 9128 37077 9137 37111
rect 9137 37077 9171 37111
rect 9171 37077 9180 37111
rect 9128 37068 9180 37077
rect 11980 37136 12032 37188
rect 31852 37136 31904 37188
rect 10784 37068 10836 37120
rect 12992 37111 13044 37120
rect 12992 37077 13001 37111
rect 13001 37077 13035 37111
rect 13035 37077 13044 37111
rect 12992 37068 13044 37077
rect 14832 37068 14884 37120
rect 16580 37068 16632 37120
rect 18052 37068 18104 37120
rect 19340 37068 19392 37120
rect 20720 37111 20772 37120
rect 20720 37077 20729 37111
rect 20729 37077 20763 37111
rect 20763 37077 20772 37111
rect 20720 37068 20772 37077
rect 21732 37068 21784 37120
rect 23848 37068 23900 37120
rect 25780 37068 25832 37120
rect 27160 37111 27212 37120
rect 27160 37077 27169 37111
rect 27169 37077 27203 37111
rect 27203 37077 27212 37111
rect 27160 37068 27212 37077
rect 29000 37068 29052 37120
rect 30012 37068 30064 37120
rect 32312 37111 32364 37120
rect 32312 37077 32321 37111
rect 32321 37077 32355 37111
rect 32355 37077 32364 37111
rect 32312 37068 32364 37077
rect 33600 37111 33652 37120
rect 33600 37077 33609 37111
rect 33609 37077 33643 37111
rect 33643 37077 33652 37111
rect 33600 37068 33652 37077
rect 35532 37136 35584 37188
rect 35900 37068 35952 37120
rect 38200 37111 38252 37120
rect 38200 37077 38209 37111
rect 38209 37077 38243 37111
rect 38243 37077 38252 37111
rect 38200 37068 38252 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 664 36864 716 36916
rect 1860 36864 1912 36916
rect 2872 36864 2924 36916
rect 5448 36864 5500 36916
rect 29736 36864 29788 36916
rect 33600 36864 33652 36916
rect 38292 36864 38344 36916
rect 2504 36771 2556 36780
rect 2504 36737 2513 36771
rect 2513 36737 2547 36771
rect 2547 36737 2556 36771
rect 2504 36728 2556 36737
rect 39304 36796 39356 36848
rect 4068 36660 4120 36712
rect 35348 36660 35400 36712
rect 36728 36567 36780 36576
rect 36728 36533 36737 36567
rect 36737 36533 36771 36567
rect 36771 36533 36780 36567
rect 36728 36524 36780 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1768 36159 1820 36168
rect 1768 36125 1777 36159
rect 1777 36125 1811 36159
rect 1811 36125 1820 36159
rect 1768 36116 1820 36125
rect 38016 36116 38068 36168
rect 2688 35980 2740 36032
rect 34520 35980 34572 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 2504 35819 2556 35828
rect 2504 35785 2513 35819
rect 2513 35785 2547 35819
rect 2547 35785 2556 35819
rect 2504 35776 2556 35785
rect 2412 35683 2464 35692
rect 2412 35649 2421 35683
rect 2421 35649 2455 35683
rect 2455 35649 2464 35683
rect 2412 35640 2464 35649
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4068 35232 4120 35284
rect 14924 35232 14976 35284
rect 16856 35232 16908 35284
rect 18144 35232 18196 35284
rect 22928 35232 22980 35284
rect 24676 35232 24728 35284
rect 7196 35028 7248 35080
rect 12992 35028 13044 35080
rect 15660 35028 15712 35080
rect 16672 35071 16724 35080
rect 16672 35037 16681 35071
rect 16681 35037 16715 35071
rect 16715 35037 16724 35071
rect 16672 35028 16724 35037
rect 17592 35071 17644 35080
rect 17592 35037 17601 35071
rect 17601 35037 17635 35071
rect 17635 35037 17644 35071
rect 17592 35028 17644 35037
rect 19984 35028 20036 35080
rect 22008 35028 22060 35080
rect 31852 35028 31904 35080
rect 35440 35028 35492 35080
rect 11704 34892 11756 34944
rect 30564 34935 30616 34944
rect 30564 34901 30573 34935
rect 30573 34901 30607 34935
rect 30607 34901 30616 34935
rect 30564 34892 30616 34901
rect 38200 34935 38252 34944
rect 38200 34901 38209 34935
rect 38209 34901 38243 34935
rect 38243 34901 38252 34935
rect 38200 34892 38252 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 6736 34688 6788 34740
rect 19432 34688 19484 34740
rect 27804 34688 27856 34740
rect 4068 34552 4120 34604
rect 9864 34552 9916 34604
rect 11980 34595 12032 34604
rect 11980 34561 11989 34595
rect 11989 34561 12023 34595
rect 12023 34561 12032 34595
rect 11980 34552 12032 34561
rect 18512 34595 18564 34604
rect 18512 34561 18521 34595
rect 18521 34561 18555 34595
rect 18555 34561 18564 34595
rect 18512 34552 18564 34561
rect 20720 34552 20772 34604
rect 27344 34595 27396 34604
rect 27344 34561 27353 34595
rect 27353 34561 27387 34595
rect 27387 34561 27396 34595
rect 27344 34552 27396 34561
rect 34520 34552 34572 34604
rect 12164 34484 12216 34536
rect 19064 34484 19116 34536
rect 33324 34527 33376 34536
rect 33324 34493 33333 34527
rect 33333 34493 33367 34527
rect 33367 34493 33376 34527
rect 33324 34484 33376 34493
rect 1768 34391 1820 34400
rect 1768 34357 1777 34391
rect 1777 34357 1811 34391
rect 1811 34357 1820 34391
rect 1768 34348 1820 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 7196 34187 7248 34196
rect 7196 34153 7205 34187
rect 7205 34153 7239 34187
rect 7239 34153 7248 34187
rect 7196 34144 7248 34153
rect 27344 34144 27396 34196
rect 35348 34144 35400 34196
rect 7104 33983 7156 33992
rect 7104 33949 7113 33983
rect 7113 33949 7147 33983
rect 7147 33949 7156 33983
rect 7104 33940 7156 33949
rect 21732 33983 21784 33992
rect 21732 33949 21741 33983
rect 21741 33949 21775 33983
rect 21775 33949 21784 33983
rect 21732 33940 21784 33949
rect 23204 33940 23256 33992
rect 29736 33983 29788 33992
rect 29736 33949 29745 33983
rect 29745 33949 29779 33983
rect 29779 33949 29788 33983
rect 29736 33940 29788 33949
rect 30104 33940 30156 33992
rect 21824 33847 21876 33856
rect 21824 33813 21833 33847
rect 21833 33813 21867 33847
rect 21867 33813 21876 33847
rect 21824 33804 21876 33813
rect 29828 33847 29880 33856
rect 29828 33813 29837 33847
rect 29837 33813 29871 33847
rect 29871 33813 29880 33847
rect 29828 33804 29880 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 19340 33600 19392 33652
rect 29828 33600 29880 33652
rect 10784 33507 10836 33516
rect 10784 33473 10793 33507
rect 10793 33473 10827 33507
rect 10827 33473 10836 33507
rect 10784 33464 10836 33473
rect 35348 33464 35400 33516
rect 38200 33371 38252 33380
rect 38200 33337 38209 33371
rect 38209 33337 38243 33371
rect 38243 33337 38252 33371
rect 38200 33328 38252 33337
rect 10140 33260 10192 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1768 32895 1820 32904
rect 1768 32861 1777 32895
rect 1777 32861 1811 32895
rect 1811 32861 1820 32895
rect 1768 32852 1820 32861
rect 5540 32716 5592 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 35532 32512 35584 32564
rect 6552 32419 6604 32428
rect 6552 32385 6561 32419
rect 6561 32385 6595 32419
rect 6595 32385 6604 32419
rect 6552 32376 6604 32385
rect 7104 32376 7156 32428
rect 20168 32376 20220 32428
rect 27160 32376 27212 32428
rect 29920 32376 29972 32428
rect 29000 32308 29052 32360
rect 30012 32308 30064 32360
rect 6644 32215 6696 32224
rect 6644 32181 6653 32215
rect 6653 32181 6687 32215
rect 6687 32181 6696 32215
rect 6644 32172 6696 32181
rect 18788 32172 18840 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 9864 32011 9916 32020
rect 9864 31977 9873 32011
rect 9873 31977 9907 32011
rect 9907 31977 9916 32011
rect 9864 31968 9916 31977
rect 18420 31900 18472 31952
rect 5448 31764 5500 31816
rect 8852 31764 8904 31816
rect 9128 31807 9180 31816
rect 9128 31773 9137 31807
rect 9137 31773 9171 31807
rect 9171 31773 9180 31807
rect 9128 31764 9180 31773
rect 9312 31764 9364 31816
rect 10876 31764 10928 31816
rect 29000 31832 29052 31884
rect 25228 31807 25280 31816
rect 25228 31773 25237 31807
rect 25237 31773 25271 31807
rect 25271 31773 25280 31807
rect 25228 31764 25280 31773
rect 32312 31968 32364 32020
rect 37004 31900 37056 31952
rect 29828 31875 29880 31884
rect 29828 31841 29837 31875
rect 29837 31841 29871 31875
rect 29871 31841 29880 31875
rect 29828 31832 29880 31841
rect 35900 31764 35952 31816
rect 38292 31807 38344 31816
rect 38292 31773 38301 31807
rect 38301 31773 38335 31807
rect 38335 31773 38344 31807
rect 38292 31764 38344 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 36728 31288 36780 31340
rect 20444 31084 20496 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 4068 30880 4120 30932
rect 16672 30880 16724 30932
rect 35440 30880 35492 30932
rect 1768 30719 1820 30728
rect 1768 30685 1777 30719
rect 1777 30685 1811 30719
rect 1811 30685 1820 30719
rect 1768 30676 1820 30685
rect 6092 30676 6144 30728
rect 17408 30676 17460 30728
rect 30012 30676 30064 30728
rect 3792 30540 3844 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 15660 30311 15712 30320
rect 15660 30277 15669 30311
rect 15669 30277 15703 30311
rect 15703 30277 15712 30311
rect 15660 30268 15712 30277
rect 16028 30200 16080 30252
rect 38292 30243 38344 30252
rect 38292 30209 38301 30243
rect 38301 30209 38335 30243
rect 38335 30209 38344 30243
rect 38292 30200 38344 30209
rect 34152 29996 34204 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 6092 29835 6144 29844
rect 6092 29801 6101 29835
rect 6101 29801 6135 29835
rect 6135 29801 6144 29835
rect 6092 29792 6144 29801
rect 17592 29792 17644 29844
rect 19984 29792 20036 29844
rect 22008 29835 22060 29844
rect 22008 29801 22017 29835
rect 22017 29801 22051 29835
rect 22051 29801 22060 29835
rect 22008 29792 22060 29801
rect 35348 29792 35400 29844
rect 2688 29588 2740 29640
rect 7656 29588 7708 29640
rect 17592 29588 17644 29640
rect 2780 29520 2832 29572
rect 16764 29520 16816 29572
rect 20628 29588 20680 29640
rect 34704 29588 34756 29640
rect 1768 29495 1820 29504
rect 1768 29461 1777 29495
rect 1777 29461 1811 29495
rect 1811 29461 1820 29495
rect 1768 29452 1820 29461
rect 4068 29495 4120 29504
rect 4068 29461 4077 29495
rect 4077 29461 4111 29495
rect 4111 29461 4120 29495
rect 4068 29452 4120 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 18512 29248 18564 29300
rect 30104 29248 30156 29300
rect 17960 29155 18012 29164
rect 17960 29121 17969 29155
rect 17969 29121 18003 29155
rect 18003 29121 18012 29155
rect 17960 29112 18012 29121
rect 29092 29155 29144 29164
rect 29092 29121 29101 29155
rect 29101 29121 29135 29155
rect 29135 29121 29144 29155
rect 29092 29112 29144 29121
rect 38016 29155 38068 29164
rect 38016 29121 38025 29155
rect 38025 29121 38059 29155
rect 38059 29121 38068 29155
rect 38016 29112 38068 29121
rect 2780 28976 2832 29028
rect 38200 29019 38252 29028
rect 38200 28985 38209 29019
rect 38209 28985 38243 29019
rect 38243 28985 38252 29019
rect 38200 28976 38252 28985
rect 4068 28908 4120 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 29920 28704 29972 28756
rect 5540 28500 5592 28552
rect 29736 28543 29788 28552
rect 29736 28509 29745 28543
rect 29745 28509 29779 28543
rect 29779 28509 29788 28543
rect 29736 28500 29788 28509
rect 7012 28407 7064 28416
rect 7012 28373 7021 28407
rect 7021 28373 7055 28407
rect 7055 28373 7064 28407
rect 7012 28364 7064 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 1768 28067 1820 28076
rect 1768 28033 1777 28067
rect 1777 28033 1811 28067
rect 1811 28033 1820 28067
rect 1768 28024 1820 28033
rect 37004 28024 37056 28076
rect 3884 27820 3936 27872
rect 32404 27863 32456 27872
rect 32404 27829 32413 27863
rect 32413 27829 32447 27863
rect 32447 27829 32456 27863
rect 32404 27820 32456 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3792 27412 3844 27464
rect 34152 27455 34204 27464
rect 34152 27421 34161 27455
rect 34161 27421 34195 27455
rect 34195 27421 34204 27455
rect 34152 27412 34204 27421
rect 8576 27276 8628 27328
rect 20720 27276 20772 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 34796 26936 34848 26988
rect 38200 26775 38252 26784
rect 38200 26741 38209 26775
rect 38209 26741 38243 26775
rect 38243 26741 38252 26775
rect 38200 26732 38252 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 30012 26528 30064 26580
rect 5080 26460 5132 26512
rect 1768 26367 1820 26376
rect 1768 26333 1777 26367
rect 1777 26333 1811 26367
rect 1811 26333 1820 26367
rect 1768 26324 1820 26333
rect 29644 26324 29696 26376
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4068 26027 4120 26036
rect 4068 25993 4077 26027
rect 4077 25993 4111 26027
rect 4111 25993 4120 26027
rect 4068 25984 4120 25993
rect 4620 25848 4672 25900
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 34704 25440 34756 25492
rect 28724 25279 28776 25288
rect 28724 25245 28733 25279
rect 28733 25245 28767 25279
rect 28767 25245 28776 25279
rect 28724 25236 28776 25245
rect 38292 25279 38344 25288
rect 38292 25245 38301 25279
rect 38301 25245 38335 25279
rect 38335 25245 38344 25279
rect 38292 25236 38344 25245
rect 34612 25100 34664 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 5448 24760 5500 24812
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 32036 24760 32088 24812
rect 17132 24735 17184 24744
rect 17132 24701 17141 24735
rect 17141 24701 17175 24735
rect 17175 24701 17184 24735
rect 17132 24692 17184 24701
rect 18144 24692 18196 24744
rect 19984 24692 20036 24744
rect 38016 24624 38068 24676
rect 1768 24599 1820 24608
rect 1768 24565 1777 24599
rect 1777 24565 1811 24599
rect 1811 24565 1820 24599
rect 1768 24556 1820 24565
rect 19432 24599 19484 24608
rect 19432 24565 19441 24599
rect 19441 24565 19475 24599
rect 19475 24565 19484 24599
rect 19432 24556 19484 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 18144 24395 18196 24404
rect 18144 24361 18153 24395
rect 18153 24361 18187 24395
rect 18187 24361 18196 24395
rect 18144 24352 18196 24361
rect 19984 24259 20036 24268
rect 19984 24225 19993 24259
rect 19993 24225 20027 24259
rect 20027 24225 20036 24259
rect 19984 24216 20036 24225
rect 20628 24259 20680 24268
rect 20628 24225 20637 24259
rect 20637 24225 20671 24259
rect 20671 24225 20680 24259
rect 20628 24216 20680 24225
rect 16120 24148 16172 24200
rect 16948 24148 17000 24200
rect 18052 24191 18104 24200
rect 18052 24157 18061 24191
rect 18061 24157 18095 24191
rect 18095 24157 18104 24191
rect 18052 24148 18104 24157
rect 18328 24148 18380 24200
rect 17224 24012 17276 24064
rect 17500 24012 17552 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 16120 23851 16172 23860
rect 16120 23817 16129 23851
rect 16129 23817 16163 23851
rect 16163 23817 16172 23851
rect 16120 23808 16172 23817
rect 18328 23851 18380 23860
rect 18328 23817 18337 23851
rect 18337 23817 18371 23851
rect 18371 23817 18380 23851
rect 18328 23808 18380 23817
rect 34796 23851 34848 23860
rect 34796 23817 34805 23851
rect 34805 23817 34839 23851
rect 34839 23817 34848 23851
rect 34796 23808 34848 23817
rect 17132 23783 17184 23792
rect 17132 23749 17141 23783
rect 17141 23749 17175 23783
rect 17175 23749 17184 23783
rect 17132 23740 17184 23749
rect 17224 23783 17276 23792
rect 17224 23749 17233 23783
rect 17233 23749 17267 23783
rect 17267 23749 17276 23783
rect 17224 23740 17276 23749
rect 20628 23740 20680 23792
rect 3884 23672 3936 23724
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 9496 23604 9548 23656
rect 16948 23672 17000 23724
rect 18512 23715 18564 23724
rect 18512 23681 18521 23715
rect 18521 23681 18555 23715
rect 18555 23681 18564 23715
rect 18512 23672 18564 23681
rect 31760 23672 31812 23724
rect 38292 23715 38344 23724
rect 38292 23681 38301 23715
rect 38301 23681 38335 23715
rect 38335 23681 38344 23715
rect 38292 23672 38344 23681
rect 17408 23647 17460 23656
rect 17408 23613 17417 23647
rect 17417 23613 17451 23647
rect 17451 23613 17460 23647
rect 17408 23604 17460 23613
rect 19432 23604 19484 23656
rect 9588 23468 9640 23520
rect 12900 23468 12952 23520
rect 15200 23468 15252 23520
rect 34520 23468 34572 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 9220 23128 9272 23180
rect 18052 23264 18104 23316
rect 19432 23264 19484 23316
rect 17408 23196 17460 23248
rect 21088 23239 21140 23248
rect 12900 23103 12952 23112
rect 12900 23069 12909 23103
rect 12909 23069 12943 23103
rect 12943 23069 12952 23103
rect 12900 23060 12952 23069
rect 13360 23103 13412 23112
rect 13360 23069 13369 23103
rect 13369 23069 13403 23103
rect 13403 23069 13412 23103
rect 13360 23060 13412 23069
rect 14556 23103 14608 23112
rect 14556 23069 14565 23103
rect 14565 23069 14599 23103
rect 14599 23069 14608 23103
rect 14556 23060 14608 23069
rect 15200 23103 15252 23112
rect 15200 23069 15209 23103
rect 15209 23069 15243 23103
rect 15243 23069 15252 23103
rect 15200 23060 15252 23069
rect 15844 23103 15896 23112
rect 15844 23069 15853 23103
rect 15853 23069 15887 23103
rect 15887 23069 15896 23103
rect 15844 23060 15896 23069
rect 13176 22992 13228 23044
rect 14004 22992 14056 23044
rect 21088 23205 21097 23239
rect 21097 23205 21131 23239
rect 21131 23205 21140 23239
rect 21088 23196 21140 23205
rect 20720 23171 20772 23180
rect 20720 23137 20729 23171
rect 20729 23137 20763 23171
rect 20763 23137 20772 23171
rect 20720 23128 20772 23137
rect 20904 23103 20956 23112
rect 17500 23035 17552 23044
rect 17500 23001 17509 23035
rect 17509 23001 17543 23035
rect 17543 23001 17552 23035
rect 17500 22992 17552 23001
rect 12072 22967 12124 22976
rect 12072 22933 12081 22967
rect 12081 22933 12115 22967
rect 12115 22933 12124 22967
rect 12072 22924 12124 22933
rect 12716 22967 12768 22976
rect 12716 22933 12725 22967
rect 12725 22933 12759 22967
rect 12759 22933 12768 22967
rect 12716 22924 12768 22933
rect 13452 22967 13504 22976
rect 13452 22933 13461 22967
rect 13461 22933 13495 22967
rect 13495 22933 13504 22967
rect 13452 22924 13504 22933
rect 14372 22967 14424 22976
rect 14372 22933 14381 22967
rect 14381 22933 14415 22967
rect 14415 22933 14424 22967
rect 14372 22924 14424 22933
rect 15016 22967 15068 22976
rect 15016 22933 15025 22967
rect 15025 22933 15059 22967
rect 15059 22933 15068 22967
rect 15016 22924 15068 22933
rect 15660 22967 15712 22976
rect 15660 22933 15669 22967
rect 15669 22933 15703 22967
rect 15703 22933 15712 22967
rect 15660 22924 15712 22933
rect 20904 23069 20913 23103
rect 20913 23069 20947 23103
rect 20947 23069 20956 23103
rect 20904 23060 20956 23069
rect 21180 22992 21232 23044
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 5448 22763 5500 22772
rect 5448 22729 5457 22763
rect 5457 22729 5491 22763
rect 5491 22729 5500 22763
rect 5448 22720 5500 22729
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 8208 22584 8260 22636
rect 8576 22584 8628 22636
rect 12072 22627 12124 22636
rect 12072 22593 12081 22627
rect 12081 22593 12115 22627
rect 12115 22593 12124 22627
rect 12072 22584 12124 22593
rect 14556 22720 14608 22772
rect 15016 22720 15068 22772
rect 20904 22720 20956 22772
rect 21088 22763 21140 22772
rect 21088 22729 21097 22763
rect 21097 22729 21131 22763
rect 21131 22729 21140 22763
rect 21088 22720 21140 22729
rect 21180 22720 21232 22772
rect 21548 22720 21600 22772
rect 29828 22720 29880 22772
rect 17592 22695 17644 22704
rect 17592 22661 17601 22695
rect 17601 22661 17635 22695
rect 17635 22661 17644 22695
rect 17592 22652 17644 22661
rect 13728 22448 13780 22500
rect 14372 22584 14424 22636
rect 18696 22627 18748 22636
rect 18696 22593 18705 22627
rect 18705 22593 18739 22627
rect 18739 22593 18748 22627
rect 18696 22584 18748 22593
rect 19800 22627 19852 22636
rect 19800 22593 19809 22627
rect 19809 22593 19843 22627
rect 19843 22593 19852 22627
rect 19800 22584 19852 22593
rect 20444 22627 20496 22636
rect 20444 22593 20453 22627
rect 20453 22593 20487 22627
rect 20487 22593 20496 22627
rect 20444 22584 20496 22593
rect 15752 22516 15804 22568
rect 18144 22516 18196 22568
rect 18236 22516 18288 22568
rect 20628 22559 20680 22568
rect 20628 22525 20637 22559
rect 20637 22525 20671 22559
rect 20671 22525 20680 22559
rect 20628 22516 20680 22525
rect 15476 22448 15528 22500
rect 17592 22448 17644 22500
rect 5540 22380 5592 22432
rect 13268 22380 13320 22432
rect 14464 22380 14516 22432
rect 16212 22380 16264 22432
rect 18512 22423 18564 22432
rect 18512 22389 18521 22423
rect 18521 22389 18555 22423
rect 18555 22389 18564 22423
rect 18512 22380 18564 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 13268 22219 13320 22228
rect 13268 22185 13277 22219
rect 13277 22185 13311 22219
rect 13311 22185 13320 22219
rect 13268 22176 13320 22185
rect 18144 22176 18196 22228
rect 18604 22219 18656 22228
rect 18604 22185 18613 22219
rect 18613 22185 18647 22219
rect 18647 22185 18656 22219
rect 18604 22176 18656 22185
rect 20628 22176 20680 22228
rect 4620 22040 4672 22092
rect 8208 22040 8260 22092
rect 12716 22040 12768 22092
rect 13820 22108 13872 22160
rect 19800 22108 19852 22160
rect 16764 22040 16816 22092
rect 18236 22083 18288 22092
rect 18236 22049 18245 22083
rect 18245 22049 18279 22083
rect 18279 22049 18288 22083
rect 18236 22040 18288 22049
rect 18512 22040 18564 22092
rect 4804 21972 4856 22024
rect 7840 21972 7892 22024
rect 11152 22015 11204 22024
rect 11152 21981 11161 22015
rect 11161 21981 11195 22015
rect 11195 21981 11204 22015
rect 11152 21972 11204 21981
rect 11520 21972 11572 22024
rect 12256 22015 12308 22024
rect 12256 21981 12265 22015
rect 12265 21981 12299 22015
rect 12299 21981 12308 22015
rect 12256 21972 12308 21981
rect 11244 21904 11296 21956
rect 17684 21972 17736 22024
rect 31760 22040 31812 22092
rect 10324 21836 10376 21888
rect 10968 21879 11020 21888
rect 10968 21845 10977 21879
rect 10977 21845 11011 21879
rect 11011 21845 11020 21879
rect 10968 21836 11020 21845
rect 11612 21879 11664 21888
rect 11612 21845 11621 21879
rect 11621 21845 11655 21879
rect 11655 21845 11664 21879
rect 11612 21836 11664 21845
rect 14464 21947 14516 21956
rect 14464 21913 14473 21947
rect 14473 21913 14507 21947
rect 14507 21913 14516 21947
rect 16120 21947 16172 21956
rect 14464 21904 14516 21913
rect 16120 21913 16129 21947
rect 16129 21913 16163 21947
rect 16163 21913 16172 21947
rect 16120 21904 16172 21913
rect 16212 21947 16264 21956
rect 16212 21913 16221 21947
rect 16221 21913 16255 21947
rect 16255 21913 16264 21947
rect 16212 21904 16264 21913
rect 18788 21904 18840 21956
rect 18696 21836 18748 21888
rect 19432 21836 19484 21888
rect 24860 21972 24912 22024
rect 38292 22015 38344 22024
rect 38292 21981 38301 22015
rect 38301 21981 38335 22015
rect 38335 21981 38344 22015
rect 38292 21972 38344 21981
rect 38108 21879 38160 21888
rect 38108 21845 38117 21879
rect 38117 21845 38151 21879
rect 38151 21845 38160 21879
rect 38108 21836 38160 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 11152 21632 11204 21684
rect 13360 21632 13412 21684
rect 15844 21632 15896 21684
rect 18604 21632 18656 21684
rect 4896 21496 4948 21548
rect 5080 21539 5132 21548
rect 5080 21505 5089 21539
rect 5089 21505 5123 21539
rect 5123 21505 5132 21539
rect 5080 21496 5132 21505
rect 9036 21496 9088 21548
rect 10048 21496 10100 21548
rect 10508 21539 10560 21548
rect 10508 21505 10517 21539
rect 10517 21505 10551 21539
rect 10551 21505 10560 21539
rect 10508 21496 10560 21505
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 12164 21496 12216 21548
rect 13452 21496 13504 21548
rect 17684 21564 17736 21616
rect 15660 21496 15712 21548
rect 17316 21539 17368 21548
rect 17316 21505 17325 21539
rect 17325 21505 17359 21539
rect 17359 21505 17368 21539
rect 17316 21496 17368 21505
rect 8760 21471 8812 21480
rect 8760 21437 8769 21471
rect 8769 21437 8803 21471
rect 8803 21437 8812 21471
rect 8760 21428 8812 21437
rect 15476 21428 15528 21480
rect 15568 21471 15620 21480
rect 15568 21437 15577 21471
rect 15577 21437 15611 21471
rect 15611 21437 15620 21471
rect 15568 21428 15620 21437
rect 16948 21428 17000 21480
rect 19432 21496 19484 21548
rect 34520 21496 34572 21548
rect 34612 21539 34664 21548
rect 34612 21505 34621 21539
rect 34621 21505 34655 21539
rect 34655 21505 34664 21539
rect 34612 21496 34664 21505
rect 18696 21428 18748 21480
rect 19984 21428 20036 21480
rect 20444 21428 20496 21480
rect 22560 21471 22612 21480
rect 22560 21437 22569 21471
rect 22569 21437 22603 21471
rect 22603 21437 22612 21471
rect 22560 21428 22612 21437
rect 6276 21360 6328 21412
rect 8024 21360 8076 21412
rect 13728 21360 13780 21412
rect 15752 21360 15804 21412
rect 17040 21360 17092 21412
rect 19800 21360 19852 21412
rect 1768 21335 1820 21344
rect 1768 21301 1777 21335
rect 1777 21301 1811 21335
rect 1811 21301 1820 21335
rect 1768 21292 1820 21301
rect 5540 21292 5592 21344
rect 9772 21335 9824 21344
rect 9772 21301 9781 21335
rect 9781 21301 9815 21335
rect 9815 21301 9824 21335
rect 9772 21292 9824 21301
rect 12072 21335 12124 21344
rect 12072 21301 12081 21335
rect 12081 21301 12115 21335
rect 12115 21301 12124 21335
rect 12072 21292 12124 21301
rect 17132 21335 17184 21344
rect 17132 21301 17141 21335
rect 17141 21301 17175 21335
rect 17175 21301 17184 21335
rect 17132 21292 17184 21301
rect 17868 21335 17920 21344
rect 17868 21301 17877 21335
rect 17877 21301 17911 21335
rect 17911 21301 17920 21335
rect 17868 21292 17920 21301
rect 20904 21292 20956 21344
rect 34704 21335 34756 21344
rect 34704 21301 34713 21335
rect 34713 21301 34747 21335
rect 34747 21301 34756 21335
rect 34704 21292 34756 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6368 21088 6420 21140
rect 9036 21088 9088 21140
rect 12256 21088 12308 21140
rect 15200 21131 15252 21140
rect 15200 21097 15209 21131
rect 15209 21097 15243 21131
rect 15243 21097 15252 21131
rect 15200 21088 15252 21097
rect 16120 21131 16172 21140
rect 16120 21097 16129 21131
rect 16129 21097 16163 21131
rect 16163 21097 16172 21131
rect 16120 21088 16172 21097
rect 18696 21131 18748 21140
rect 18696 21097 18705 21131
rect 18705 21097 18739 21131
rect 18739 21097 18748 21131
rect 18696 21088 18748 21097
rect 19800 21131 19852 21140
rect 19800 21097 19809 21131
rect 19809 21097 19843 21131
rect 19843 21097 19852 21131
rect 19800 21088 19852 21097
rect 32036 21088 32088 21140
rect 12072 21020 12124 21072
rect 17868 21020 17920 21072
rect 9772 20995 9824 21004
rect 9772 20961 9781 20995
rect 9781 20961 9815 20995
rect 9815 20961 9824 20995
rect 9772 20952 9824 20961
rect 10968 20952 11020 21004
rect 19340 20952 19392 21004
rect 22560 20995 22612 21004
rect 22560 20961 22569 20995
rect 22569 20961 22603 20995
rect 22603 20961 22612 20995
rect 22560 20952 22612 20961
rect 23204 20995 23256 21004
rect 23204 20961 23213 20995
rect 23213 20961 23247 20995
rect 23247 20961 23256 20995
rect 23204 20952 23256 20961
rect 11244 20927 11296 20936
rect 10048 20816 10100 20868
rect 11244 20893 11253 20927
rect 11253 20893 11287 20927
rect 11287 20893 11296 20927
rect 11244 20884 11296 20893
rect 14464 20884 14516 20936
rect 13820 20816 13872 20868
rect 15568 20884 15620 20936
rect 15936 20927 15988 20936
rect 15936 20893 15945 20927
rect 15945 20893 15979 20927
rect 15979 20893 15988 20927
rect 15936 20884 15988 20893
rect 16856 20927 16908 20936
rect 16856 20893 16865 20927
rect 16865 20893 16899 20927
rect 16899 20893 16908 20927
rect 16856 20884 16908 20893
rect 18236 20884 18288 20936
rect 18420 20884 18472 20936
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 18052 20816 18104 20868
rect 19340 20816 19392 20868
rect 22376 20884 22428 20936
rect 28816 20927 28868 20936
rect 28816 20893 28825 20927
rect 28825 20893 28859 20927
rect 28859 20893 28868 20927
rect 28816 20884 28868 20893
rect 8944 20748 8996 20800
rect 15108 20748 15160 20800
rect 20628 20791 20680 20800
rect 20628 20757 20637 20791
rect 20637 20757 20671 20791
rect 20671 20757 20680 20791
rect 20628 20748 20680 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4896 20544 4948 20596
rect 5816 20544 5868 20596
rect 9588 20476 9640 20528
rect 15936 20544 15988 20596
rect 18052 20587 18104 20596
rect 18052 20553 18061 20587
rect 18061 20553 18095 20587
rect 18095 20553 18104 20587
rect 18052 20544 18104 20553
rect 18880 20544 18932 20596
rect 5540 20408 5592 20460
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 8944 20451 8996 20460
rect 8944 20417 8953 20451
rect 8953 20417 8987 20451
rect 8987 20417 8996 20451
rect 8944 20408 8996 20417
rect 10140 20451 10192 20460
rect 10140 20417 10149 20451
rect 10149 20417 10183 20451
rect 10183 20417 10192 20451
rect 10140 20408 10192 20417
rect 10324 20451 10376 20460
rect 10324 20417 10333 20451
rect 10333 20417 10367 20451
rect 10367 20417 10376 20451
rect 10324 20408 10376 20417
rect 11612 20408 11664 20460
rect 16948 20476 17000 20528
rect 13912 20451 13964 20460
rect 13912 20417 13921 20451
rect 13921 20417 13955 20451
rect 13955 20417 13964 20451
rect 13912 20408 13964 20417
rect 14004 20408 14056 20460
rect 14372 20451 14424 20460
rect 14372 20417 14381 20451
rect 14381 20417 14415 20451
rect 14415 20417 14424 20451
rect 14372 20408 14424 20417
rect 15016 20451 15068 20460
rect 15016 20417 15025 20451
rect 15025 20417 15059 20451
rect 15059 20417 15068 20451
rect 15016 20408 15068 20417
rect 15108 20408 15160 20460
rect 17132 20408 17184 20460
rect 21824 20544 21876 20596
rect 22376 20544 22428 20596
rect 20812 20519 20864 20528
rect 20812 20485 20821 20519
rect 20821 20485 20855 20519
rect 20855 20485 20864 20519
rect 20812 20476 20864 20485
rect 9864 20340 9916 20392
rect 9036 20272 9088 20324
rect 17040 20340 17092 20392
rect 14924 20272 14976 20324
rect 17224 20272 17276 20324
rect 10600 20247 10652 20256
rect 10600 20213 10609 20247
rect 10609 20213 10643 20247
rect 10643 20213 10652 20247
rect 10600 20204 10652 20213
rect 13728 20247 13780 20256
rect 13728 20213 13737 20247
rect 13737 20213 13771 20247
rect 13771 20213 13780 20247
rect 13728 20204 13780 20213
rect 15200 20204 15252 20256
rect 16580 20204 16632 20256
rect 17500 20272 17552 20324
rect 19984 20340 20036 20392
rect 21824 20340 21876 20392
rect 22008 20340 22060 20392
rect 24584 20340 24636 20392
rect 25228 20272 25280 20324
rect 20260 20204 20312 20256
rect 22836 20247 22888 20256
rect 22836 20213 22845 20247
rect 22845 20213 22879 20247
rect 22879 20213 22888 20247
rect 22836 20204 22888 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7012 20000 7064 20052
rect 10508 20000 10560 20052
rect 12992 20000 13044 20052
rect 14464 20043 14516 20052
rect 14464 20009 14473 20043
rect 14473 20009 14507 20043
rect 14507 20009 14516 20043
rect 14464 20000 14516 20009
rect 16120 20043 16172 20052
rect 16120 20009 16129 20043
rect 16129 20009 16163 20043
rect 16163 20009 16172 20043
rect 16120 20000 16172 20009
rect 1768 19839 1820 19848
rect 1768 19805 1777 19839
rect 1777 19805 1811 19839
rect 1811 19805 1820 19839
rect 1768 19796 1820 19805
rect 7840 19796 7892 19848
rect 9220 19796 9272 19848
rect 9864 19839 9916 19848
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 13268 19932 13320 19984
rect 22836 20000 22888 20052
rect 24584 20043 24636 20052
rect 24584 20009 24593 20043
rect 24593 20009 24627 20043
rect 24627 20009 24636 20043
rect 24584 20000 24636 20009
rect 13728 19864 13780 19916
rect 11520 19796 11572 19848
rect 11796 19796 11848 19848
rect 13820 19796 13872 19848
rect 15016 19796 15068 19848
rect 15476 19796 15528 19848
rect 19340 19796 19392 19848
rect 5540 19660 5592 19712
rect 12808 19728 12860 19780
rect 14280 19728 14332 19780
rect 7932 19660 7984 19712
rect 10600 19660 10652 19712
rect 13452 19660 13504 19712
rect 15384 19728 15436 19780
rect 16672 19728 16724 19780
rect 17224 19771 17276 19780
rect 17224 19737 17233 19771
rect 17233 19737 17267 19771
rect 17267 19737 17276 19771
rect 17224 19728 17276 19737
rect 18144 19728 18196 19780
rect 16764 19660 16816 19712
rect 16856 19660 16908 19712
rect 20076 19660 20128 19712
rect 23204 19907 23256 19916
rect 23204 19873 23213 19907
rect 23213 19873 23247 19907
rect 23247 19873 23256 19907
rect 23204 19864 23256 19873
rect 21548 19839 21600 19848
rect 21548 19805 21557 19839
rect 21557 19805 21591 19839
rect 21591 19805 21600 19839
rect 21548 19796 21600 19805
rect 23848 19839 23900 19848
rect 23848 19805 23857 19839
rect 23857 19805 23891 19839
rect 23891 19805 23900 19839
rect 23848 19796 23900 19805
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 25412 19839 25464 19848
rect 25412 19805 25421 19839
rect 25421 19805 25455 19839
rect 25455 19805 25464 19839
rect 25412 19796 25464 19805
rect 38292 19839 38344 19848
rect 38292 19805 38301 19839
rect 38301 19805 38335 19839
rect 38335 19805 38344 19839
rect 38292 19796 38344 19805
rect 22744 19771 22796 19780
rect 22744 19737 22753 19771
rect 22753 19737 22787 19771
rect 22787 19737 22796 19771
rect 22744 19728 22796 19737
rect 22836 19771 22888 19780
rect 22836 19737 22845 19771
rect 22845 19737 22879 19771
rect 22879 19737 22888 19771
rect 22836 19728 22888 19737
rect 24860 19660 24912 19712
rect 25228 19703 25280 19712
rect 25228 19669 25237 19703
rect 25237 19669 25271 19703
rect 25271 19669 25280 19703
rect 25228 19660 25280 19669
rect 37004 19660 37056 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 5632 19320 5684 19372
rect 7748 19320 7800 19372
rect 9220 19363 9272 19372
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 10600 19320 10652 19372
rect 10508 19295 10560 19304
rect 10508 19261 10517 19295
rect 10517 19261 10551 19295
rect 10551 19261 10560 19295
rect 10508 19252 10560 19261
rect 12992 19388 13044 19440
rect 13912 19456 13964 19508
rect 14924 19456 14976 19508
rect 16672 19456 16724 19508
rect 16856 19499 16908 19508
rect 16856 19465 16865 19499
rect 16865 19465 16899 19499
rect 16899 19465 16908 19499
rect 16856 19456 16908 19465
rect 17500 19499 17552 19508
rect 17500 19465 17509 19499
rect 17509 19465 17543 19499
rect 17543 19465 17552 19499
rect 17500 19456 17552 19465
rect 18144 19499 18196 19508
rect 18144 19465 18153 19499
rect 18153 19465 18187 19499
rect 18187 19465 18196 19499
rect 18144 19456 18196 19465
rect 13084 19320 13136 19372
rect 15292 19388 15344 19440
rect 20904 19456 20956 19508
rect 22836 19456 22888 19508
rect 25412 19456 25464 19508
rect 20076 19431 20128 19440
rect 14924 19363 14976 19372
rect 14924 19329 14933 19363
rect 14933 19329 14967 19363
rect 14967 19329 14976 19363
rect 14924 19320 14976 19329
rect 11060 19252 11112 19304
rect 13820 19252 13872 19304
rect 13912 19295 13964 19304
rect 13912 19261 13921 19295
rect 13921 19261 13955 19295
rect 13955 19261 13964 19295
rect 20076 19397 20085 19431
rect 20085 19397 20119 19431
rect 20119 19397 20128 19431
rect 20076 19388 20128 19397
rect 21364 19388 21416 19440
rect 22008 19388 22060 19440
rect 16764 19320 16816 19372
rect 17132 19320 17184 19372
rect 18788 19363 18840 19372
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 19432 19363 19484 19372
rect 19432 19329 19441 19363
rect 19441 19329 19475 19363
rect 19475 19329 19484 19363
rect 19432 19320 19484 19329
rect 21732 19320 21784 19372
rect 22928 19388 22980 19440
rect 25228 19388 25280 19440
rect 24676 19363 24728 19372
rect 24676 19329 24685 19363
rect 24685 19329 24719 19363
rect 24719 19329 24728 19363
rect 24676 19320 24728 19329
rect 13912 19252 13964 19261
rect 18972 19295 19024 19304
rect 11244 19184 11296 19236
rect 11336 19184 11388 19236
rect 7472 19116 7524 19168
rect 12256 19116 12308 19168
rect 12808 19184 12860 19236
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 20076 19252 20128 19304
rect 23664 19252 23716 19304
rect 29736 19252 29788 19304
rect 20444 19184 20496 19236
rect 28724 19184 28776 19236
rect 13268 19116 13320 19168
rect 13360 19116 13412 19168
rect 14372 19116 14424 19168
rect 14924 19116 14976 19168
rect 21180 19159 21232 19168
rect 21180 19125 21189 19159
rect 21189 19125 21223 19159
rect 21223 19125 21232 19159
rect 21180 19116 21232 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 10600 18912 10652 18964
rect 9772 18844 9824 18896
rect 6644 18640 6696 18692
rect 9036 18640 9088 18692
rect 10784 18708 10836 18760
rect 9680 18640 9732 18692
rect 7104 18572 7156 18624
rect 11704 18572 11756 18624
rect 12256 18912 12308 18964
rect 11980 18844 12032 18896
rect 13360 18844 13412 18896
rect 13452 18844 13504 18896
rect 12532 18572 12584 18624
rect 14004 18776 14056 18828
rect 14280 18819 14332 18828
rect 14280 18785 14289 18819
rect 14289 18785 14323 18819
rect 14323 18785 14332 18819
rect 14280 18776 14332 18785
rect 15660 18751 15712 18760
rect 15660 18717 15669 18751
rect 15669 18717 15703 18751
rect 15703 18717 15712 18751
rect 15660 18708 15712 18717
rect 17132 18912 17184 18964
rect 17316 18912 17368 18964
rect 24768 18912 24820 18964
rect 20260 18844 20312 18896
rect 20444 18887 20496 18896
rect 20444 18853 20453 18887
rect 20453 18853 20487 18887
rect 20487 18853 20496 18887
rect 20444 18844 20496 18853
rect 20168 18776 20220 18828
rect 30564 18844 30616 18896
rect 21180 18819 21232 18828
rect 21180 18785 21189 18819
rect 21189 18785 21223 18819
rect 21223 18785 21232 18819
rect 21180 18776 21232 18785
rect 23664 18819 23716 18828
rect 23664 18785 23673 18819
rect 23673 18785 23707 18819
rect 23707 18785 23716 18819
rect 23664 18776 23716 18785
rect 17132 18708 17184 18760
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 13820 18572 13872 18624
rect 17868 18572 17920 18624
rect 20628 18640 20680 18692
rect 21180 18572 21232 18624
rect 37004 18708 37056 18760
rect 38292 18751 38344 18760
rect 38292 18717 38301 18751
rect 38301 18717 38335 18751
rect 38335 18717 38344 18751
rect 38292 18708 38344 18717
rect 23020 18683 23072 18692
rect 23020 18649 23029 18683
rect 23029 18649 23063 18683
rect 23063 18649 23072 18683
rect 23020 18640 23072 18649
rect 23112 18683 23164 18692
rect 23112 18649 23121 18683
rect 23121 18649 23155 18683
rect 23155 18649 23164 18683
rect 23112 18640 23164 18649
rect 23848 18572 23900 18624
rect 33140 18615 33192 18624
rect 33140 18581 33149 18615
rect 33149 18581 33183 18615
rect 33183 18581 33192 18615
rect 33140 18572 33192 18581
rect 34520 18572 34572 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 7656 18368 7708 18420
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 9680 18411 9732 18420
rect 9680 18377 9689 18411
rect 9689 18377 9723 18411
rect 9723 18377 9732 18411
rect 9680 18368 9732 18377
rect 7104 18343 7156 18352
rect 7104 18309 7113 18343
rect 7113 18309 7147 18343
rect 7147 18309 7156 18343
rect 7104 18300 7156 18309
rect 7196 18343 7248 18352
rect 7196 18309 7205 18343
rect 7205 18309 7239 18343
rect 7239 18309 7248 18343
rect 7196 18300 7248 18309
rect 8668 18300 8720 18352
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 8576 18275 8628 18284
rect 8576 18241 8585 18275
rect 8585 18241 8619 18275
rect 8619 18241 8628 18275
rect 8576 18232 8628 18241
rect 9220 18275 9272 18284
rect 9220 18241 9229 18275
rect 9229 18241 9263 18275
rect 9263 18241 9272 18275
rect 9220 18232 9272 18241
rect 13360 18368 13412 18420
rect 7748 18164 7800 18216
rect 11336 18300 11388 18352
rect 18972 18368 19024 18420
rect 21180 18411 21232 18420
rect 21180 18377 21189 18411
rect 21189 18377 21223 18411
rect 21223 18377 21232 18411
rect 21180 18368 21232 18377
rect 23112 18368 23164 18420
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 3056 18028 3108 18080
rect 3976 18028 4028 18080
rect 8944 18028 8996 18080
rect 11796 18275 11848 18284
rect 11796 18241 11805 18275
rect 11805 18241 11839 18275
rect 11839 18241 11848 18275
rect 11796 18232 11848 18241
rect 12992 18232 13044 18284
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 11244 18164 11296 18216
rect 12256 18096 12308 18148
rect 12348 18096 12400 18148
rect 12532 18096 12584 18148
rect 13360 18164 13412 18216
rect 17592 18232 17644 18284
rect 13084 18028 13136 18080
rect 14096 18028 14148 18080
rect 14832 18071 14884 18080
rect 14832 18037 14841 18071
rect 14841 18037 14875 18071
rect 14875 18037 14884 18071
rect 14832 18028 14884 18037
rect 15292 18164 15344 18216
rect 16948 18207 17000 18216
rect 16948 18173 16957 18207
rect 16957 18173 16991 18207
rect 16991 18173 17000 18207
rect 16948 18164 17000 18173
rect 21548 18232 21600 18284
rect 19064 18207 19116 18216
rect 19064 18173 19073 18207
rect 19073 18173 19107 18207
rect 19107 18173 19116 18207
rect 19064 18164 19116 18173
rect 20720 18207 20772 18216
rect 18144 18028 18196 18080
rect 20352 18028 20404 18080
rect 20720 18173 20729 18207
rect 20729 18173 20763 18207
rect 20763 18173 20772 18207
rect 20720 18164 20772 18173
rect 22652 18207 22704 18216
rect 22652 18173 22661 18207
rect 22661 18173 22695 18207
rect 22695 18173 22704 18207
rect 22652 18164 22704 18173
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 24400 18275 24452 18284
rect 23572 18232 23624 18241
rect 24400 18241 24409 18275
rect 24409 18241 24443 18275
rect 24443 18241 24452 18275
rect 24400 18232 24452 18241
rect 33324 18164 33376 18216
rect 29644 18096 29696 18148
rect 21640 18028 21692 18080
rect 22744 18028 22796 18080
rect 24216 18071 24268 18080
rect 24216 18037 24225 18071
rect 24225 18037 24259 18071
rect 24259 18037 24268 18071
rect 24216 18028 24268 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 7196 17824 7248 17876
rect 9220 17824 9272 17876
rect 13820 17824 13872 17876
rect 16948 17867 17000 17876
rect 16948 17833 16957 17867
rect 16957 17833 16991 17867
rect 16991 17833 17000 17867
rect 16948 17824 17000 17833
rect 10140 17756 10192 17808
rect 14464 17756 14516 17808
rect 16120 17756 16172 17808
rect 16304 17756 16356 17808
rect 2320 17620 2372 17672
rect 2780 17620 2832 17672
rect 3240 17663 3292 17672
rect 3240 17629 3249 17663
rect 3249 17629 3283 17663
rect 3283 17629 3292 17663
rect 3240 17620 3292 17629
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 7012 17620 7064 17672
rect 7840 17688 7892 17740
rect 8852 17688 8904 17740
rect 9772 17688 9824 17740
rect 10876 17731 10928 17740
rect 10876 17697 10885 17731
rect 10885 17697 10919 17731
rect 10919 17697 10928 17731
rect 10876 17688 10928 17697
rect 10968 17620 11020 17672
rect 12992 17688 13044 17740
rect 13544 17688 13596 17740
rect 15384 17731 15436 17740
rect 15384 17697 15393 17731
rect 15393 17697 15427 17731
rect 15427 17697 15436 17731
rect 15384 17688 15436 17697
rect 16028 17731 16080 17740
rect 16028 17697 16037 17731
rect 16037 17697 16071 17731
rect 16071 17697 16080 17731
rect 16028 17688 16080 17697
rect 12348 17620 12400 17672
rect 12716 17620 12768 17672
rect 14832 17663 14884 17672
rect 14832 17629 14841 17663
rect 14841 17629 14875 17663
rect 14875 17629 14884 17663
rect 14832 17620 14884 17629
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 18236 17824 18288 17876
rect 19064 17824 19116 17876
rect 20720 17824 20772 17876
rect 1860 17484 1912 17536
rect 2504 17527 2556 17536
rect 2504 17493 2513 17527
rect 2513 17493 2547 17527
rect 2547 17493 2556 17527
rect 2504 17484 2556 17493
rect 2596 17484 2648 17536
rect 4712 17484 4764 17536
rect 9772 17552 9824 17604
rect 10232 17595 10284 17604
rect 10232 17561 10241 17595
rect 10241 17561 10275 17595
rect 10275 17561 10284 17595
rect 10232 17552 10284 17561
rect 8300 17484 8352 17536
rect 15476 17595 15528 17604
rect 15476 17561 15485 17595
rect 15485 17561 15519 17595
rect 15519 17561 15528 17595
rect 15476 17552 15528 17561
rect 17868 17620 17920 17672
rect 16856 17552 16908 17604
rect 21180 17688 21232 17740
rect 21640 17824 21692 17876
rect 22652 17824 22704 17876
rect 22744 17799 22796 17808
rect 22744 17765 22753 17799
rect 22753 17765 22787 17799
rect 22787 17765 22796 17799
rect 22744 17756 22796 17765
rect 22284 17688 22336 17740
rect 24216 17688 24268 17740
rect 21732 17663 21784 17672
rect 21732 17629 21741 17663
rect 21741 17629 21775 17663
rect 21775 17629 21784 17663
rect 21732 17620 21784 17629
rect 23296 17663 23348 17672
rect 23296 17629 23305 17663
rect 23305 17629 23339 17663
rect 23339 17629 23348 17663
rect 23296 17620 23348 17629
rect 38108 17688 38160 17740
rect 34520 17620 34572 17672
rect 29092 17552 29144 17604
rect 18236 17527 18288 17536
rect 18236 17493 18245 17527
rect 18245 17493 18279 17527
rect 18279 17493 18288 17527
rect 18236 17484 18288 17493
rect 20444 17484 20496 17536
rect 31576 17527 31628 17536
rect 31576 17493 31585 17527
rect 31585 17493 31619 17527
rect 31619 17493 31628 17527
rect 31576 17484 31628 17493
rect 33232 17527 33284 17536
rect 33232 17493 33241 17527
rect 33241 17493 33275 17527
rect 33275 17493 33284 17527
rect 33232 17484 33284 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 8576 17323 8628 17332
rect 8576 17289 8585 17323
rect 8585 17289 8619 17323
rect 8619 17289 8628 17323
rect 8576 17280 8628 17289
rect 10232 17280 10284 17332
rect 11060 17323 11112 17332
rect 11060 17289 11069 17323
rect 11069 17289 11103 17323
rect 11103 17289 11112 17323
rect 11060 17280 11112 17289
rect 4712 17255 4764 17264
rect 4712 17221 4721 17255
rect 4721 17221 4755 17255
rect 4755 17221 4764 17255
rect 4712 17212 4764 17221
rect 11796 17212 11848 17264
rect 16488 17280 16540 17332
rect 16948 17280 17000 17332
rect 19432 17280 19484 17332
rect 19984 17323 20036 17332
rect 19984 17289 19993 17323
rect 19993 17289 20027 17323
rect 20027 17289 20036 17323
rect 19984 17280 20036 17289
rect 20812 17280 20864 17332
rect 23020 17280 23072 17332
rect 24400 17280 24452 17332
rect 2412 17144 2464 17196
rect 2780 17144 2832 17196
rect 3148 17144 3200 17196
rect 7288 17144 7340 17196
rect 8852 17144 8904 17196
rect 8944 17144 8996 17196
rect 10968 17187 11020 17196
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 14372 17212 14424 17264
rect 15292 17212 15344 17264
rect 12440 17144 12492 17153
rect 13268 17144 13320 17196
rect 16764 17144 16816 17196
rect 17224 17144 17276 17196
rect 20076 17212 20128 17264
rect 20260 17212 20312 17264
rect 18972 17144 19024 17196
rect 31576 17212 31628 17264
rect 23112 17144 23164 17196
rect 23296 17187 23348 17196
rect 23296 17153 23305 17187
rect 23305 17153 23339 17187
rect 23339 17153 23348 17187
rect 23296 17144 23348 17153
rect 23848 17144 23900 17196
rect 24584 17187 24636 17196
rect 24584 17153 24593 17187
rect 24593 17153 24627 17187
rect 24627 17153 24636 17187
rect 24584 17144 24636 17153
rect 35900 17144 35952 17196
rect 4620 17119 4672 17128
rect 4620 17085 4629 17119
rect 4629 17085 4663 17119
rect 4663 17085 4672 17119
rect 4620 17076 4672 17085
rect 4804 17076 4856 17128
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 9312 17076 9364 17128
rect 14280 17076 14332 17128
rect 3332 17051 3384 17060
rect 3332 17017 3341 17051
rect 3341 17017 3375 17051
rect 3375 17017 3384 17051
rect 3332 17008 3384 17017
rect 11428 17008 11480 17060
rect 11612 17008 11664 17060
rect 14464 17076 14516 17128
rect 2136 16940 2188 16992
rect 2688 16983 2740 16992
rect 2688 16949 2697 16983
rect 2697 16949 2731 16983
rect 2731 16949 2740 16983
rect 2688 16940 2740 16949
rect 6460 16940 6512 16992
rect 6920 16940 6972 16992
rect 9680 16983 9732 16992
rect 9680 16949 9689 16983
rect 9689 16949 9723 16983
rect 9723 16949 9732 16983
rect 9680 16940 9732 16949
rect 15476 17008 15528 17060
rect 19340 17119 19392 17128
rect 19340 17085 19349 17119
rect 19349 17085 19383 17119
rect 19383 17085 19392 17119
rect 19340 17076 19392 17085
rect 19432 17076 19484 17128
rect 22008 17119 22060 17128
rect 22008 17085 22017 17119
rect 22017 17085 22051 17119
rect 22051 17085 22060 17119
rect 22008 17076 22060 17085
rect 22836 17076 22888 17128
rect 38200 17051 38252 17060
rect 38200 17017 38209 17051
rect 38209 17017 38243 17051
rect 38243 17017 38252 17051
rect 38200 17008 38252 17017
rect 16856 16940 16908 16992
rect 17316 16940 17368 16992
rect 22008 16940 22060 16992
rect 23480 16940 23532 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 11612 16779 11664 16788
rect 11612 16745 11621 16779
rect 11621 16745 11655 16779
rect 11655 16745 11664 16779
rect 11612 16736 11664 16745
rect 12440 16736 12492 16788
rect 16764 16779 16816 16788
rect 16764 16745 16773 16779
rect 16773 16745 16807 16779
rect 16807 16745 16816 16779
rect 16764 16736 16816 16745
rect 22836 16779 22888 16788
rect 22836 16745 22845 16779
rect 22845 16745 22879 16779
rect 22879 16745 22888 16779
rect 22836 16736 22888 16745
rect 8484 16711 8536 16720
rect 8484 16677 8493 16711
rect 8493 16677 8527 16711
rect 8527 16677 8536 16711
rect 8484 16668 8536 16677
rect 13360 16668 13412 16720
rect 16028 16711 16080 16720
rect 16028 16677 16037 16711
rect 16037 16677 16071 16711
rect 16071 16677 16080 16711
rect 16028 16668 16080 16677
rect 20444 16668 20496 16720
rect 1676 16532 1728 16584
rect 2412 16532 2464 16584
rect 2964 16575 3016 16584
rect 2964 16541 2973 16575
rect 2973 16541 3007 16575
rect 3007 16541 3016 16575
rect 2964 16532 3016 16541
rect 4620 16600 4672 16652
rect 5540 16600 5592 16652
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 6460 16643 6512 16652
rect 6460 16609 6469 16643
rect 6469 16609 6503 16643
rect 6503 16609 6512 16643
rect 6460 16600 6512 16609
rect 7932 16643 7984 16652
rect 7932 16609 7941 16643
rect 7941 16609 7975 16643
rect 7975 16609 7984 16643
rect 7932 16600 7984 16609
rect 8300 16600 8352 16652
rect 9036 16532 9088 16584
rect 12716 16600 12768 16652
rect 17408 16600 17460 16652
rect 18512 16600 18564 16652
rect 20904 16668 20956 16720
rect 21272 16600 21324 16652
rect 10416 16532 10468 16584
rect 2780 16464 2832 16516
rect 1768 16439 1820 16448
rect 1768 16405 1777 16439
rect 1777 16405 1811 16439
rect 1811 16405 1820 16439
rect 1768 16396 1820 16405
rect 2872 16396 2924 16448
rect 3332 16396 3384 16448
rect 5724 16439 5776 16448
rect 5724 16405 5733 16439
rect 5733 16405 5767 16439
rect 5767 16405 5776 16439
rect 5724 16396 5776 16405
rect 6920 16439 6972 16448
rect 6920 16405 6929 16439
rect 6929 16405 6963 16439
rect 6963 16405 6972 16439
rect 6920 16396 6972 16405
rect 7196 16396 7248 16448
rect 9680 16396 9732 16448
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 13636 16532 13688 16584
rect 12992 16464 13044 16516
rect 16856 16532 16908 16584
rect 17592 16575 17644 16584
rect 11796 16396 11848 16448
rect 15568 16507 15620 16516
rect 15568 16473 15577 16507
rect 15577 16473 15611 16507
rect 15611 16473 15620 16507
rect 15568 16464 15620 16473
rect 15752 16464 15804 16516
rect 16764 16464 16816 16516
rect 17592 16541 17601 16575
rect 17601 16541 17635 16575
rect 17635 16541 17644 16575
rect 17592 16532 17644 16541
rect 19340 16532 19392 16584
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 33232 16600 33284 16652
rect 23480 16532 23532 16584
rect 23664 16575 23716 16584
rect 23664 16541 23673 16575
rect 23673 16541 23707 16575
rect 23707 16541 23716 16575
rect 23664 16532 23716 16541
rect 19432 16396 19484 16448
rect 20076 16396 20128 16448
rect 20904 16396 20956 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 5172 16192 5224 16244
rect 5724 16192 5776 16244
rect 2964 16124 3016 16176
rect 2044 16056 2096 16108
rect 2412 16056 2464 16108
rect 5264 16124 5316 16176
rect 7012 16124 7064 16176
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 5540 16099 5592 16108
rect 5540 16065 5549 16099
rect 5549 16065 5583 16099
rect 5583 16065 5592 16099
rect 5540 16056 5592 16065
rect 7288 16056 7340 16108
rect 7840 16056 7892 16108
rect 3976 15988 4028 16040
rect 1492 15852 1544 15904
rect 2688 15852 2740 15904
rect 3516 15852 3568 15904
rect 5632 15852 5684 15904
rect 8024 15852 8076 15904
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 9772 16192 9824 16244
rect 10784 16192 10836 16244
rect 9312 16124 9364 16176
rect 10876 16124 10928 16176
rect 12624 16192 12676 16244
rect 21180 16235 21232 16244
rect 9864 16099 9916 16108
rect 9864 16065 9873 16099
rect 9873 16065 9907 16099
rect 9907 16065 9916 16099
rect 9864 16056 9916 16065
rect 12348 16099 12400 16108
rect 12348 16065 12357 16099
rect 12357 16065 12391 16099
rect 12391 16065 12400 16099
rect 12348 16056 12400 16065
rect 20628 16124 20680 16176
rect 21180 16201 21189 16235
rect 21189 16201 21223 16235
rect 21223 16201 21232 16235
rect 21180 16192 21232 16201
rect 23020 16192 23072 16244
rect 23112 16192 23164 16244
rect 21732 16124 21784 16176
rect 13360 16056 13412 16108
rect 15660 16099 15712 16108
rect 11612 15988 11664 16040
rect 13452 16031 13504 16040
rect 13452 15997 13461 16031
rect 13461 15997 13495 16031
rect 13495 15997 13504 16031
rect 13452 15988 13504 15997
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 17868 16056 17920 16108
rect 16948 15988 17000 16040
rect 12440 15920 12492 15972
rect 13636 15920 13688 15972
rect 16672 15920 16724 15972
rect 20904 16056 20956 16108
rect 21548 16056 21600 16108
rect 23848 16099 23900 16108
rect 23848 16065 23857 16099
rect 23857 16065 23891 16099
rect 23891 16065 23900 16099
rect 23848 16056 23900 16065
rect 38108 16056 38160 16108
rect 9956 15852 10008 15904
rect 10692 15852 10744 15904
rect 12624 15852 12676 15904
rect 13176 15852 13228 15904
rect 14556 15852 14608 15904
rect 17500 15920 17552 15972
rect 19616 15920 19668 15972
rect 20812 15988 20864 16040
rect 17224 15895 17276 15904
rect 17224 15861 17233 15895
rect 17233 15861 17267 15895
rect 17267 15861 17276 15895
rect 17224 15852 17276 15861
rect 20444 15895 20496 15904
rect 20444 15861 20453 15895
rect 20453 15861 20487 15895
rect 20487 15861 20496 15895
rect 20444 15852 20496 15861
rect 23112 15852 23164 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 7196 15691 7248 15700
rect 7196 15657 7205 15691
rect 7205 15657 7239 15691
rect 7239 15657 7248 15691
rect 7196 15648 7248 15657
rect 9312 15691 9364 15700
rect 9312 15657 9321 15691
rect 9321 15657 9355 15691
rect 9355 15657 9364 15691
rect 9312 15648 9364 15657
rect 10692 15648 10744 15700
rect 12532 15648 12584 15700
rect 13176 15648 13228 15700
rect 15568 15648 15620 15700
rect 17224 15648 17276 15700
rect 7104 15580 7156 15632
rect 8484 15623 8536 15632
rect 8484 15589 8493 15623
rect 8493 15589 8527 15623
rect 8527 15589 8536 15623
rect 8484 15580 8536 15589
rect 13452 15580 13504 15632
rect 21456 15623 21508 15632
rect 9680 15512 9732 15564
rect 12624 15512 12676 15564
rect 15016 15512 15068 15564
rect 16212 15512 16264 15564
rect 21456 15589 21465 15623
rect 21465 15589 21499 15623
rect 21499 15589 21508 15623
rect 21456 15580 21508 15589
rect 23664 15648 23716 15700
rect 35900 15648 35952 15700
rect 38108 15691 38160 15700
rect 38108 15657 38117 15691
rect 38117 15657 38151 15691
rect 38151 15657 38160 15691
rect 38108 15648 38160 15657
rect 32404 15580 32456 15632
rect 19616 15512 19668 15564
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 2596 15444 2648 15496
rect 3608 15444 3660 15496
rect 5172 15444 5224 15496
rect 5356 15487 5408 15496
rect 5356 15453 5365 15487
rect 5365 15453 5399 15487
rect 5399 15453 5408 15487
rect 5356 15444 5408 15453
rect 7012 15444 7064 15496
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 9772 15444 9824 15496
rect 8392 15376 8444 15428
rect 9680 15376 9732 15428
rect 10416 15444 10468 15496
rect 10600 15444 10652 15496
rect 12072 15444 12124 15496
rect 12716 15444 12768 15496
rect 13176 15444 13228 15496
rect 16304 15444 16356 15496
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 16488 15444 16540 15453
rect 16672 15487 16724 15496
rect 16672 15453 16681 15487
rect 16681 15453 16715 15487
rect 16715 15453 16724 15487
rect 16672 15444 16724 15453
rect 16948 15444 17000 15496
rect 14740 15376 14792 15428
rect 22560 15512 22612 15564
rect 22928 15444 22980 15496
rect 23112 15512 23164 15564
rect 33140 15512 33192 15564
rect 31944 15444 31996 15496
rect 38292 15487 38344 15496
rect 38292 15453 38301 15487
rect 38301 15453 38335 15487
rect 38335 15453 38344 15487
rect 38292 15444 38344 15453
rect 2688 15308 2740 15360
rect 3056 15351 3108 15360
rect 3056 15317 3065 15351
rect 3065 15317 3099 15351
rect 3099 15317 3108 15351
rect 3056 15308 3108 15317
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 4620 15308 4672 15317
rect 4804 15308 4856 15360
rect 6276 15351 6328 15360
rect 6276 15317 6285 15351
rect 6285 15317 6319 15351
rect 6319 15317 6328 15351
rect 6276 15308 6328 15317
rect 7840 15308 7892 15360
rect 11336 15308 11388 15360
rect 13176 15308 13228 15360
rect 13636 15308 13688 15360
rect 17040 15308 17092 15360
rect 20260 15308 20312 15360
rect 24584 15376 24636 15428
rect 20628 15308 20680 15360
rect 23480 15351 23532 15360
rect 23480 15317 23489 15351
rect 23489 15317 23523 15351
rect 23523 15317 23532 15351
rect 23480 15308 23532 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 5356 15104 5408 15156
rect 7380 15104 7432 15156
rect 7564 15104 7616 15156
rect 8392 15104 8444 15156
rect 1584 14968 1636 15020
rect 2136 14968 2188 15020
rect 3148 14968 3200 15020
rect 6276 15036 6328 15088
rect 5172 14968 5224 15020
rect 5540 14968 5592 15020
rect 5816 14968 5868 15020
rect 8024 15011 8076 15020
rect 6276 14900 6328 14952
rect 8024 14977 8033 15011
rect 8033 14977 8067 15011
rect 8067 14977 8076 15011
rect 8024 14968 8076 14977
rect 12532 15104 12584 15156
rect 14556 15104 14608 15156
rect 16212 15147 16264 15156
rect 16212 15113 16221 15147
rect 16221 15113 16255 15147
rect 16255 15113 16264 15147
rect 16212 15104 16264 15113
rect 16396 15104 16448 15156
rect 11704 15036 11756 15088
rect 19340 15104 19392 15156
rect 20444 15104 20496 15156
rect 21272 15147 21324 15156
rect 21272 15113 21281 15147
rect 21281 15113 21315 15147
rect 21315 15113 21324 15147
rect 21272 15104 21324 15113
rect 22928 15104 22980 15156
rect 17500 15036 17552 15088
rect 20720 15036 20772 15088
rect 9404 14943 9456 14952
rect 9404 14909 9413 14943
rect 9413 14909 9447 14943
rect 9447 14909 9456 14943
rect 9404 14900 9456 14909
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 11888 14900 11940 14952
rect 12164 14943 12216 14952
rect 12164 14909 12173 14943
rect 12173 14909 12207 14943
rect 12207 14909 12216 14943
rect 12164 14900 12216 14909
rect 13820 14968 13872 15020
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 16304 14968 16356 15020
rect 17868 14968 17920 15020
rect 10968 14832 11020 14884
rect 11060 14832 11112 14884
rect 17224 14943 17276 14952
rect 17224 14909 17234 14943
rect 17234 14909 17268 14943
rect 17268 14909 17276 14943
rect 18420 14943 18472 14952
rect 17224 14900 17276 14909
rect 18420 14909 18429 14943
rect 18429 14909 18463 14943
rect 18463 14909 18472 14943
rect 18420 14900 18472 14909
rect 20260 14968 20312 15020
rect 22560 15036 22612 15088
rect 19984 14900 20036 14952
rect 22652 14900 22704 14952
rect 23480 14968 23532 15020
rect 33416 14900 33468 14952
rect 16580 14832 16632 14884
rect 17684 14832 17736 14884
rect 19432 14832 19484 14884
rect 20168 14832 20220 14884
rect 21456 14832 21508 14884
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 3424 14764 3476 14816
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 4712 14764 4764 14816
rect 5356 14764 5408 14816
rect 6736 14764 6788 14816
rect 8576 14764 8628 14816
rect 11152 14764 11204 14816
rect 12164 14764 12216 14816
rect 17868 14764 17920 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2320 14560 2372 14612
rect 4528 14560 4580 14612
rect 2688 14492 2740 14544
rect 3056 14424 3108 14476
rect 3424 14399 3476 14408
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 8484 14492 8536 14544
rect 10692 14560 10744 14612
rect 11060 14603 11112 14612
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 11704 14603 11756 14612
rect 11704 14569 11713 14603
rect 11713 14569 11747 14603
rect 11747 14569 11756 14603
rect 11704 14560 11756 14569
rect 12348 14560 12400 14612
rect 14832 14560 14884 14612
rect 15016 14603 15068 14612
rect 15016 14569 15025 14603
rect 15025 14569 15059 14603
rect 15059 14569 15068 14603
rect 15016 14560 15068 14569
rect 15108 14560 15160 14612
rect 16856 14560 16908 14612
rect 17592 14560 17644 14612
rect 20076 14560 20128 14612
rect 20812 14603 20864 14612
rect 20812 14569 20821 14603
rect 20821 14569 20855 14603
rect 20855 14569 20864 14603
rect 20812 14560 20864 14569
rect 22652 14603 22704 14612
rect 22652 14569 22661 14603
rect 22661 14569 22695 14603
rect 22695 14569 22704 14603
rect 22652 14560 22704 14569
rect 31944 14560 31996 14612
rect 4620 14424 4672 14476
rect 4896 14424 4948 14476
rect 8576 14467 8628 14476
rect 8576 14433 8585 14467
rect 8585 14433 8619 14467
rect 8619 14433 8628 14467
rect 8576 14424 8628 14433
rect 7932 14399 7984 14408
rect 4896 14288 4948 14340
rect 5356 14331 5408 14340
rect 5356 14297 5365 14331
rect 5365 14297 5399 14331
rect 5399 14297 5408 14331
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 5356 14288 5408 14297
rect 9588 14288 9640 14340
rect 10692 14356 10744 14408
rect 11520 14356 11572 14408
rect 12716 14424 12768 14476
rect 16488 14424 16540 14476
rect 16580 14424 16632 14476
rect 13912 14356 13964 14408
rect 14924 14399 14976 14408
rect 14924 14365 14933 14399
rect 14933 14365 14967 14399
rect 14967 14365 14976 14399
rect 14924 14356 14976 14365
rect 17592 14399 17644 14408
rect 17592 14365 17601 14399
rect 17601 14365 17635 14399
rect 17635 14365 17644 14399
rect 17592 14356 17644 14365
rect 17960 14424 18012 14476
rect 19892 14424 19944 14476
rect 20076 14467 20128 14476
rect 20076 14433 20085 14467
rect 20085 14433 20119 14467
rect 20119 14433 20128 14467
rect 20076 14424 20128 14433
rect 20996 14424 21048 14476
rect 18052 14356 18104 14408
rect 19340 14356 19392 14408
rect 19432 14356 19484 14408
rect 20720 14399 20772 14408
rect 20720 14365 20729 14399
rect 20729 14365 20763 14399
rect 20763 14365 20772 14399
rect 20720 14356 20772 14365
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 22560 14399 22612 14408
rect 22560 14365 22569 14399
rect 22569 14365 22603 14399
rect 22603 14365 22612 14399
rect 22560 14356 22612 14365
rect 23756 14424 23808 14476
rect 23480 14356 23532 14408
rect 1768 14263 1820 14272
rect 1768 14229 1777 14263
rect 1777 14229 1811 14263
rect 1811 14229 1820 14263
rect 1768 14220 1820 14229
rect 4068 14220 4120 14272
rect 6552 14220 6604 14272
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 13820 14288 13872 14340
rect 14004 14288 14056 14340
rect 13636 14263 13688 14272
rect 13636 14229 13645 14263
rect 13645 14229 13679 14263
rect 13679 14229 13688 14263
rect 13636 14220 13688 14229
rect 15016 14220 15068 14272
rect 16580 14288 16632 14340
rect 18604 14288 18656 14340
rect 17776 14220 17828 14272
rect 19340 14220 19392 14272
rect 19432 14220 19484 14272
rect 22376 14220 22428 14272
rect 22468 14220 22520 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1676 14016 1728 14068
rect 6000 14016 6052 14068
rect 7932 14016 7984 14068
rect 9404 14016 9456 14068
rect 10600 14016 10652 14068
rect 13636 14016 13688 14068
rect 2136 13948 2188 14000
rect 2872 13948 2924 14000
rect 4068 13923 4120 13932
rect 4068 13889 4077 13923
rect 4077 13889 4111 13923
rect 4111 13889 4120 13923
rect 4068 13880 4120 13889
rect 7380 13948 7432 14000
rect 5356 13880 5408 13932
rect 6184 13880 6236 13932
rect 7288 13880 7340 13932
rect 8484 13948 8536 14000
rect 8576 13880 8628 13932
rect 9588 13880 9640 13932
rect 9772 13880 9824 13932
rect 10600 13880 10652 13932
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 13820 13948 13872 14000
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 1952 13812 2004 13864
rect 8024 13812 8076 13864
rect 10140 13812 10192 13864
rect 12440 13812 12492 13864
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 14096 13948 14148 14000
rect 15016 13948 15068 14000
rect 18236 14016 18288 14068
rect 19984 14016 20036 14068
rect 14832 13880 14884 13932
rect 17684 13948 17736 14000
rect 28816 14016 28868 14068
rect 23204 13948 23256 14000
rect 5448 13744 5500 13796
rect 3148 13676 3200 13728
rect 5080 13676 5132 13728
rect 8208 13676 8260 13728
rect 10324 13719 10376 13728
rect 10324 13685 10333 13719
rect 10333 13685 10367 13719
rect 10367 13685 10376 13719
rect 10324 13676 10376 13685
rect 11060 13719 11112 13728
rect 11060 13685 11069 13719
rect 11069 13685 11103 13719
rect 11103 13685 11112 13719
rect 11060 13676 11112 13685
rect 11428 13744 11480 13796
rect 11704 13744 11756 13796
rect 12072 13787 12124 13796
rect 12072 13753 12081 13787
rect 12081 13753 12115 13787
rect 12115 13753 12124 13787
rect 12072 13744 12124 13753
rect 13268 13744 13320 13796
rect 13728 13744 13780 13796
rect 14096 13812 14148 13864
rect 15384 13812 15436 13864
rect 16672 13880 16724 13932
rect 19984 13923 20036 13932
rect 15292 13744 15344 13796
rect 16488 13812 16540 13864
rect 18420 13855 18472 13864
rect 18420 13821 18429 13855
rect 18429 13821 18463 13855
rect 18463 13821 18472 13855
rect 18420 13812 18472 13821
rect 19984 13889 19993 13923
rect 19993 13889 20027 13923
rect 20027 13889 20036 13923
rect 19984 13880 20036 13889
rect 22468 13880 22520 13932
rect 20444 13812 20496 13864
rect 22192 13855 22244 13864
rect 22192 13821 22201 13855
rect 22201 13821 22235 13855
rect 22235 13821 22244 13855
rect 22192 13812 22244 13821
rect 24400 13923 24452 13932
rect 24400 13889 24409 13923
rect 24409 13889 24443 13923
rect 24443 13889 24452 13923
rect 24400 13880 24452 13889
rect 34244 13880 34296 13932
rect 16396 13744 16448 13796
rect 22376 13787 22428 13796
rect 22376 13753 22385 13787
rect 22385 13753 22419 13787
rect 22419 13753 22428 13787
rect 22376 13744 22428 13753
rect 34704 13812 34756 13864
rect 12164 13676 12216 13728
rect 14556 13676 14608 13728
rect 16580 13676 16632 13728
rect 38200 13719 38252 13728
rect 38200 13685 38209 13719
rect 38209 13685 38243 13719
rect 38243 13685 38252 13719
rect 38200 13676 38252 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 5816 13472 5868 13524
rect 8116 13472 8168 13524
rect 7564 13404 7616 13456
rect 9680 13472 9732 13524
rect 12900 13472 12952 13524
rect 13268 13472 13320 13524
rect 13636 13472 13688 13524
rect 14556 13472 14608 13524
rect 15384 13472 15436 13524
rect 17776 13472 17828 13524
rect 18604 13515 18656 13524
rect 18604 13481 18613 13515
rect 18613 13481 18647 13515
rect 18647 13481 18656 13515
rect 18604 13472 18656 13481
rect 19984 13472 20036 13524
rect 21640 13472 21692 13524
rect 24400 13472 24452 13524
rect 33416 13515 33468 13524
rect 33416 13481 33425 13515
rect 33425 13481 33459 13515
rect 33459 13481 33468 13515
rect 33416 13472 33468 13481
rect 8760 13404 8812 13456
rect 11152 13404 11204 13456
rect 14464 13404 14516 13456
rect 15660 13404 15712 13456
rect 18236 13404 18288 13456
rect 20076 13447 20128 13456
rect 20076 13413 20085 13447
rect 20085 13413 20119 13447
rect 20119 13413 20128 13447
rect 20076 13404 20128 13413
rect 22376 13404 22428 13456
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 5356 13336 5408 13388
rect 6460 13336 6512 13388
rect 9220 13336 9272 13388
rect 10876 13336 10928 13388
rect 11060 13336 11112 13388
rect 12440 13336 12492 13388
rect 14924 13336 14976 13388
rect 17040 13379 17092 13388
rect 4988 13311 5040 13320
rect 4988 13277 4997 13311
rect 4997 13277 5031 13311
rect 5031 13277 5040 13311
rect 4988 13268 5040 13277
rect 7104 13268 7156 13320
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10416 13268 10468 13320
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 11704 13268 11756 13320
rect 11980 13268 12032 13320
rect 1952 13200 2004 13252
rect 3700 13200 3752 13252
rect 4436 13132 4488 13184
rect 10232 13200 10284 13252
rect 15108 13268 15160 13320
rect 15660 13311 15712 13320
rect 15660 13277 15669 13311
rect 15669 13277 15703 13311
rect 15703 13277 15712 13311
rect 15660 13268 15712 13277
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 17040 13345 17049 13379
rect 17049 13345 17083 13379
rect 17083 13345 17092 13379
rect 17040 13336 17092 13345
rect 20352 13336 20404 13388
rect 20628 13336 20680 13388
rect 23480 13336 23532 13388
rect 24032 13336 24084 13388
rect 17224 13311 17276 13320
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 18328 13268 18380 13320
rect 20720 13268 20772 13320
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 23756 13311 23808 13320
rect 23756 13277 23765 13311
rect 23765 13277 23799 13311
rect 23799 13277 23808 13311
rect 23756 13268 23808 13277
rect 34612 13268 34664 13320
rect 5356 13132 5408 13184
rect 5632 13132 5684 13184
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 10508 13132 10560 13184
rect 10692 13132 10744 13184
rect 11060 13132 11112 13184
rect 11152 13132 11204 13184
rect 11336 13132 11388 13184
rect 11520 13132 11572 13184
rect 11980 13132 12032 13184
rect 12164 13132 12216 13184
rect 12440 13132 12492 13184
rect 12624 13132 12676 13184
rect 13636 13132 13688 13184
rect 17776 13132 17828 13184
rect 19984 13200 20036 13252
rect 22560 13243 22612 13252
rect 22560 13209 22569 13243
rect 22569 13209 22603 13243
rect 22603 13209 22612 13243
rect 22560 13200 22612 13209
rect 21640 13132 21692 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3332 12860 3384 12912
rect 3884 12928 3936 12980
rect 4988 12928 5040 12980
rect 5080 12928 5132 12980
rect 4160 12903 4212 12912
rect 4160 12869 4169 12903
rect 4169 12869 4203 12903
rect 4203 12869 4212 12903
rect 4160 12860 4212 12869
rect 1584 12792 1636 12844
rect 3884 12835 3936 12844
rect 3884 12801 3893 12835
rect 3893 12801 3927 12835
rect 3927 12801 3936 12835
rect 3884 12792 3936 12801
rect 5264 12792 5316 12844
rect 5724 12860 5776 12912
rect 7104 12860 7156 12912
rect 7472 12860 7524 12912
rect 8944 12928 8996 12980
rect 9496 12928 9548 12980
rect 11336 12860 11388 12912
rect 3424 12724 3476 12776
rect 4528 12724 4580 12776
rect 4712 12724 4764 12776
rect 5172 12724 5224 12776
rect 5356 12724 5408 12776
rect 1676 12588 1728 12640
rect 3700 12656 3752 12708
rect 3884 12656 3936 12708
rect 7472 12724 7524 12776
rect 7840 12724 7892 12776
rect 8300 12792 8352 12844
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 8760 12724 8812 12776
rect 10416 12724 10468 12776
rect 11704 12792 11756 12844
rect 11888 12792 11940 12844
rect 12532 12860 12584 12912
rect 15292 12928 15344 12980
rect 15936 12928 15988 12980
rect 16488 12928 16540 12980
rect 18420 12928 18472 12980
rect 19340 12928 19392 12980
rect 20260 12928 20312 12980
rect 12808 12724 12860 12776
rect 13268 12724 13320 12776
rect 14096 12724 14148 12776
rect 14280 12724 14332 12776
rect 15752 12835 15804 12844
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 15752 12792 15804 12801
rect 15108 12724 15160 12776
rect 16120 12724 16172 12776
rect 5724 12588 5776 12640
rect 6828 12588 6880 12640
rect 9588 12588 9640 12640
rect 10692 12588 10744 12640
rect 10876 12656 10928 12708
rect 13636 12656 13688 12708
rect 17040 12860 17092 12912
rect 17868 12860 17920 12912
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 16672 12724 16724 12776
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 18788 12767 18840 12776
rect 18788 12733 18797 12767
rect 18797 12733 18831 12767
rect 18831 12733 18840 12767
rect 18788 12724 18840 12733
rect 19340 12724 19392 12776
rect 20996 12860 21048 12912
rect 21732 12860 21784 12912
rect 18696 12656 18748 12708
rect 22192 12928 22244 12980
rect 22100 12860 22152 12912
rect 23388 12860 23440 12912
rect 31392 12835 31444 12844
rect 31392 12801 31401 12835
rect 31401 12801 31435 12835
rect 31435 12801 31444 12835
rect 31392 12792 31444 12801
rect 23204 12724 23256 12776
rect 23756 12767 23808 12776
rect 23756 12733 23765 12767
rect 23765 12733 23799 12767
rect 23799 12733 23808 12767
rect 23756 12724 23808 12733
rect 22192 12656 22244 12708
rect 23388 12656 23440 12708
rect 16396 12588 16448 12640
rect 19984 12588 20036 12640
rect 20628 12588 20680 12640
rect 22284 12588 22336 12640
rect 23572 12588 23624 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 5816 12384 5868 12436
rect 6828 12384 6880 12436
rect 4344 12316 4396 12368
rect 5264 12316 5316 12368
rect 4804 12248 4856 12300
rect 4988 12248 5040 12300
rect 7196 12316 7248 12368
rect 8116 12316 8168 12368
rect 9956 12384 10008 12436
rect 12440 12384 12492 12436
rect 14924 12384 14976 12436
rect 8024 12248 8076 12300
rect 9496 12248 9548 12300
rect 9864 12248 9916 12300
rect 10416 12248 10468 12300
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 3792 12180 3844 12232
rect 4160 12180 4212 12232
rect 5172 12180 5224 12232
rect 4068 12112 4120 12164
rect 4896 12112 4948 12164
rect 5724 12155 5776 12164
rect 5724 12121 5733 12155
rect 5733 12121 5767 12155
rect 5767 12121 5776 12155
rect 5724 12112 5776 12121
rect 2964 12044 3016 12096
rect 3240 12044 3292 12096
rect 3516 12044 3568 12096
rect 7012 12112 7064 12164
rect 8300 12180 8352 12232
rect 10324 12180 10376 12232
rect 11612 12316 11664 12368
rect 11888 12248 11940 12300
rect 12624 12291 12676 12300
rect 12624 12257 12633 12291
rect 12633 12257 12667 12291
rect 12667 12257 12676 12291
rect 12624 12248 12676 12257
rect 12808 12248 12860 12300
rect 12992 12248 13044 12300
rect 11520 12180 11572 12232
rect 12440 12180 12492 12232
rect 16672 12316 16724 12368
rect 18328 12384 18380 12436
rect 19432 12384 19484 12436
rect 20168 12384 20220 12436
rect 20352 12316 20404 12368
rect 20628 12316 20680 12368
rect 16304 12291 16356 12300
rect 16304 12257 16313 12291
rect 16313 12257 16347 12291
rect 16347 12257 16356 12291
rect 16304 12248 16356 12257
rect 16580 12291 16632 12300
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 18236 12248 18288 12300
rect 23480 12316 23532 12368
rect 24032 12291 24084 12300
rect 24032 12257 24041 12291
rect 24041 12257 24075 12291
rect 24075 12257 24084 12291
rect 24032 12248 24084 12257
rect 14648 12180 14700 12232
rect 16120 12180 16172 12232
rect 18420 12180 18472 12232
rect 19984 12180 20036 12232
rect 21548 12223 21600 12232
rect 9588 12112 9640 12164
rect 9680 12112 9732 12164
rect 7196 12087 7248 12096
rect 7196 12053 7205 12087
rect 7205 12053 7239 12087
rect 7239 12053 7248 12087
rect 7196 12044 7248 12053
rect 7288 12044 7340 12096
rect 12256 12112 12308 12164
rect 12440 12044 12492 12096
rect 13268 12155 13320 12164
rect 13268 12121 13277 12155
rect 13277 12121 13311 12155
rect 13311 12121 13320 12155
rect 13268 12112 13320 12121
rect 13452 12112 13504 12164
rect 15200 12112 15252 12164
rect 16580 12112 16632 12164
rect 18512 12112 18564 12164
rect 21548 12189 21557 12223
rect 21557 12189 21591 12223
rect 21591 12189 21600 12223
rect 21548 12180 21600 12189
rect 21732 12180 21784 12232
rect 24124 12180 24176 12232
rect 24676 12112 24728 12164
rect 14004 12044 14056 12096
rect 14740 12044 14792 12096
rect 15568 12044 15620 12096
rect 16304 12044 16356 12096
rect 20444 12044 20496 12096
rect 21180 12044 21232 12096
rect 23848 12044 23900 12096
rect 36452 12044 36504 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2964 11840 3016 11892
rect 2044 11772 2096 11824
rect 4068 11772 4120 11824
rect 5080 11840 5132 11892
rect 5356 11840 5408 11892
rect 5816 11840 5868 11892
rect 6276 11772 6328 11824
rect 1952 11704 2004 11756
rect 4252 11704 4304 11756
rect 5080 11704 5132 11756
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 6920 11772 6972 11824
rect 7288 11772 7340 11824
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 7012 11704 7064 11756
rect 7932 11704 7984 11756
rect 1676 11636 1728 11688
rect 3056 11636 3108 11688
rect 3608 11636 3660 11688
rect 4804 11679 4856 11688
rect 4804 11645 4813 11679
rect 4813 11645 4847 11679
rect 4847 11645 4856 11679
rect 4804 11636 4856 11645
rect 5724 11636 5776 11688
rect 6092 11636 6144 11688
rect 6460 11636 6512 11688
rect 8668 11636 8720 11688
rect 9588 11636 9640 11688
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 12440 11840 12492 11892
rect 12624 11840 12676 11892
rect 13176 11840 13228 11892
rect 14188 11840 14240 11892
rect 13820 11772 13872 11824
rect 15016 11840 15068 11892
rect 16580 11840 16632 11892
rect 17224 11840 17276 11892
rect 17960 11840 18012 11892
rect 20076 11840 20128 11892
rect 21732 11840 21784 11892
rect 22100 11883 22152 11892
rect 22100 11849 22109 11883
rect 22109 11849 22143 11883
rect 22143 11849 22152 11883
rect 22100 11840 22152 11849
rect 22560 11840 22612 11892
rect 24676 11883 24728 11892
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 34244 11883 34296 11892
rect 34244 11849 34253 11883
rect 34253 11849 34287 11883
rect 34287 11849 34296 11883
rect 34244 11840 34296 11849
rect 34612 11840 34664 11892
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 14740 11704 14792 11756
rect 10232 11636 10284 11688
rect 10784 11636 10836 11688
rect 13360 11679 13412 11688
rect 13360 11645 13369 11679
rect 13369 11645 13403 11679
rect 13403 11645 13412 11679
rect 13360 11636 13412 11645
rect 13452 11636 13504 11688
rect 4344 11568 4396 11620
rect 6736 11568 6788 11620
rect 3608 11500 3660 11552
rect 5080 11500 5132 11552
rect 7656 11500 7708 11552
rect 14188 11568 14240 11620
rect 10324 11500 10376 11552
rect 10416 11500 10468 11552
rect 11980 11500 12032 11552
rect 14096 11500 14148 11552
rect 14556 11636 14608 11688
rect 15752 11679 15804 11688
rect 15752 11645 15761 11679
rect 15761 11645 15795 11679
rect 15795 11645 15804 11679
rect 15752 11636 15804 11645
rect 14832 11568 14884 11620
rect 17776 11747 17828 11756
rect 17776 11713 17785 11747
rect 17785 11713 17819 11747
rect 17819 11713 17828 11747
rect 17776 11704 17828 11713
rect 18696 11704 18748 11756
rect 19432 11704 19484 11756
rect 21180 11772 21232 11824
rect 24584 11772 24636 11824
rect 20536 11704 20588 11756
rect 20904 11704 20956 11756
rect 21548 11704 21600 11756
rect 20168 11679 20220 11688
rect 20168 11645 20177 11679
rect 20177 11645 20211 11679
rect 20211 11645 20220 11679
rect 20168 11636 20220 11645
rect 20720 11636 20772 11688
rect 20352 11568 20404 11620
rect 22836 11704 22888 11756
rect 24216 11704 24268 11756
rect 30380 11704 30432 11756
rect 38292 11747 38344 11756
rect 38292 11713 38301 11747
rect 38301 11713 38335 11747
rect 38335 11713 38344 11747
rect 38292 11704 38344 11713
rect 23664 11568 23716 11620
rect 23756 11568 23808 11620
rect 24308 11568 24360 11620
rect 17592 11500 17644 11552
rect 19524 11543 19576 11552
rect 19524 11509 19533 11543
rect 19533 11509 19567 11543
rect 19567 11509 19576 11543
rect 19524 11500 19576 11509
rect 20444 11500 20496 11552
rect 20720 11500 20772 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3608 11228 3660 11280
rect 7196 11296 7248 11348
rect 9128 11296 9180 11348
rect 13360 11296 13412 11348
rect 13912 11296 13964 11348
rect 14280 11296 14332 11348
rect 15108 11296 15160 11348
rect 16304 11296 16356 11348
rect 16488 11296 16540 11348
rect 18420 11339 18472 11348
rect 18420 11305 18429 11339
rect 18429 11305 18463 11339
rect 18463 11305 18472 11339
rect 18420 11296 18472 11305
rect 19340 11296 19392 11348
rect 24216 11296 24268 11348
rect 24584 11339 24636 11348
rect 24584 11305 24593 11339
rect 24593 11305 24627 11339
rect 24627 11305 24636 11339
rect 24584 11296 24636 11305
rect 1584 11092 1636 11144
rect 3608 11024 3660 11076
rect 2780 10956 2832 11008
rect 3332 10956 3384 11008
rect 4988 11160 5040 11212
rect 6736 11160 6788 11212
rect 7564 11160 7616 11212
rect 7656 11160 7708 11212
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 9036 11160 9088 11212
rect 11520 11228 11572 11280
rect 13084 11228 13136 11280
rect 15936 11228 15988 11280
rect 10416 11160 10468 11212
rect 10968 11160 11020 11212
rect 13912 11160 13964 11212
rect 15844 11160 15896 11212
rect 5540 11092 5592 11144
rect 9312 11092 9364 11144
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12532 11092 12584 11101
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 14832 11135 14884 11144
rect 14832 11101 14841 11135
rect 14841 11101 14875 11135
rect 14875 11101 14884 11135
rect 14832 11092 14884 11101
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 18512 11092 18564 11144
rect 19340 11160 19392 11212
rect 19524 11160 19576 11212
rect 24124 11160 24176 11212
rect 24308 11160 24360 11212
rect 20812 11092 20864 11144
rect 22836 11135 22888 11144
rect 22836 11101 22845 11135
rect 22845 11101 22879 11135
rect 22879 11101 22888 11135
rect 22836 11092 22888 11101
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 4436 11067 4488 11076
rect 4436 11033 4445 11067
rect 4445 11033 4479 11067
rect 4479 11033 4488 11067
rect 4436 11024 4488 11033
rect 7012 11024 7064 11076
rect 9128 11024 9180 11076
rect 10416 11067 10468 11076
rect 10416 11033 10425 11067
rect 10425 11033 10459 11067
rect 10459 11033 10468 11067
rect 10416 11024 10468 11033
rect 11704 11024 11756 11076
rect 17776 11067 17828 11076
rect 17776 11033 17785 11067
rect 17785 11033 17819 11067
rect 17819 11033 17828 11067
rect 17776 11024 17828 11033
rect 30840 11024 30892 11076
rect 9680 10956 9732 11008
rect 9772 10956 9824 11008
rect 12164 10956 12216 11008
rect 13176 10956 13228 11008
rect 15568 10956 15620 11008
rect 16764 10956 16816 11008
rect 17224 10956 17276 11008
rect 20720 10956 20772 11008
rect 21088 10956 21140 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1768 10752 1820 10804
rect 4804 10752 4856 10804
rect 8392 10752 8444 10804
rect 9128 10752 9180 10804
rect 2780 10684 2832 10736
rect 3148 10684 3200 10736
rect 5448 10684 5500 10736
rect 7104 10684 7156 10736
rect 14464 10752 14516 10804
rect 15752 10752 15804 10804
rect 16120 10752 16172 10804
rect 18604 10752 18656 10804
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 20168 10752 20220 10804
rect 20812 10795 20864 10804
rect 20812 10761 20821 10795
rect 20821 10761 20855 10795
rect 20855 10761 20864 10795
rect 20812 10752 20864 10761
rect 20996 10752 21048 10804
rect 23204 10752 23256 10804
rect 23848 10752 23900 10804
rect 24768 10752 24820 10804
rect 30380 10752 30432 10804
rect 10692 10684 10744 10736
rect 12440 10684 12492 10736
rect 13452 10684 13504 10736
rect 16856 10684 16908 10736
rect 16948 10684 17000 10736
rect 20444 10684 20496 10736
rect 2136 10616 2188 10668
rect 2320 10616 2372 10668
rect 5172 10659 5224 10668
rect 5172 10625 5181 10659
rect 5181 10625 5215 10659
rect 5215 10625 5224 10659
rect 5172 10616 5224 10625
rect 6000 10659 6052 10668
rect 6000 10625 6009 10659
rect 6009 10625 6043 10659
rect 6043 10625 6052 10659
rect 6000 10616 6052 10625
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 8852 10616 8904 10668
rect 9128 10616 9180 10668
rect 1584 10480 1636 10532
rect 3148 10591 3200 10600
rect 3148 10557 3157 10591
rect 3157 10557 3191 10591
rect 3191 10557 3200 10591
rect 3148 10548 3200 10557
rect 8760 10548 8812 10600
rect 9036 10548 9088 10600
rect 4436 10412 4488 10464
rect 4804 10412 4856 10464
rect 5080 10412 5132 10464
rect 8852 10480 8904 10532
rect 11152 10523 11204 10532
rect 11152 10489 11161 10523
rect 11161 10489 11195 10523
rect 11195 10489 11204 10523
rect 13176 10548 13228 10600
rect 15108 10616 15160 10668
rect 16028 10616 16080 10668
rect 16396 10616 16448 10668
rect 20352 10616 20404 10668
rect 20996 10659 21048 10668
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 21088 10616 21140 10668
rect 23572 10659 23624 10668
rect 23572 10625 23581 10659
rect 23581 10625 23615 10659
rect 23615 10625 23624 10659
rect 23572 10616 23624 10625
rect 23664 10616 23716 10668
rect 24860 10616 24912 10668
rect 30840 10616 30892 10668
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 16856 10591 16908 10600
rect 16856 10557 16865 10591
rect 16865 10557 16899 10591
rect 16899 10557 16908 10591
rect 16856 10548 16908 10557
rect 11152 10480 11204 10489
rect 9680 10455 9732 10464
rect 9680 10421 9704 10455
rect 9704 10421 9732 10455
rect 9680 10412 9732 10421
rect 10416 10412 10468 10464
rect 17224 10523 17276 10532
rect 17224 10489 17233 10523
rect 17233 10489 17267 10523
rect 17267 10489 17276 10523
rect 17224 10480 17276 10489
rect 18604 10548 18656 10600
rect 19156 10480 19208 10532
rect 24768 10480 24820 10532
rect 13636 10412 13688 10464
rect 15844 10412 15896 10464
rect 38016 10412 38068 10464
rect 38200 10455 38252 10464
rect 38200 10421 38209 10455
rect 38209 10421 38243 10455
rect 38243 10421 38252 10455
rect 38200 10412 38252 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 5356 10208 5408 10260
rect 5080 10140 5132 10192
rect 3976 10115 4028 10124
rect 3976 10081 3985 10115
rect 3985 10081 4019 10115
rect 4019 10081 4028 10115
rect 3976 10072 4028 10081
rect 4068 10072 4120 10124
rect 1584 10004 1636 10056
rect 6552 10208 6604 10260
rect 7380 10208 7432 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 12072 10208 12124 10260
rect 13084 10208 13136 10260
rect 13268 10208 13320 10260
rect 13820 10208 13872 10260
rect 14464 10208 14516 10260
rect 14648 10251 14700 10260
rect 14648 10217 14657 10251
rect 14657 10217 14691 10251
rect 14691 10217 14700 10251
rect 14648 10208 14700 10217
rect 15108 10208 15160 10260
rect 15568 10208 15620 10260
rect 16672 10208 16724 10260
rect 18604 10251 18656 10260
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 20996 10208 21048 10260
rect 23480 10251 23532 10260
rect 23480 10217 23489 10251
rect 23489 10217 23523 10251
rect 23523 10217 23532 10251
rect 23480 10208 23532 10217
rect 11888 10183 11940 10192
rect 6736 10072 6788 10124
rect 9036 10072 9088 10124
rect 11888 10149 11897 10183
rect 11897 10149 11931 10183
rect 11931 10149 11940 10183
rect 11888 10140 11940 10149
rect 12808 10072 12860 10124
rect 13176 10072 13228 10124
rect 8944 10004 8996 10056
rect 9312 10004 9364 10056
rect 9404 10004 9456 10056
rect 11980 10004 12032 10056
rect 13820 10004 13872 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 5540 9936 5592 9988
rect 6460 9936 6512 9988
rect 6920 9936 6972 9988
rect 2596 9868 2648 9920
rect 8300 9936 8352 9988
rect 10140 9936 10192 9988
rect 11704 9936 11756 9988
rect 15936 10140 15988 10192
rect 16212 10140 16264 10192
rect 18788 10140 18840 10192
rect 16488 10072 16540 10124
rect 19340 10072 19392 10124
rect 20260 10140 20312 10192
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 20260 10004 20312 10056
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 23296 10047 23348 10056
rect 8668 9868 8720 9920
rect 9128 9868 9180 9920
rect 16764 9936 16816 9988
rect 17132 9979 17184 9988
rect 17132 9945 17141 9979
rect 17141 9945 17175 9979
rect 17175 9945 17184 9979
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 36912 10004 36964 10056
rect 17132 9936 17184 9945
rect 29552 9936 29604 9988
rect 14096 9868 14148 9920
rect 14372 9868 14424 9920
rect 16120 9868 16172 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 3424 9596 3476 9648
rect 4896 9596 4948 9648
rect 7288 9664 7340 9716
rect 8852 9664 8904 9716
rect 7196 9596 7248 9648
rect 8208 9596 8260 9648
rect 8576 9596 8628 9648
rect 9588 9596 9640 9648
rect 11704 9664 11756 9716
rect 12072 9596 12124 9648
rect 12256 9639 12308 9648
rect 12256 9605 12265 9639
rect 12265 9605 12299 9639
rect 12299 9605 12308 9639
rect 12256 9596 12308 9605
rect 12808 9596 12860 9648
rect 14280 9664 14332 9716
rect 18328 9664 18380 9716
rect 19064 9664 19116 9716
rect 21548 9664 21600 9716
rect 23296 9707 23348 9716
rect 23296 9673 23305 9707
rect 23305 9673 23339 9707
rect 23339 9673 23348 9707
rect 23296 9664 23348 9673
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 10600 9528 10652 9580
rect 14372 9596 14424 9648
rect 14648 9596 14700 9648
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 3976 9460 4028 9512
rect 8484 9460 8536 9512
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 12532 9460 12584 9512
rect 1860 9324 1912 9376
rect 10416 9392 10468 9444
rect 12348 9392 12400 9444
rect 4528 9324 4580 9376
rect 5080 9324 5132 9376
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 6736 9324 6788 9376
rect 9036 9324 9088 9376
rect 9312 9324 9364 9376
rect 11152 9324 11204 9376
rect 11428 9324 11480 9376
rect 13268 9324 13320 9376
rect 13452 9324 13504 9376
rect 14832 9528 14884 9580
rect 15016 9460 15068 9512
rect 18052 9596 18104 9648
rect 17592 9528 17644 9580
rect 15292 9460 15344 9512
rect 17040 9460 17092 9512
rect 17224 9460 17276 9512
rect 22192 9460 22244 9512
rect 28264 9392 28316 9444
rect 15200 9324 15252 9376
rect 18788 9324 18840 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1952 9120 2004 9172
rect 5724 9163 5776 9172
rect 3332 9095 3384 9104
rect 3332 9061 3341 9095
rect 3341 9061 3375 9095
rect 3375 9061 3384 9095
rect 3332 9052 3384 9061
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 5908 9120 5960 9172
rect 9220 9120 9272 9172
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 3976 9027 4028 9036
rect 3976 8993 3985 9027
rect 3985 8993 4019 9027
rect 4019 8993 4028 9027
rect 3976 8984 4028 8993
rect 5264 8984 5316 9036
rect 8484 9052 8536 9104
rect 11060 9120 11112 9172
rect 14648 9120 14700 9172
rect 15752 9120 15804 9172
rect 11612 9052 11664 9104
rect 9864 8984 9916 9036
rect 10324 9027 10376 9036
rect 10324 8993 10333 9027
rect 10333 8993 10367 9027
rect 10367 8993 10376 9027
rect 10324 8984 10376 8993
rect 13544 9052 13596 9104
rect 15476 9052 15528 9104
rect 16856 9120 16908 9172
rect 17408 9120 17460 9172
rect 18052 9163 18104 9172
rect 18052 9129 18061 9163
rect 18061 9129 18095 9163
rect 18095 9129 18104 9163
rect 18052 9120 18104 9129
rect 21824 9120 21876 9172
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 6736 8916 6788 8968
rect 8208 8916 8260 8968
rect 8760 8916 8812 8968
rect 8944 8916 8996 8968
rect 9772 8916 9824 8968
rect 11888 8916 11940 8968
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 16212 9027 16264 9036
rect 16212 8993 16221 9027
rect 16221 8993 16255 9027
rect 16255 8993 16264 9027
rect 16212 8984 16264 8993
rect 16304 8984 16356 9036
rect 20076 8984 20128 9036
rect 14648 8916 14700 8968
rect 15384 8959 15436 8968
rect 15384 8925 15393 8959
rect 15393 8925 15427 8959
rect 15427 8925 15436 8959
rect 15384 8916 15436 8925
rect 15476 8916 15528 8968
rect 1860 8891 1912 8900
rect 1860 8857 1869 8891
rect 1869 8857 1903 8891
rect 1903 8857 1912 8891
rect 1860 8848 1912 8857
rect 3516 8848 3568 8900
rect 4804 8848 4856 8900
rect 3148 8780 3200 8832
rect 6092 8780 6144 8832
rect 10416 8848 10468 8900
rect 11336 8848 11388 8900
rect 14280 8848 14332 8900
rect 20996 8916 21048 8968
rect 28448 8916 28500 8968
rect 38016 8959 38068 8968
rect 38016 8925 38025 8959
rect 38025 8925 38059 8959
rect 38059 8925 38068 8959
rect 38016 8916 38068 8925
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 8760 8780 8812 8832
rect 9588 8780 9640 8832
rect 9864 8780 9916 8832
rect 13544 8780 13596 8832
rect 13820 8780 13872 8832
rect 16672 8780 16724 8832
rect 17316 8780 17368 8832
rect 17960 8780 18012 8832
rect 20352 8780 20404 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 3332 8440 3384 8492
rect 3884 8576 3936 8628
rect 4988 8508 5040 8560
rect 5908 8508 5960 8560
rect 1584 8372 1636 8424
rect 2872 8372 2924 8424
rect 4620 8440 4672 8492
rect 6092 8576 6144 8628
rect 3700 8236 3752 8288
rect 8392 8440 8444 8492
rect 6736 8372 6788 8424
rect 10140 8576 10192 8628
rect 10508 8576 10560 8628
rect 15016 8619 15068 8628
rect 9036 8440 9088 8492
rect 9772 8508 9824 8560
rect 10048 8508 10100 8560
rect 12256 8508 12308 8560
rect 13728 8508 13780 8560
rect 15016 8585 15025 8619
rect 15025 8585 15059 8619
rect 15059 8585 15068 8619
rect 15016 8576 15068 8585
rect 18236 8576 18288 8628
rect 17316 8551 17368 8560
rect 17316 8517 17325 8551
rect 17325 8517 17359 8551
rect 17359 8517 17368 8551
rect 17316 8508 17368 8517
rect 17408 8551 17460 8560
rect 17408 8517 17417 8551
rect 17417 8517 17451 8551
rect 17451 8517 17460 8551
rect 18512 8551 18564 8560
rect 17408 8508 17460 8517
rect 18512 8517 18521 8551
rect 18521 8517 18555 8551
rect 18555 8517 18564 8551
rect 18512 8508 18564 8517
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 6000 8304 6052 8356
rect 10968 8372 11020 8424
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 13452 8415 13504 8424
rect 13452 8381 13461 8415
rect 13461 8381 13495 8415
rect 13495 8381 13504 8415
rect 13452 8372 13504 8381
rect 13544 8372 13596 8424
rect 9220 8304 9272 8356
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 15752 8372 15804 8424
rect 16396 8372 16448 8424
rect 24860 8576 24912 8628
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 22008 8440 22060 8492
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 20720 8415 20772 8424
rect 16028 8304 16080 8356
rect 20720 8381 20729 8415
rect 20729 8381 20763 8415
rect 20763 8381 20772 8415
rect 20720 8372 20772 8381
rect 18052 8304 18104 8356
rect 21088 8304 21140 8356
rect 22100 8304 22152 8356
rect 30012 8304 30064 8356
rect 9312 8236 9364 8288
rect 9588 8236 9640 8288
rect 10140 8236 10192 8288
rect 11060 8236 11112 8288
rect 12440 8236 12492 8288
rect 12532 8236 12584 8288
rect 14004 8236 14056 8288
rect 16120 8236 16172 8288
rect 18880 8236 18932 8288
rect 20628 8236 20680 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1860 8032 1912 8084
rect 2596 8032 2648 8084
rect 3792 7964 3844 8016
rect 5172 8032 5224 8084
rect 11060 8032 11112 8084
rect 12716 8032 12768 8084
rect 17132 8032 17184 8084
rect 17408 8075 17460 8084
rect 17408 8041 17417 8075
rect 17417 8041 17451 8075
rect 17451 8041 17460 8075
rect 17408 8032 17460 8041
rect 17500 8032 17552 8084
rect 19432 8032 19484 8084
rect 20720 8032 20772 8084
rect 7288 8007 7340 8016
rect 7288 7973 7297 8007
rect 7297 7973 7331 8007
rect 7331 7973 7340 8007
rect 7288 7964 7340 7973
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 3608 7896 3660 7948
rect 3884 7828 3936 7880
rect 6460 7896 6512 7948
rect 8300 7896 8352 7948
rect 9312 7896 9364 7948
rect 4068 7760 4120 7812
rect 4988 7828 5040 7880
rect 9220 7828 9272 7880
rect 9772 7896 9824 7948
rect 11428 7964 11480 8016
rect 12072 7896 12124 7948
rect 12716 7896 12768 7948
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 16396 7896 16448 7948
rect 9956 7828 10008 7880
rect 11428 7828 11480 7880
rect 11704 7828 11756 7880
rect 12440 7828 12492 7880
rect 5356 7760 5408 7812
rect 5724 7760 5776 7812
rect 8300 7760 8352 7812
rect 10232 7760 10284 7812
rect 10324 7803 10376 7812
rect 10324 7769 10333 7803
rect 10333 7769 10367 7803
rect 10367 7769 10376 7803
rect 10324 7760 10376 7769
rect 3332 7735 3384 7744
rect 3332 7701 3341 7735
rect 3341 7701 3375 7735
rect 3375 7701 3384 7735
rect 3332 7692 3384 7701
rect 8208 7692 8260 7744
rect 8576 7692 8628 7744
rect 9036 7692 9088 7744
rect 9312 7692 9364 7744
rect 12716 7760 12768 7812
rect 12072 7692 12124 7744
rect 13176 7828 13228 7880
rect 13820 7828 13872 7880
rect 15016 7828 15068 7880
rect 15660 7760 15712 7812
rect 16948 7828 17000 7880
rect 18328 7964 18380 8016
rect 20628 7871 20680 7880
rect 17500 7760 17552 7812
rect 17684 7760 17736 7812
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 20812 7828 20864 7880
rect 30196 7828 30248 7880
rect 20536 7760 20588 7812
rect 22468 7760 22520 7812
rect 13636 7692 13688 7744
rect 16580 7692 16632 7744
rect 16856 7692 16908 7744
rect 17592 7692 17644 7744
rect 18328 7692 18380 7744
rect 22192 7692 22244 7744
rect 22652 7692 22704 7744
rect 23296 7692 23348 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1860 7463 1912 7472
rect 1860 7429 1869 7463
rect 1869 7429 1903 7463
rect 1903 7429 1912 7463
rect 1860 7420 1912 7429
rect 6552 7488 6604 7540
rect 6920 7488 6972 7540
rect 7748 7420 7800 7472
rect 5356 7352 5408 7404
rect 8852 7488 8904 7540
rect 9036 7488 9088 7540
rect 10600 7488 10652 7540
rect 12992 7488 13044 7540
rect 13452 7488 13504 7540
rect 8116 7420 8168 7472
rect 11060 7420 11112 7472
rect 11980 7463 12032 7472
rect 11980 7429 11989 7463
rect 11989 7429 12023 7463
rect 12023 7429 12032 7463
rect 11980 7420 12032 7429
rect 14004 7420 14056 7472
rect 15200 7420 15252 7472
rect 16212 7488 16264 7540
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 17040 7488 17092 7540
rect 18236 7531 18288 7540
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 18880 7531 18932 7540
rect 18880 7497 18889 7531
rect 18889 7497 18923 7531
rect 18923 7497 18932 7531
rect 18880 7488 18932 7497
rect 29552 7531 29604 7540
rect 29552 7497 29561 7531
rect 29561 7497 29595 7531
rect 29595 7497 29604 7531
rect 29552 7488 29604 7497
rect 33876 7531 33928 7540
rect 33876 7497 33885 7531
rect 33885 7497 33919 7531
rect 33919 7497 33928 7531
rect 33876 7488 33928 7497
rect 36912 7488 36964 7540
rect 18328 7420 18380 7472
rect 18604 7420 18656 7472
rect 20996 7420 21048 7472
rect 22192 7463 22244 7472
rect 22192 7429 22201 7463
rect 22201 7429 22235 7463
rect 22235 7429 22244 7463
rect 22192 7420 22244 7429
rect 23296 7463 23348 7472
rect 23296 7429 23305 7463
rect 23305 7429 23339 7463
rect 23339 7429 23348 7463
rect 23296 7420 23348 7429
rect 23388 7463 23440 7472
rect 23388 7429 23397 7463
rect 23397 7429 23431 7463
rect 23431 7429 23440 7463
rect 23388 7420 23440 7429
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 10324 7352 10376 7404
rect 10968 7352 11020 7404
rect 14924 7352 14976 7404
rect 15844 7352 15896 7404
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 3884 7284 3936 7336
rect 4620 7284 4672 7336
rect 5448 7284 5500 7336
rect 6736 7284 6788 7336
rect 8208 7284 8260 7336
rect 10508 7327 10560 7336
rect 7288 7259 7340 7268
rect 7288 7225 7297 7259
rect 7297 7225 7331 7259
rect 7331 7225 7340 7259
rect 7288 7216 7340 7225
rect 10508 7293 10517 7327
rect 10517 7293 10551 7327
rect 10551 7293 10560 7327
rect 10508 7284 10560 7293
rect 11152 7216 11204 7268
rect 8944 7148 8996 7200
rect 11704 7148 11756 7200
rect 13452 7284 13504 7336
rect 16764 7352 16816 7404
rect 17868 7352 17920 7404
rect 17040 7284 17092 7336
rect 19892 7352 19944 7404
rect 20076 7352 20128 7404
rect 19340 7284 19392 7336
rect 22100 7327 22152 7336
rect 22100 7293 22109 7327
rect 22109 7293 22143 7327
rect 22143 7293 22152 7327
rect 22100 7284 22152 7293
rect 29552 7284 29604 7336
rect 35716 7352 35768 7404
rect 38292 7395 38344 7404
rect 38292 7361 38301 7395
rect 38301 7361 38335 7395
rect 38335 7361 38344 7395
rect 38292 7352 38344 7361
rect 34704 7284 34756 7336
rect 16488 7216 16540 7268
rect 16948 7216 17000 7268
rect 17592 7216 17644 7268
rect 13452 7191 13504 7200
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 17868 7148 17920 7200
rect 20996 7148 21048 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3332 6944 3384 6996
rect 4620 6944 4672 6996
rect 7748 6944 7800 6996
rect 10048 6944 10100 6996
rect 13452 6944 13504 6996
rect 13636 6944 13688 6996
rect 16212 6944 16264 6996
rect 17500 6944 17552 6996
rect 23388 6944 23440 6996
rect 1584 6740 1636 6792
rect 3884 6808 3936 6860
rect 4988 6808 5040 6860
rect 6736 6808 6788 6860
rect 7104 6808 7156 6860
rect 9772 6808 9824 6860
rect 10324 6851 10376 6860
rect 10324 6817 10333 6851
rect 10333 6817 10367 6851
rect 10367 6817 10376 6851
rect 10324 6808 10376 6817
rect 12072 6876 12124 6928
rect 14556 6876 14608 6928
rect 11336 6808 11388 6860
rect 5540 6740 5592 6792
rect 5724 6740 5776 6792
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 2228 6672 2280 6724
rect 5264 6672 5316 6724
rect 2320 6604 2372 6656
rect 4160 6604 4212 6656
rect 5724 6604 5776 6656
rect 7288 6604 7340 6656
rect 7564 6672 7616 6724
rect 7840 6604 7892 6656
rect 8116 6604 8168 6656
rect 10232 6672 10284 6724
rect 10508 6672 10560 6724
rect 11152 6672 11204 6724
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 9496 6604 9548 6656
rect 13176 6808 13228 6860
rect 15384 6808 15436 6860
rect 19432 6876 19484 6928
rect 20444 6876 20496 6928
rect 20996 6851 21048 6860
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 16856 6740 16908 6792
rect 16948 6783 17000 6792
rect 16948 6749 16957 6783
rect 16957 6749 16991 6783
rect 16991 6749 17000 6783
rect 16948 6740 17000 6749
rect 17868 6740 17920 6792
rect 18052 6740 18104 6792
rect 18604 6740 18656 6792
rect 11980 6672 12032 6724
rect 14372 6672 14424 6724
rect 19984 6740 20036 6792
rect 20996 6817 21005 6851
rect 21005 6817 21039 6851
rect 21039 6817 21048 6851
rect 20996 6808 21048 6817
rect 22100 6808 22152 6860
rect 24584 6808 24636 6860
rect 22652 6783 22704 6792
rect 20720 6672 20772 6724
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 31208 6672 31260 6724
rect 12072 6647 12124 6656
rect 12072 6613 12081 6647
rect 12081 6613 12115 6647
rect 12115 6613 12124 6647
rect 12072 6604 12124 6613
rect 13084 6604 13136 6656
rect 15016 6604 15068 6656
rect 17040 6604 17092 6656
rect 21456 6604 21508 6656
rect 33876 6740 33928 6792
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2504 6400 2556 6452
rect 2688 6400 2740 6452
rect 4160 6332 4212 6384
rect 1584 6196 1636 6248
rect 2780 6196 2832 6248
rect 7104 6332 7156 6384
rect 7288 6375 7340 6384
rect 7288 6341 7297 6375
rect 7297 6341 7331 6375
rect 7331 6341 7340 6375
rect 7288 6332 7340 6341
rect 9864 6400 9916 6452
rect 11980 6400 12032 6452
rect 12716 6400 12768 6452
rect 16396 6400 16448 6452
rect 18696 6400 18748 6452
rect 19248 6400 19300 6452
rect 21640 6400 21692 6452
rect 13912 6332 13964 6384
rect 14280 6332 14332 6384
rect 17040 6375 17092 6384
rect 17040 6341 17049 6375
rect 17049 6341 17083 6375
rect 17083 6341 17092 6375
rect 17040 6332 17092 6341
rect 20076 6375 20128 6384
rect 20076 6341 20085 6375
rect 20085 6341 20119 6375
rect 20119 6341 20128 6375
rect 20076 6332 20128 6341
rect 4620 6196 4672 6248
rect 5448 6196 5500 6248
rect 6460 6264 6512 6316
rect 8024 6264 8076 6316
rect 11060 6264 11112 6316
rect 11428 6264 11480 6316
rect 15292 6264 15344 6316
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 17684 6264 17736 6316
rect 19340 6307 19392 6316
rect 19340 6273 19349 6307
rect 19349 6273 19383 6307
rect 19383 6273 19392 6307
rect 19340 6264 19392 6273
rect 19984 6307 20036 6316
rect 19984 6273 19993 6307
rect 19993 6273 20027 6307
rect 20027 6273 20036 6307
rect 20628 6307 20680 6316
rect 19984 6264 20036 6273
rect 20628 6273 20637 6307
rect 20637 6273 20671 6307
rect 20671 6273 20680 6307
rect 20628 6264 20680 6273
rect 24216 6264 24268 6316
rect 29552 6307 29604 6316
rect 29552 6273 29561 6307
rect 29561 6273 29595 6307
rect 29595 6273 29604 6307
rect 29552 6264 29604 6273
rect 5632 6128 5684 6180
rect 2412 6060 2464 6112
rect 6736 6196 6788 6248
rect 10048 6196 10100 6248
rect 10324 6196 10376 6248
rect 11980 6239 12032 6248
rect 6828 6060 6880 6112
rect 10876 6128 10928 6180
rect 11612 6128 11664 6180
rect 8760 6060 8812 6112
rect 9404 6060 9456 6112
rect 11704 6060 11756 6112
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 13912 6239 13964 6248
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 16488 6196 16540 6248
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 17224 6196 17276 6205
rect 19156 6196 19208 6248
rect 21456 6196 21508 6248
rect 13452 6171 13504 6180
rect 13452 6137 13461 6171
rect 13461 6137 13495 6171
rect 13495 6137 13504 6171
rect 13452 6128 13504 6137
rect 15292 6128 15344 6180
rect 21364 6171 21416 6180
rect 13820 6060 13872 6112
rect 16028 6060 16080 6112
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 21364 6137 21373 6171
rect 21373 6137 21407 6171
rect 21407 6137 21416 6171
rect 21364 6128 21416 6137
rect 29644 6103 29696 6112
rect 29644 6069 29653 6103
rect 29653 6069 29687 6103
rect 29687 6069 29696 6103
rect 29644 6060 29696 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4068 5856 4120 5908
rect 6552 5856 6604 5908
rect 2964 5788 3016 5840
rect 8576 5856 8628 5908
rect 9312 5899 9364 5908
rect 9312 5865 9321 5899
rect 9321 5865 9355 5899
rect 9355 5865 9364 5899
rect 9312 5856 9364 5865
rect 9588 5856 9640 5908
rect 10784 5856 10836 5908
rect 10968 5856 11020 5908
rect 11244 5856 11296 5908
rect 11888 5856 11940 5908
rect 12072 5856 12124 5908
rect 19432 5856 19484 5908
rect 20904 5856 20956 5908
rect 21272 5856 21324 5908
rect 22100 5899 22152 5908
rect 22100 5865 22109 5899
rect 22109 5865 22143 5899
rect 22143 5865 22152 5899
rect 22100 5856 22152 5865
rect 6552 5720 6604 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 4068 5652 4120 5704
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 4988 5652 5040 5704
rect 8024 5652 8076 5704
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 6736 5584 6788 5636
rect 7288 5584 7340 5636
rect 8484 5652 8536 5704
rect 9128 5652 9180 5704
rect 8392 5584 8444 5636
rect 10324 5720 10376 5772
rect 12072 5720 12124 5772
rect 12348 5720 12400 5772
rect 13084 5763 13136 5772
rect 13084 5729 13093 5763
rect 13093 5729 13127 5763
rect 13127 5729 13136 5763
rect 13084 5720 13136 5729
rect 13820 5720 13872 5772
rect 13912 5720 13964 5772
rect 18604 5788 18656 5840
rect 16028 5763 16080 5772
rect 16028 5729 16037 5763
rect 16037 5729 16071 5763
rect 16071 5729 16080 5763
rect 16028 5720 16080 5729
rect 16488 5763 16540 5772
rect 16488 5729 16497 5763
rect 16497 5729 16531 5763
rect 16531 5729 16540 5763
rect 16488 5720 16540 5729
rect 17224 5720 17276 5772
rect 23388 5720 23440 5772
rect 16304 5652 16356 5704
rect 17960 5652 18012 5704
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 18420 5652 18472 5661
rect 19340 5652 19392 5704
rect 19524 5652 19576 5704
rect 19984 5652 20036 5704
rect 20168 5652 20220 5704
rect 20628 5652 20680 5704
rect 24768 5695 24820 5704
rect 10692 5584 10744 5636
rect 10784 5627 10836 5636
rect 10784 5593 10793 5627
rect 10793 5593 10827 5627
rect 10827 5593 10836 5627
rect 10784 5584 10836 5593
rect 4068 5516 4120 5525
rect 4712 5516 4764 5568
rect 5540 5516 5592 5568
rect 8668 5516 8720 5568
rect 9588 5516 9640 5568
rect 9680 5516 9732 5568
rect 10508 5516 10560 5568
rect 11428 5516 11480 5568
rect 14556 5627 14608 5636
rect 13912 5516 13964 5568
rect 14556 5593 14565 5627
rect 14565 5593 14599 5627
rect 14599 5593 14608 5627
rect 14556 5584 14608 5593
rect 24768 5661 24777 5695
rect 24777 5661 24811 5695
rect 24811 5661 24820 5695
rect 24768 5652 24820 5661
rect 29644 5652 29696 5704
rect 22192 5584 22244 5636
rect 19432 5516 19484 5568
rect 19984 5516 20036 5568
rect 25688 5516 25740 5568
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3976 5312 4028 5364
rect 7012 5312 7064 5364
rect 1492 5176 1544 5228
rect 3792 5176 3844 5228
rect 2688 5151 2740 5160
rect 1584 5040 1636 5092
rect 2688 5117 2697 5151
rect 2697 5117 2731 5151
rect 2731 5117 2740 5151
rect 2688 5108 2740 5117
rect 6920 5244 6972 5296
rect 8208 5244 8260 5296
rect 9036 5244 9088 5296
rect 4620 5176 4672 5228
rect 10324 5312 10376 5364
rect 11704 5312 11756 5364
rect 11980 5287 12032 5296
rect 11980 5253 11989 5287
rect 11989 5253 12023 5287
rect 12023 5253 12032 5287
rect 11980 5244 12032 5253
rect 12256 5244 12308 5296
rect 13452 5244 13504 5296
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 13636 5244 13688 5296
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7472 5108 7524 5160
rect 13544 5108 13596 5160
rect 4068 4972 4120 5024
rect 4988 4972 5040 5024
rect 6000 4972 6052 5024
rect 6552 4972 6604 5024
rect 11612 5040 11664 5092
rect 15200 5312 15252 5364
rect 17040 5312 17092 5364
rect 17316 5312 17368 5364
rect 17868 5244 17920 5296
rect 19524 5287 19576 5296
rect 19524 5253 19533 5287
rect 19533 5253 19567 5287
rect 19567 5253 19576 5287
rect 19524 5244 19576 5253
rect 20076 5312 20128 5364
rect 21180 5312 21232 5364
rect 23388 5244 23440 5296
rect 15476 5176 15528 5228
rect 15660 5176 15712 5228
rect 16120 5176 16172 5228
rect 16580 5176 16632 5228
rect 18144 5219 18196 5228
rect 18144 5185 18153 5219
rect 18153 5185 18187 5219
rect 18187 5185 18196 5219
rect 18144 5176 18196 5185
rect 19064 5176 19116 5228
rect 19616 5176 19668 5228
rect 20076 5219 20128 5228
rect 14096 5151 14148 5160
rect 14096 5117 14105 5151
rect 14105 5117 14139 5151
rect 14139 5117 14148 5151
rect 14096 5108 14148 5117
rect 10508 4972 10560 5024
rect 11060 4972 11112 5024
rect 13820 5040 13872 5092
rect 18052 5108 18104 5160
rect 19340 5108 19392 5160
rect 20076 5185 20085 5219
rect 20085 5185 20119 5219
rect 20119 5185 20128 5219
rect 20076 5176 20128 5185
rect 20720 5219 20772 5228
rect 20720 5185 20729 5219
rect 20729 5185 20763 5219
rect 20763 5185 20772 5219
rect 20720 5176 20772 5185
rect 22652 5219 22704 5228
rect 22652 5185 22661 5219
rect 22661 5185 22695 5219
rect 22695 5185 22704 5219
rect 22652 5176 22704 5185
rect 31116 5219 31168 5228
rect 31116 5185 31125 5219
rect 31125 5185 31159 5219
rect 31159 5185 31168 5219
rect 31116 5176 31168 5185
rect 31208 5219 31260 5228
rect 31208 5185 31217 5219
rect 31217 5185 31251 5219
rect 31251 5185 31260 5219
rect 31208 5176 31260 5185
rect 30012 5108 30064 5160
rect 14464 5040 14516 5092
rect 14740 5040 14792 5092
rect 22100 5083 22152 5092
rect 22100 5049 22109 5083
rect 22109 5049 22143 5083
rect 22143 5049 22152 5083
rect 22100 5040 22152 5049
rect 31116 5040 31168 5092
rect 34428 5040 34480 5092
rect 13636 4972 13688 5024
rect 15476 4972 15528 5024
rect 15936 4972 15988 5024
rect 20628 4972 20680 5024
rect 22376 4972 22428 5024
rect 35808 4972 35860 5024
rect 38016 4972 38068 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 6552 4768 6604 4820
rect 8392 4768 8444 4820
rect 9404 4768 9456 4820
rect 15936 4768 15988 4820
rect 16120 4811 16172 4820
rect 16120 4777 16129 4811
rect 16129 4777 16163 4811
rect 16163 4777 16172 4811
rect 16120 4768 16172 4777
rect 17500 4811 17552 4820
rect 17500 4777 17509 4811
rect 17509 4777 17543 4811
rect 17543 4777 17552 4811
rect 17500 4768 17552 4777
rect 20352 4768 20404 4820
rect 21088 4768 21140 4820
rect 21548 4768 21600 4820
rect 2320 4632 2372 4684
rect 2688 4632 2740 4684
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 8944 4632 8996 4684
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 2964 4564 3016 4616
rect 4068 4564 4120 4616
rect 7748 4564 7800 4616
rect 8300 4564 8352 4616
rect 3148 4539 3200 4548
rect 3148 4505 3157 4539
rect 3157 4505 3191 4539
rect 3191 4505 3200 4539
rect 3148 4496 3200 4505
rect 6460 4496 6512 4548
rect 7104 4496 7156 4548
rect 9036 4564 9088 4616
rect 9404 4632 9456 4684
rect 10140 4632 10192 4684
rect 10324 4632 10376 4684
rect 12348 4700 12400 4752
rect 12992 4632 13044 4684
rect 9312 4564 9364 4616
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 12256 4564 12308 4616
rect 13820 4700 13872 4752
rect 15384 4700 15436 4752
rect 21916 4700 21968 4752
rect 13912 4632 13964 4684
rect 6368 4428 6420 4480
rect 9036 4428 9088 4480
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 10968 4496 11020 4548
rect 12716 4496 12768 4548
rect 15016 4607 15068 4616
rect 15016 4573 15025 4607
rect 15025 4573 15059 4607
rect 15059 4573 15068 4607
rect 15016 4564 15068 4573
rect 16212 4564 16264 4616
rect 18144 4632 18196 4684
rect 20444 4632 20496 4684
rect 16764 4607 16816 4616
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 16948 4564 17000 4616
rect 17960 4564 18012 4616
rect 18420 4564 18472 4616
rect 18788 4607 18840 4616
rect 18788 4573 18797 4607
rect 18797 4573 18831 4607
rect 18831 4573 18840 4607
rect 18788 4564 18840 4573
rect 13636 4428 13688 4480
rect 14740 4496 14792 4548
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 19064 4496 19116 4548
rect 15476 4428 15528 4480
rect 19432 4428 19484 4480
rect 19616 4428 19668 4480
rect 20076 4428 20128 4480
rect 22192 4564 22244 4616
rect 23112 4564 23164 4616
rect 22100 4539 22152 4548
rect 22100 4505 22109 4539
rect 22109 4505 22143 4539
rect 22143 4505 22152 4539
rect 22100 4496 22152 4505
rect 22008 4428 22060 4480
rect 22744 4471 22796 4480
rect 22744 4437 22753 4471
rect 22753 4437 22787 4471
rect 22787 4437 22796 4471
rect 22744 4428 22796 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 3148 4224 3200 4276
rect 5172 4156 5224 4208
rect 6368 4224 6420 4276
rect 8024 4224 8076 4276
rect 11980 4224 12032 4276
rect 12072 4224 12124 4276
rect 13452 4224 13504 4276
rect 7656 4156 7708 4208
rect 9588 4156 9640 4208
rect 9772 4156 9824 4208
rect 12256 4156 12308 4208
rect 22744 4224 22796 4276
rect 13636 4156 13688 4208
rect 17132 4156 17184 4208
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2964 4131 3016 4140
rect 2964 4097 2973 4131
rect 2973 4097 3007 4131
rect 3007 4097 3016 4131
rect 2964 4088 3016 4097
rect 5724 4088 5776 4140
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 9312 4088 9364 4140
rect 11060 4131 11112 4140
rect 11060 4097 11069 4131
rect 11069 4097 11103 4131
rect 11103 4097 11112 4131
rect 11704 4131 11756 4140
rect 11060 4088 11112 4097
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 17684 4088 17736 4140
rect 3240 4063 3292 4072
rect 3240 4029 3249 4063
rect 3249 4029 3283 4063
rect 3283 4029 3292 4063
rect 3240 4020 3292 4029
rect 4068 4020 4120 4072
rect 6000 4020 6052 4072
rect 7472 4020 7524 4072
rect 9680 4020 9732 4072
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 9956 4020 10008 4072
rect 11428 4020 11480 4072
rect 11980 4063 12032 4072
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 13728 4020 13780 4072
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 7288 3952 7340 4004
rect 10232 3952 10284 4004
rect 17592 4020 17644 4072
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 18420 4088 18472 4097
rect 17868 4020 17920 4072
rect 19432 4156 19484 4208
rect 19064 4131 19116 4140
rect 19064 4097 19073 4131
rect 19073 4097 19107 4131
rect 19107 4097 19116 4131
rect 19064 4088 19116 4097
rect 19340 4020 19392 4072
rect 20720 4088 20772 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22652 4131 22704 4140
rect 22008 4088 22060 4097
rect 22652 4097 22661 4131
rect 22661 4097 22695 4131
rect 22695 4097 22704 4131
rect 22652 4088 22704 4097
rect 26700 4088 26752 4140
rect 19800 4020 19852 4072
rect 26608 4020 26660 4072
rect 4620 3884 4672 3936
rect 5448 3884 5500 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 10416 3884 10468 3936
rect 11060 3884 11112 3936
rect 12440 3884 12492 3936
rect 12532 3884 12584 3936
rect 14372 3884 14424 3936
rect 14464 3884 14516 3936
rect 16856 3952 16908 4004
rect 19432 3952 19484 4004
rect 20812 3952 20864 4004
rect 15660 3884 15712 3936
rect 19156 3927 19208 3936
rect 19156 3893 19165 3927
rect 19165 3893 19199 3927
rect 19199 3893 19208 3927
rect 19156 3884 19208 3893
rect 19248 3884 19300 3936
rect 20536 3884 20588 3936
rect 20904 3884 20956 3936
rect 22284 3884 22336 3936
rect 28908 3884 28960 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 10232 3680 10284 3732
rect 10324 3680 10376 3732
rect 3240 3612 3292 3664
rect 13728 3655 13780 3664
rect 5632 3544 5684 3596
rect 6000 3587 6052 3596
rect 6000 3553 6009 3587
rect 6009 3553 6043 3587
rect 6043 3553 6052 3587
rect 6000 3544 6052 3553
rect 9772 3544 9824 3596
rect 2596 3519 2648 3528
rect 2596 3485 2605 3519
rect 2605 3485 2639 3519
rect 2639 3485 2648 3519
rect 2596 3476 2648 3485
rect 2964 3476 3016 3528
rect 5724 3476 5776 3528
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 9312 3476 9364 3528
rect 11520 3587 11572 3596
rect 11520 3553 11529 3587
rect 11529 3553 11563 3587
rect 11563 3553 11572 3587
rect 11520 3544 11572 3553
rect 11704 3544 11756 3596
rect 13728 3621 13737 3655
rect 13737 3621 13771 3655
rect 13771 3621 13780 3655
rect 13728 3612 13780 3621
rect 16028 3655 16080 3664
rect 16028 3621 16037 3655
rect 16037 3621 16071 3655
rect 16071 3621 16080 3655
rect 16028 3612 16080 3621
rect 13452 3544 13504 3596
rect 5080 3408 5132 3460
rect 1860 3340 1912 3392
rect 3516 3340 3568 3392
rect 5816 3408 5868 3460
rect 7840 3408 7892 3460
rect 9772 3451 9824 3460
rect 9772 3417 9781 3451
rect 9781 3417 9815 3451
rect 9815 3417 9824 3451
rect 9772 3408 9824 3417
rect 11428 3408 11480 3460
rect 12164 3408 12216 3460
rect 12256 3451 12308 3460
rect 12256 3417 12265 3451
rect 12265 3417 12299 3451
rect 12299 3417 12308 3451
rect 12256 3408 12308 3417
rect 13544 3408 13596 3460
rect 10416 3340 10468 3392
rect 10692 3340 10744 3392
rect 14004 3476 14056 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 17408 3680 17460 3732
rect 19248 3680 19300 3732
rect 19524 3723 19576 3732
rect 19524 3689 19533 3723
rect 19533 3689 19567 3723
rect 19567 3689 19576 3723
rect 19524 3680 19576 3689
rect 21456 3723 21508 3732
rect 21456 3689 21465 3723
rect 21465 3689 21499 3723
rect 21499 3689 21508 3723
rect 21456 3680 21508 3689
rect 22468 3723 22520 3732
rect 22468 3689 22477 3723
rect 22477 3689 22511 3723
rect 22511 3689 22520 3723
rect 22468 3680 22520 3689
rect 23204 3680 23256 3732
rect 26700 3723 26752 3732
rect 26700 3689 26709 3723
rect 26709 3689 26743 3723
rect 26743 3689 26752 3723
rect 26700 3680 26752 3689
rect 31392 3680 31444 3732
rect 16856 3612 16908 3664
rect 19800 3612 19852 3664
rect 18236 3544 18288 3596
rect 16856 3476 16908 3528
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 18420 3476 18472 3528
rect 13728 3408 13780 3460
rect 14464 3408 14516 3460
rect 14832 3408 14884 3460
rect 19340 3476 19392 3528
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 22100 3587 22152 3596
rect 22100 3553 22109 3587
rect 22109 3553 22143 3587
rect 22143 3553 22152 3587
rect 22100 3544 22152 3553
rect 23480 3519 23532 3528
rect 23480 3485 23489 3519
rect 23489 3485 23523 3519
rect 23523 3485 23532 3519
rect 23480 3476 23532 3485
rect 26608 3519 26660 3528
rect 26608 3485 26617 3519
rect 26617 3485 26651 3519
rect 26651 3485 26660 3519
rect 26608 3476 26660 3485
rect 38292 3519 38344 3528
rect 38292 3485 38301 3519
rect 38301 3485 38335 3519
rect 38335 3485 38344 3519
rect 38292 3476 38344 3485
rect 17960 3383 18012 3392
rect 17960 3349 17969 3383
rect 17969 3349 18003 3383
rect 18003 3349 18012 3383
rect 17960 3340 18012 3349
rect 20076 3340 20128 3392
rect 20352 3340 20404 3392
rect 22836 3383 22888 3392
rect 22836 3349 22845 3383
rect 22845 3349 22879 3383
rect 22879 3349 22888 3383
rect 22836 3340 22888 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 7104 3136 7156 3188
rect 3884 3068 3936 3120
rect 8116 3068 8168 3120
rect 12164 3136 12216 3188
rect 12348 3136 12400 3188
rect 12992 3136 13044 3188
rect 13360 3136 13412 3188
rect 13636 3136 13688 3188
rect 18328 3136 18380 3188
rect 23940 3179 23992 3188
rect 23940 3145 23949 3179
rect 23949 3145 23983 3179
rect 23983 3145 23992 3179
rect 23940 3136 23992 3145
rect 35716 3136 35768 3188
rect 10232 3068 10284 3120
rect 4068 3000 4120 3052
rect 1308 2932 1360 2984
rect 3424 2932 3476 2984
rect 3516 2932 3568 2984
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 7472 3000 7524 3052
rect 10140 3000 10192 3052
rect 10692 3068 10744 3120
rect 11520 3068 11572 3120
rect 13268 3068 13320 3120
rect 14372 3068 14424 3120
rect 17960 3068 18012 3120
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 13084 3000 13136 3052
rect 16672 3000 16724 3052
rect 9956 2975 10008 2984
rect 4160 2864 4212 2916
rect 9956 2941 9965 2975
rect 9965 2941 9999 2975
rect 9999 2941 10008 2975
rect 9956 2932 10008 2941
rect 10508 2932 10560 2984
rect 13728 2932 13780 2984
rect 14004 2975 14056 2984
rect 14004 2941 14036 2975
rect 14036 2941 14056 2975
rect 14004 2932 14056 2941
rect 14372 2932 14424 2984
rect 17868 3000 17920 3052
rect 19340 3000 19392 3052
rect 23112 3043 23164 3052
rect 23112 3009 23121 3043
rect 23121 3009 23155 3043
rect 23155 3009 23164 3043
rect 23112 3000 23164 3009
rect 23572 3000 23624 3052
rect 37280 3000 37332 3052
rect 38016 3043 38068 3052
rect 38016 3009 38025 3043
rect 38025 3009 38059 3043
rect 38059 3009 38068 3043
rect 38016 3000 38068 3009
rect 11612 2864 11664 2916
rect 15752 2907 15804 2916
rect 15752 2873 15761 2907
rect 15761 2873 15795 2907
rect 15795 2873 15804 2907
rect 15752 2864 15804 2873
rect 15844 2864 15896 2916
rect 18604 2864 18656 2916
rect 22192 2864 22244 2916
rect 7656 2796 7708 2848
rect 10140 2796 10192 2848
rect 13636 2796 13688 2848
rect 13820 2796 13872 2848
rect 18880 2839 18932 2848
rect 18880 2805 18889 2839
rect 18889 2805 18923 2839
rect 18923 2805 18932 2839
rect 18880 2796 18932 2805
rect 18972 2796 19024 2848
rect 20168 2839 20220 2848
rect 20168 2805 20177 2839
rect 20177 2805 20211 2839
rect 20211 2805 20220 2839
rect 20168 2796 20220 2805
rect 20720 2796 20772 2848
rect 22100 2839 22152 2848
rect 22100 2805 22109 2839
rect 22109 2805 22143 2839
rect 22143 2805 22152 2839
rect 38200 2839 38252 2848
rect 22100 2796 22152 2805
rect 38200 2805 38209 2839
rect 38209 2805 38243 2839
rect 38243 2805 38252 2839
rect 38200 2796 38252 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 4988 2592 5040 2644
rect 9772 2592 9824 2644
rect 4068 2524 4120 2576
rect 5908 2524 5960 2576
rect 11152 2592 11204 2644
rect 1308 2388 1360 2440
rect 6000 2456 6052 2508
rect 7472 2456 7524 2508
rect 9312 2499 9364 2508
rect 9312 2465 9321 2499
rect 9321 2465 9355 2499
rect 9355 2465 9364 2499
rect 9312 2456 9364 2465
rect 11704 2499 11756 2508
rect 11704 2465 11713 2499
rect 11713 2465 11747 2499
rect 11747 2465 11756 2499
rect 14280 2499 14332 2508
rect 11704 2456 11756 2465
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 14648 2592 14700 2644
rect 16764 2592 16816 2644
rect 19340 2592 19392 2644
rect 20168 2592 20220 2644
rect 20260 2592 20312 2644
rect 24216 2592 24268 2644
rect 28448 2592 28500 2644
rect 30196 2592 30248 2644
rect 34704 2592 34756 2644
rect 17224 2524 17276 2576
rect 22836 2524 22888 2576
rect 24584 2567 24636 2576
rect 24584 2533 24593 2567
rect 24593 2533 24627 2567
rect 24627 2533 24636 2567
rect 24584 2524 24636 2533
rect 34428 2524 34480 2576
rect 35624 2524 35676 2576
rect 15568 2456 15620 2508
rect 18972 2456 19024 2508
rect 19432 2456 19484 2508
rect 22744 2499 22796 2508
rect 16764 2388 16816 2440
rect 18604 2431 18656 2440
rect 1952 2363 2004 2372
rect 1952 2329 1961 2363
rect 1961 2329 1995 2363
rect 1995 2329 2004 2363
rect 1952 2320 2004 2329
rect 4436 2363 4488 2372
rect 4436 2329 4445 2363
rect 4445 2329 4479 2363
rect 4479 2329 4488 2363
rect 4436 2320 4488 2329
rect 6828 2320 6880 2372
rect 8484 2320 8536 2372
rect 8576 2363 8628 2372
rect 8576 2329 8585 2363
rect 8585 2329 8619 2363
rect 8619 2329 8628 2363
rect 9588 2363 9640 2372
rect 8576 2320 8628 2329
rect 9588 2329 9597 2363
rect 9597 2329 9631 2363
rect 9631 2329 9640 2363
rect 9588 2320 9640 2329
rect 10048 2320 10100 2372
rect 10876 2320 10928 2372
rect 14464 2320 14516 2372
rect 14556 2363 14608 2372
rect 14556 2329 14565 2363
rect 14565 2329 14599 2363
rect 14599 2329 14608 2363
rect 14556 2320 14608 2329
rect 16120 2320 16172 2372
rect 18604 2397 18613 2431
rect 18613 2397 18647 2431
rect 18647 2397 18656 2431
rect 18604 2388 18656 2397
rect 18788 2388 18840 2440
rect 22744 2465 22753 2499
rect 22753 2465 22787 2499
rect 22787 2465 22796 2499
rect 22744 2456 22796 2465
rect 25688 2456 25740 2508
rect 5448 2252 5500 2304
rect 6920 2252 6972 2304
rect 10968 2252 11020 2304
rect 21272 2388 21324 2440
rect 23112 2388 23164 2440
rect 21916 2320 21968 2372
rect 24492 2388 24544 2440
rect 26424 2388 26476 2440
rect 28908 2456 28960 2508
rect 29000 2388 29052 2440
rect 35808 2456 35860 2508
rect 32220 2388 32272 2440
rect 34152 2388 34204 2440
rect 35440 2388 35492 2440
rect 33876 2320 33928 2372
rect 35624 2320 35676 2372
rect 38660 2320 38712 2372
rect 15292 2252 15344 2304
rect 15568 2252 15620 2304
rect 18512 2252 18564 2304
rect 18696 2252 18748 2304
rect 19432 2295 19484 2304
rect 19432 2261 19441 2295
rect 19441 2261 19475 2295
rect 19475 2261 19484 2295
rect 19432 2252 19484 2261
rect 19984 2252 20036 2304
rect 20444 2295 20496 2304
rect 20444 2261 20453 2295
rect 20453 2261 20487 2295
rect 20487 2261 20496 2295
rect 20444 2252 20496 2261
rect 20812 2295 20864 2304
rect 20812 2261 20821 2295
rect 20821 2261 20855 2295
rect 20855 2261 20864 2295
rect 20812 2252 20864 2261
rect 23204 2252 23256 2304
rect 27712 2252 27764 2304
rect 30932 2252 30984 2304
rect 37372 2252 37424 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 4436 2048 4488 2100
rect 9956 2048 10008 2100
rect 14464 2048 14516 2100
rect 17224 2048 17276 2100
rect 8484 1980 8536 2032
rect 13268 1980 13320 2032
rect 13452 1980 13504 2032
rect 20352 1980 20404 2032
rect 5816 1912 5868 1964
rect 20444 1912 20496 1964
rect 11612 1844 11664 1896
rect 20812 1844 20864 1896
rect 8300 1776 8352 1828
rect 19340 1776 19392 1828
rect 12256 1708 12308 1760
rect 18788 1708 18840 1760
rect 9588 1640 9640 1692
rect 15660 1640 15712 1692
rect 5540 1572 5592 1624
rect 13268 1572 13320 1624
rect 20720 1572 20772 1624
rect 20536 1436 20588 1488
rect 8576 1368 8628 1420
rect 14556 1368 14608 1420
rect 15476 1368 15528 1420
rect 16120 1368 16172 1420
rect 20 1300 72 1352
rect 4712 1300 4764 1352
rect 3792 1232 3844 1284
rect 20076 1300 20128 1352
rect 3976 1096 4028 1148
rect 18880 1232 18932 1284
rect 4988 1164 5040 1216
rect 20628 1164 20680 1216
rect 7564 1096 7616 1148
rect 22376 1096 22428 1148
rect 5264 1028 5316 1080
rect 19156 1028 19208 1080
rect 6644 960 6696 1012
rect 20260 960 20312 1012
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 2778 39536 2834 39545
rect 2778 39471 2834 39480
rect 676 36922 704 39200
rect 1964 37262 1992 39200
rect 1860 37256 1912 37262
rect 1860 37198 1912 37204
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 1872 36922 1900 37198
rect 2792 37194 2820 39471
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 16224 39222 16528 39250
rect 3146 37496 3202 37505
rect 3146 37431 3202 37440
rect 3160 37262 3188 37431
rect 3148 37256 3200 37262
rect 3148 37198 3200 37204
rect 2780 37188 2832 37194
rect 2780 37130 2832 37136
rect 3896 37126 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 2872 37120 2924 37126
rect 2872 37062 2924 37068
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 2884 36922 2912 37062
rect 664 36916 716 36922
rect 664 36858 716 36864
rect 1860 36916 1912 36922
rect 1860 36858 1912 36864
rect 2872 36916 2924 36922
rect 2872 36858 2924 36864
rect 2504 36780 2556 36786
rect 2504 36722 2556 36728
rect 1768 36168 1820 36174
rect 1766 36136 1768 36145
rect 1820 36136 1822 36145
rect 1766 36071 1822 36080
rect 2516 35834 2544 36722
rect 2688 36032 2740 36038
rect 2688 35974 2740 35980
rect 2504 35828 2556 35834
rect 2504 35770 2556 35776
rect 2412 35692 2464 35698
rect 2412 35634 2464 35640
rect 1768 34400 1820 34406
rect 1768 34342 1820 34348
rect 1780 34105 1808 34342
rect 1766 34096 1822 34105
rect 1766 34031 1822 34040
rect 1768 32904 1820 32910
rect 1768 32846 1820 32852
rect 1780 32745 1808 32846
rect 1766 32736 1822 32745
rect 1766 32671 1822 32680
rect 1768 30728 1820 30734
rect 1766 30696 1768 30705
rect 1820 30696 1822 30705
rect 1766 30631 1822 30640
rect 1768 29504 1820 29510
rect 1768 29446 1820 29452
rect 1780 29345 1808 29446
rect 1766 29336 1822 29345
rect 1766 29271 1822 29280
rect 1768 28076 1820 28082
rect 1768 28018 1820 28024
rect 1780 27985 1808 28018
rect 1766 27976 1822 27985
rect 1766 27911 1822 27920
rect 1768 26376 1820 26382
rect 1768 26318 1820 26324
rect 1780 25945 1808 26318
rect 1766 25936 1822 25945
rect 1766 25871 1822 25880
rect 1768 24608 1820 24614
rect 1766 24576 1768 24585
rect 1820 24576 1822 24585
rect 1766 24511 1822 24520
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1780 22545 1808 22578
rect 1766 22536 1822 22545
rect 1766 22471 1822 22480
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1780 21185 1808 21286
rect 1766 21176 1822 21185
rect 1766 21111 1822 21120
rect 2424 20369 2452 35634
rect 2700 29646 2728 35974
rect 3792 30592 3844 30598
rect 3792 30534 3844 30540
rect 2688 29640 2740 29646
rect 2688 29582 2740 29588
rect 2780 29572 2832 29578
rect 2780 29514 2832 29520
rect 2792 29034 2820 29514
rect 2780 29028 2832 29034
rect 2780 28970 2832 28976
rect 3804 27470 3832 30534
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 3896 23730 3924 27814
rect 3884 23724 3936 23730
rect 3884 23666 3936 23672
rect 2410 20360 2466 20369
rect 2410 20295 2466 20304
rect 1768 19848 1820 19854
rect 1766 19816 1768 19825
rect 1820 19816 1822 19825
rect 1766 19751 1822 19760
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 5234 1532 15846
rect 1596 15026 1624 18022
rect 1780 17785 1808 18226
rect 3988 18086 4016 37198
rect 5184 37126 5212 39200
rect 7116 37330 7144 39200
rect 7104 37324 7156 37330
rect 7104 37266 7156 37272
rect 8404 37262 8432 39200
rect 10336 37262 10364 39200
rect 11624 37262 11652 39200
rect 12912 37262 12940 39200
rect 6736 37256 6788 37262
rect 6736 37198 6788 37204
rect 7472 37256 7524 37262
rect 7472 37198 7524 37204
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 10324 37256 10376 37262
rect 10324 37198 10376 37204
rect 11612 37256 11664 37262
rect 11612 37198 11664 37204
rect 12900 37256 12952 37262
rect 12900 37198 12952 37204
rect 6552 37188 6604 37194
rect 6552 37130 6604 37136
rect 5172 37120 5224 37126
rect 5172 37062 5224 37068
rect 5448 36916 5500 36922
rect 5448 36858 5500 36864
rect 4068 36712 4120 36718
rect 4068 36654 4120 36660
rect 4080 35290 4108 36654
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 35284 4120 35290
rect 4068 35226 4120 35232
rect 4068 34604 4120 34610
rect 4068 34546 4120 34552
rect 4080 30938 4108 34546
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 5460 31822 5488 36858
rect 5540 32768 5592 32774
rect 5540 32710 5592 32716
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4068 30932 4120 30938
rect 4068 30874 4120 30880
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 4080 29073 4108 29446
rect 4066 29064 4122 29073
rect 4066 28999 4122 29008
rect 4068 28960 4120 28966
rect 4068 28902 4120 28908
rect 4080 26042 4108 28902
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5552 28558 5580 32710
rect 6564 32434 6592 37130
rect 6748 34746 6776 37198
rect 7484 36553 7512 37198
rect 11980 37188 12032 37194
rect 11980 37130 12032 37136
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 10784 37120 10836 37126
rect 10784 37062 10836 37068
rect 7470 36544 7526 36553
rect 7470 36479 7526 36488
rect 7196 35080 7248 35086
rect 7196 35022 7248 35028
rect 6736 34740 6788 34746
rect 6736 34682 6788 34688
rect 7208 34202 7236 35022
rect 7196 34196 7248 34202
rect 7196 34138 7248 34144
rect 7104 33992 7156 33998
rect 7104 33934 7156 33940
rect 7116 32434 7144 33934
rect 6552 32428 6604 32434
rect 6552 32370 6604 32376
rect 7104 32428 7156 32434
rect 7104 32370 7156 32376
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6092 30728 6144 30734
rect 6092 30670 6144 30676
rect 6104 29850 6132 30670
rect 6092 29844 6144 29850
rect 6092 29786 6144 29792
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5080 26512 5132 26518
rect 5080 26454 5132 26460
rect 4068 26036 4120 26042
rect 4068 25978 4120 25984
rect 4620 25900 4672 25906
rect 4620 25842 4672 25848
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22098 4660 25842
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 1766 17776 1822 17785
rect 1766 17711 1822 17720
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1688 14074 1716 16526
rect 1768 16448 1820 16454
rect 1766 16416 1768 16425
rect 1820 16416 1822 16425
rect 1766 16351 1822 16360
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 14385 1808 15438
rect 1766 14376 1822 14385
rect 1766 14311 1822 14320
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 13394 1624 13806
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1596 12850 1624 13330
rect 1780 13025 1808 14214
rect 1766 13016 1822 13025
rect 1766 12951 1822 12960
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 12322 1624 12786
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12434 1716 12582
rect 1688 12406 1808 12434
rect 1596 12294 1716 12322
rect 1688 12238 1716 12294
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1688 11694 1716 12174
rect 1676 11688 1728 11694
rect 1596 11648 1676 11676
rect 1596 11150 1624 11648
rect 1676 11630 1728 11636
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10538 1624 11086
rect 1780 10810 1808 12406
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1584 10532 1636 10538
rect 1584 10474 1636 10480
rect 1596 10062 1624 10474
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9518 1624 9998
rect 1872 9674 1900 17478
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2148 16574 2176 16934
rect 2148 16546 2268 16574
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 13870 1992 14758
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 1964 12753 1992 13194
rect 1950 12744 2006 12753
rect 1950 12679 2006 12688
rect 2056 11830 2084 16050
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2148 14006 2176 14962
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 2044 11824 2096 11830
rect 2044 11766 2096 11772
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1780 9646 1900 9674
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 8974 1624 9454
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8430 1624 8910
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 7886 1624 8366
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7342 1624 7822
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 6798 1624 7278
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 6254 1624 6734
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1596 5710 1624 6190
rect 1780 5817 1808 9646
rect 1860 9512 1912 9518
rect 1858 9480 1860 9489
rect 1912 9480 1914 9489
rect 1858 9415 1914 9424
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1872 8906 1900 9318
rect 1964 9178 1992 11698
rect 2148 10674 2176 13942
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1872 7478 1900 8026
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 2240 6730 2268 16546
rect 2332 14618 2360 17614
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2424 16590 2452 17138
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2424 16114 2452 16526
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2332 6662 2360 10610
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2424 6118 2452 16050
rect 2516 6458 2544 17478
rect 2608 15502 2636 17478
rect 2792 17202 2820 17614
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2700 16833 2728 16934
rect 2686 16824 2742 16833
rect 2686 16759 2742 16768
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2596 15496 2648 15502
rect 2700 15473 2728 15846
rect 2596 15438 2648 15444
rect 2686 15464 2742 15473
rect 2686 15399 2742 15408
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2700 14550 2728 15302
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2792 12288 2820 16458
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2884 14006 2912 16390
rect 2976 16182 3004 16526
rect 2964 16176 3016 16182
rect 2964 16118 3016 16124
rect 3068 15994 3096 18022
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 2976 15966 3096 15994
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2976 12434 3004 15966
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 3068 14482 3096 15302
rect 3160 15178 3188 17138
rect 3252 15337 3280 17614
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4724 17270 4752 17478
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 4816 17134 4844 21966
rect 5092 21554 5120 26454
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5460 22778 5488 24754
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5552 22094 5580 22374
rect 5552 22066 5672 22094
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 4908 20602 4936 21490
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 4896 20596 4948 20602
rect 4896 20538 4948 20544
rect 5552 20466 5580 21286
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4620 17128 4672 17134
rect 3330 17096 3386 17105
rect 4620 17070 4672 17076
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 3330 17031 3332 17040
rect 3384 17031 3386 17040
rect 3332 17002 3384 17008
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16658 4660 17070
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3238 15328 3294 15337
rect 3238 15263 3294 15272
rect 3160 15150 3280 15178
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3160 13734 3188 14962
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 2700 12260 2820 12288
rect 2884 12406 3004 12434
rect 2700 11665 2728 12260
rect 2778 12200 2834 12209
rect 2778 12135 2834 12144
rect 2686 11656 2742 11665
rect 2686 11591 2742 11600
rect 2686 11112 2742 11121
rect 2686 11047 2742 11056
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2608 8090 2636 9862
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2700 6458 2728 11047
rect 2792 11014 2820 12135
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2792 6254 2820 10678
rect 2884 8430 2912 12406
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 3054 12064 3110 12073
rect 2976 11898 3004 12038
rect 3054 11999 3110 12008
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3068 11694 3096 11999
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3068 9874 3096 11630
rect 3160 10742 3188 13670
rect 3252 12209 3280 15150
rect 3344 12918 3372 16390
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 3976 16040 4028 16046
rect 4448 16017 4476 16050
rect 3976 15982 4028 15988
rect 4434 16008 4490 16017
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3436 14414 3464 14758
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3238 12200 3294 12209
rect 3238 12135 3294 12144
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 3148 10600 3200 10606
rect 3252 10588 3280 12038
rect 3436 11778 3464 12718
rect 3528 12102 3556 15846
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3620 11880 3648 15438
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3712 12714 3740 13194
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3804 12238 3832 14758
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3896 12850 3924 12922
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3620 11852 3740 11880
rect 3436 11750 3648 11778
rect 3620 11694 3648 11750
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11286 3648 11494
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3606 11112 3662 11121
rect 3606 11047 3608 11056
rect 3660 11047 3662 11056
rect 3608 11018 3660 11024
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3606 10976 3662 10985
rect 3200 10560 3280 10588
rect 3148 10542 3200 10548
rect 2976 9846 3096 9874
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5896 2452 6054
rect 2332 5868 2452 5896
rect 1766 5808 1822 5817
rect 1766 5743 1822 5752
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1596 5098 1624 5646
rect 1584 5092 1636 5098
rect 1584 5034 1636 5040
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4865 1808 4966
rect 1766 4856 1822 4865
rect 1766 4791 1822 4800
rect 2332 4690 2360 5868
rect 2976 5846 3004 9846
rect 3054 9752 3110 9761
rect 3054 9687 3110 9696
rect 3068 6225 3096 9687
rect 3160 8838 3188 10542
rect 3344 10418 3372 10950
rect 3606 10911 3662 10920
rect 3252 10390 3372 10418
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3252 7018 3280 10390
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3332 9104 3384 9110
rect 3330 9072 3332 9081
rect 3384 9072 3386 9081
rect 3330 9007 3386 9016
rect 3330 8528 3386 8537
rect 3330 8463 3332 8472
rect 3384 8463 3386 8472
rect 3332 8434 3384 8440
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3160 6990 3280 7018
rect 3344 7002 3372 7686
rect 3332 6996 3384 7002
rect 3054 6216 3110 6225
rect 3054 6151 3110 6160
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2700 4690 2728 5102
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 1872 4146 1900 4558
rect 2976 4146 3004 4558
rect 3160 4554 3188 6990
rect 3332 6938 3384 6944
rect 3436 6361 3464 9590
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3422 6352 3478 6361
rect 3422 6287 3478 6296
rect 3528 6225 3556 8842
rect 3620 7954 3648 10911
rect 3712 8378 3740 11852
rect 3896 10010 3924 12650
rect 3988 10130 4016 15982
rect 4434 15943 4490 15952
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4816 15450 4844 17070
rect 5184 16250 5212 17614
rect 5552 16658 5580 19654
rect 5644 19378 5672 22066
rect 6276 21412 6328 21418
rect 6276 21354 6328 21360
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16250 5764 16390
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5264 16176 5316 16182
rect 5264 16118 5316 16124
rect 5172 15496 5224 15502
rect 4816 15422 4936 15450
rect 5172 15438 5224 15444
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4080 13938 4108 14214
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4540 13818 4568 14554
rect 4632 14482 4660 15302
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4540 13790 4660 13818
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4158 13288 4214 13297
rect 4632 13274 4660 13790
rect 4158 13223 4214 13232
rect 4540 13246 4660 13274
rect 4172 12918 4200 13223
rect 4436 13184 4488 13190
rect 4434 13152 4436 13161
rect 4488 13152 4490 13161
rect 4434 13087 4490 13096
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4540 12782 4568 13246
rect 4724 13172 4752 14758
rect 4632 13144 4752 13172
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4160 12232 4212 12238
rect 4066 12200 4122 12209
rect 4160 12174 4212 12180
rect 4066 12135 4068 12144
rect 4120 12135 4122 12144
rect 4068 12106 4120 12112
rect 4068 11824 4120 11830
rect 4066 11792 4068 11801
rect 4120 11792 4122 11801
rect 4066 11727 4122 11736
rect 4172 11540 4200 12174
rect 4250 11928 4306 11937
rect 4250 11863 4306 11872
rect 4264 11762 4292 11863
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4356 11626 4384 12310
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4080 11512 4200 11540
rect 4080 10130 4108 11512
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4448 10470 4476 11018
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4526 10160 4582 10169
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 4068 10124 4120 10130
rect 4526 10095 4582 10104
rect 4068 10066 4120 10072
rect 3896 9982 4016 10010
rect 3988 9674 4016 9982
rect 3988 9646 4108 9674
rect 3882 9616 3938 9625
rect 3882 9551 3938 9560
rect 3896 8634 3924 9551
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 9042 4016 9454
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3712 8350 3832 8378
rect 3700 8288 3752 8294
rect 3698 8256 3700 8265
rect 3752 8256 3754 8265
rect 3698 8191 3754 8200
rect 3804 8022 3832 8350
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3882 7984 3938 7993
rect 3608 7948 3660 7954
rect 4080 7970 4108 9646
rect 4540 9382 4568 10095
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4526 9072 4582 9081
rect 4526 9007 4582 9016
rect 4540 8276 4568 9007
rect 4632 8498 4660 13144
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4724 9058 4752 12718
rect 4816 12306 4844 15302
rect 4908 14482 4936 15422
rect 5184 15026 5212 15438
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4896 14340 4948 14346
rect 4896 14282 4948 14288
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4908 12170 4936 14282
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5000 12986 5028 13262
rect 5092 12986 5120 13670
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5000 12306 5028 12922
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4894 11656 4950 11665
rect 4816 10810 4844 11630
rect 4894 11591 4950 11600
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4816 9489 4844 10406
rect 4908 9654 4936 11591
rect 5000 11218 5028 12242
rect 5092 11898 5120 12922
rect 5184 12782 5212 14962
rect 5276 13025 5304 16118
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5368 15162 5396 15438
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5552 15026 5580 16050
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 14346 5396 14758
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5644 14226 5672 15846
rect 5828 15144 5856 20538
rect 6288 16658 6316 21354
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 5552 14198 5672 14226
rect 5736 15116 5856 15144
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5368 13394 5396 13874
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5460 13297 5488 13738
rect 5446 13288 5502 13297
rect 5446 13223 5502 13232
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5262 13016 5318 13025
rect 5262 12951 5318 12960
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5276 12617 5304 12786
rect 5368 12782 5396 13126
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5262 12608 5318 12617
rect 5262 12543 5318 12552
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 5446 12336 5502 12345
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5092 11558 5120 11698
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5184 11098 5212 12174
rect 5000 11070 5212 11098
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4802 9480 4858 9489
rect 4802 9415 4858 9424
rect 4724 9030 4936 9058
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4540 8248 4660 8276
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3882 7919 3938 7928
rect 3988 7942 4108 7970
rect 3608 7890 3660 7896
rect 3896 7886 3924 7919
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3896 6866 3924 7278
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3514 6216 3570 6225
rect 3514 6151 3570 6160
rect 3988 5370 4016 7942
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4080 6497 4108 7754
rect 4632 7342 4660 8248
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4618 7168 4674 7177
rect 4214 7100 4522 7109
rect 4618 7103 4674 7112
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 7002 4660 7103
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 4172 6390 4200 6598
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4172 6100 4200 6326
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4080 6072 4200 6100
rect 4080 5914 4108 6072
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4158 5808 4214 5817
rect 4158 5743 4214 5752
rect 4172 5710 4200 5743
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4080 5574 4108 5646
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4632 5234 4660 6190
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3160 4282 3188 4490
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 1872 3398 1900 4082
rect 2976 3534 3004 4082
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3252 3670 3280 4014
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 1320 2446 1348 2926
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 20 1352 72 1358
rect 20 1294 72 1300
rect 32 800 60 1294
rect 1320 800 1348 2382
rect 1952 2372 2004 2378
rect 1952 2314 2004 2320
rect 1964 2281 1992 2314
rect 1950 2272 2006 2281
rect 1950 2207 2006 2216
rect 2608 800 2636 3470
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 2990 3556 3334
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3436 2650 3464 2926
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3804 1290 3832 5170
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4622 4108 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4080 4078 4108 4558
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3896 2774 3924 3062
rect 4080 3058 4108 4014
rect 4632 3942 4660 5170
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4618 3632 4674 3641
rect 4618 3567 4674 3576
rect 4158 3360 4214 3369
rect 4158 3295 4214 3304
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3896 2746 4016 2774
rect 3792 1284 3844 1290
rect 3792 1226 3844 1232
rect 3988 1154 4016 2746
rect 4080 2582 4108 2994
rect 4172 2922 4200 3295
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 4448 2106 4476 2314
rect 4436 2100 4488 2106
rect 4436 2042 4488 2048
rect 3976 1148 4028 1154
rect 3976 1090 4028 1096
rect 4632 1034 4660 3567
rect 4724 1358 4752 5510
rect 4816 1986 4844 8842
rect 4908 2774 4936 9030
rect 5000 8566 5028 11070
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5092 10198 5120 10406
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5000 6866 5028 7822
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 5000 5710 5028 6802
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 5030 5028 5646
rect 4988 5024 5040 5030
rect 5092 5001 5120 9318
rect 5184 8090 5212 10610
rect 5276 9042 5304 12310
rect 5446 12271 5502 12280
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5368 10266 5396 11834
rect 5460 10826 5488 12271
rect 5552 11150 5580 14198
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5460 10798 5580 10826
rect 5448 10736 5500 10742
rect 5446 10704 5448 10713
rect 5500 10704 5502 10713
rect 5446 10639 5502 10648
rect 5552 10588 5580 10798
rect 5460 10560 5580 10588
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5368 7818 5396 10202
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 4988 4966 5040 4972
rect 5078 4992 5134 5001
rect 5078 4927 5134 4936
rect 5092 3466 5120 4927
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 4908 2746 5028 2774
rect 5000 2650 5028 2746
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4816 1958 5028 1986
rect 4712 1352 4764 1358
rect 4712 1294 4764 1300
rect 5000 1222 5028 1958
rect 5184 1329 5212 4150
rect 5170 1320 5226 1329
rect 5170 1255 5226 1264
rect 4988 1216 5040 1222
rect 4988 1158 5040 1164
rect 5276 1086 5304 6666
rect 5368 5273 5396 7346
rect 5460 7342 5488 10560
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5460 6254 5488 7278
rect 5552 6798 5580 9930
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5644 6186 5672 13126
rect 5736 13002 5764 15116
rect 6288 15094 6316 15302
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5828 13530 5856 14962
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5736 12974 5948 13002
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5736 12646 5764 12854
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11694 5764 12106
rect 5828 11898 5856 12378
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5724 11688 5776 11694
rect 5828 11665 5856 11698
rect 5724 11630 5776 11636
rect 5814 11656 5870 11665
rect 5814 11591 5870 11600
rect 5920 9466 5948 12974
rect 6012 10674 6040 14010
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5998 10432 6054 10441
rect 5998 10367 6054 10376
rect 5828 9438 5948 9466
rect 5828 9382 5856 9438
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5722 9208 5778 9217
rect 5722 9143 5724 9152
rect 5776 9143 5778 9152
rect 5724 9114 5776 9120
rect 5736 7818 5764 9114
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6662 5764 6734
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5354 5264 5410 5273
rect 5354 5199 5410 5208
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5460 2310 5488 3878
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5552 1630 5580 5510
rect 5630 4312 5686 4321
rect 5630 4247 5686 4256
rect 5644 3602 5672 4247
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5736 3534 5764 4082
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5828 3466 5856 9318
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5920 8566 5948 9114
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 6012 8362 6040 10367
rect 6104 8922 6132 11630
rect 6196 11529 6224 13874
rect 6288 11937 6316 14894
rect 6274 11928 6330 11937
rect 6274 11863 6330 11872
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6182 11520 6238 11529
rect 6182 11455 6238 11464
rect 6104 8894 6224 8922
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6104 8634 6132 8774
rect 6196 8650 6224 8894
rect 6288 8809 6316 11766
rect 6274 8800 6330 8809
rect 6274 8735 6330 8744
rect 6092 8628 6144 8634
rect 6196 8622 6316 8650
rect 6092 8570 6144 8576
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 6012 6798 6040 8298
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4078 6040 4966
rect 6288 4185 6316 8622
rect 6380 4486 6408 21082
rect 6656 18698 6684 32166
rect 9140 31822 9168 37062
rect 9864 34604 9916 34610
rect 9864 34546 9916 34552
rect 9876 32026 9904 34546
rect 10796 33522 10824 37062
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 10784 33516 10836 33522
rect 10784 33458 10836 33464
rect 10140 33312 10192 33318
rect 10140 33254 10192 33260
rect 9864 32020 9916 32026
rect 9864 31962 9916 31968
rect 8852 31816 8904 31822
rect 8852 31758 8904 31764
rect 9128 31816 9180 31822
rect 9128 31758 9180 31764
rect 9312 31816 9364 31822
rect 9312 31758 9364 31764
rect 7656 29640 7708 29646
rect 7656 29582 7708 29588
rect 7012 28416 7064 28422
rect 7012 28358 7064 28364
rect 7024 20058 7052 28358
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18358 7144 18566
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7208 17882 7236 18294
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6472 16658 6500 16934
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6932 16454 6960 16934
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6472 11694 6500 13330
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6564 10266 6592 14214
rect 6642 11928 6698 11937
rect 6642 11863 6698 11872
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6656 10146 6684 11863
rect 6748 11762 6776 14758
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12442 6868 12582
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6932 11830 6960 16390
rect 7024 16182 7052 17614
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 7208 15706 7236 16390
rect 7300 16114 7328 17138
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7024 12170 7052 15438
rect 7116 13326 7144 15574
rect 7300 13938 7328 16050
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7392 15162 7420 15438
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 14006 7420 14214
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7484 12918 7512 19110
rect 7668 18426 7696 29582
rect 8576 27328 8628 27334
rect 8576 27270 8628 27276
rect 8588 22642 8616 27270
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8220 22098 8248 22578
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7852 19854 7880 21966
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8024 21412 8076 21418
rect 8024 21354 8076 21360
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7760 18222 7788 19314
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7576 15162 7604 17070
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7576 13161 7604 13398
rect 7562 13152 7618 13161
rect 7562 13087 7618 13096
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6748 11218 6776 11562
rect 7024 11506 7052 11698
rect 6840 11478 7052 11506
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 10674 6776 11154
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6564 10118 6684 10146
rect 6748 10130 6776 10610
rect 6736 10124 6788 10130
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6472 9897 6500 9930
rect 6458 9888 6514 9897
rect 6458 9823 6514 9832
rect 6564 9466 6592 10118
rect 6736 10066 6788 10072
rect 6644 9580 6696 9586
rect 6748 9568 6776 10066
rect 6696 9540 6776 9568
rect 6644 9522 6696 9528
rect 6564 9438 6684 9466
rect 6458 7984 6514 7993
rect 6458 7919 6460 7928
rect 6512 7919 6514 7928
rect 6460 7890 6512 7896
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6472 5760 6500 6258
rect 6564 5914 6592 7482
rect 6656 5930 6684 9438
rect 6748 9382 6776 9540
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 8974 6776 9318
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8430 6776 8910
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 7342 6776 8366
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6748 6866 6776 7278
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 6254 6776 6802
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6840 6118 6868 11478
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6932 7546 6960 9930
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6552 5908 6604 5914
rect 6656 5902 6868 5930
rect 6552 5850 6604 5856
rect 6552 5772 6604 5778
rect 6472 5732 6552 5760
rect 6552 5714 6604 5720
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6564 4826 6592 4966
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6564 4690 6592 4762
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6458 4584 6514 4593
rect 6458 4519 6460 4528
rect 6512 4519 6514 4528
rect 6460 4490 6512 4496
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6380 4282 6408 4422
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6274 4176 6330 4185
rect 6274 4111 6330 4120
rect 6000 4072 6052 4078
rect 5906 4040 5962 4049
rect 6000 4014 6052 4020
rect 5906 3975 5962 3984
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5920 2990 5948 3975
rect 6012 3602 6040 4014
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5920 2582 5948 2926
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 6012 2514 6040 3538
rect 6748 2774 6776 5578
rect 6840 3369 6868 5902
rect 6918 5400 6974 5409
rect 7024 5370 7052 11018
rect 7116 10742 7144 12854
rect 7472 12776 7524 12782
rect 7378 12744 7434 12753
rect 7472 12718 7524 12724
rect 7378 12679 7434 12688
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7208 12102 7236 12310
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7208 11506 7236 12038
rect 7300 11830 7328 12038
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7208 11478 7328 11506
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7208 9654 7236 11290
rect 7300 9722 7328 11478
rect 7392 10266 7420 12679
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7286 8120 7342 8129
rect 7286 8055 7342 8064
rect 7300 8022 7328 8055
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7286 7304 7342 7313
rect 7286 7239 7288 7248
rect 7340 7239 7342 7248
rect 7288 7210 7340 7216
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7116 6390 7144 6802
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6390 7328 6598
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 6918 5335 6974 5344
rect 7012 5364 7064 5370
rect 6932 5302 6960 5335
rect 7012 5306 7064 5312
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6826 3360 6882 3369
rect 6826 3295 6882 3304
rect 6656 2746 6776 2774
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5816 1964 5868 1970
rect 5816 1906 5868 1912
rect 5540 1624 5592 1630
rect 5540 1566 5592 1572
rect 4540 1006 4660 1034
rect 5264 1080 5316 1086
rect 5264 1022 5316 1028
rect 4540 800 4568 1006
rect 5828 800 5856 1906
rect 6656 1018 6684 2746
rect 6826 2408 6882 2417
rect 6826 2343 6828 2352
rect 6880 2343 6882 2352
rect 6828 2314 6880 2320
rect 6932 2310 6960 5102
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 4146 7144 4490
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7116 3194 7144 4082
rect 7300 4010 7328 5578
rect 7484 5166 7512 12718
rect 7576 11218 7604 13087
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11218 7696 11494
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7668 6905 7696 10202
rect 7760 7478 7788 18158
rect 7852 17746 7880 19790
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7944 16658 7972 19654
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7852 15366 7880 16050
rect 8036 15994 8064 21354
rect 8772 20466 8800 21422
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8312 16658 8340 17478
rect 8588 17338 8616 18226
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 7944 15966 8064 15994
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7944 14498 7972 15966
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8036 15026 8064 15846
rect 8496 15638 8524 16662
rect 8680 16046 8708 18294
rect 8864 18170 8892 31758
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 9232 22094 9260 23122
rect 9140 22066 9260 22094
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 9048 21146 9076 21490
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8956 20466 8984 20742
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 9048 20330 9076 21082
rect 9036 20324 9088 20330
rect 9036 20266 9088 20272
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 9048 18426 9076 18634
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8864 18142 9076 18170
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8864 17202 8892 17682
rect 8956 17202 8984 18022
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 8206 15192 8262 15201
rect 8404 15162 8432 15370
rect 8206 15127 8262 15136
rect 8392 15156 8444 15162
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 7852 14470 7972 14498
rect 7852 12782 7880 14470
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 7944 14074 7972 14350
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 8036 12306 8064 13806
rect 8128 13530 8156 14350
rect 8220 13818 8248 15127
rect 8392 15098 8444 15104
rect 8496 14550 8524 15574
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8588 14482 8616 14758
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8484 14000 8536 14006
rect 8484 13942 8536 13948
rect 8220 13790 8340 13818
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8220 13326 8248 13670
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8312 13172 8340 13790
rect 8128 13144 8340 13172
rect 8128 12374 8156 13144
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8312 12434 8340 12786
rect 8312 12406 8432 12434
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7838 10296 7894 10305
rect 7838 10231 7894 10240
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7760 7002 7788 7414
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7654 6896 7710 6905
rect 7654 6831 7710 6840
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7484 3058 7512 4014
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7484 2514 7512 2994
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7576 1154 7604 6666
rect 7852 6662 7880 10231
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7668 3913 7696 4150
rect 7654 3904 7710 3913
rect 7654 3839 7710 3848
rect 7656 2848 7708 2854
rect 7654 2816 7656 2825
rect 7708 2816 7710 2825
rect 7654 2751 7710 2760
rect 7564 1148 7616 1154
rect 7564 1090 7616 1096
rect 6644 1012 6696 1018
rect 6644 954 6696 960
rect 7760 800 7788 4558
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7852 2553 7880 3402
rect 7944 3233 7972 11698
rect 8114 11520 8170 11529
rect 8114 11455 8170 11464
rect 8128 7478 8156 11455
rect 8312 9994 8340 12174
rect 8404 10810 8432 12406
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8496 9874 8524 13942
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8588 11218 8616 13874
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8772 12782 8800 13398
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8312 9846 8524 9874
rect 8208 9648 8260 9654
rect 8206 9616 8208 9625
rect 8260 9616 8262 9625
rect 8206 9551 8262 9560
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8673 8248 8910
rect 8206 8664 8262 8673
rect 8206 8599 8262 8608
rect 8312 7954 8340 9846
rect 8588 9654 8616 11154
rect 8680 10418 8708 11630
rect 8772 10606 8800 12718
rect 8864 10674 8892 17138
rect 9048 16590 9076 18142
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9048 13569 9076 16526
rect 9034 13560 9090 13569
rect 9034 13495 9090 13504
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8680 10390 8800 10418
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8496 9110 8524 9454
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 8401 8432 8434
rect 8390 8392 8446 8401
rect 8390 8327 8446 8336
rect 8588 8129 8616 8774
rect 8574 8120 8630 8129
rect 8574 8055 8630 8064
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8128 6662 8156 7414
rect 8220 7342 8248 7686
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8312 6769 8340 7754
rect 8576 7744 8628 7750
rect 8496 7704 8576 7732
rect 8298 6760 8354 6769
rect 8298 6695 8354 6704
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8036 5710 8064 6258
rect 8206 5808 8262 5817
rect 8206 5743 8262 5752
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8220 5302 8248 5743
rect 8496 5710 8524 7704
rect 8576 7686 8628 7692
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 5914 8616 6598
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8404 4826 8432 5578
rect 8680 5574 8708 9862
rect 8772 8974 8800 10390
rect 8864 9722 8892 10474
rect 8956 10062 8984 12922
rect 9140 11354 9168 22066
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9232 19417 9260 19790
rect 9218 19408 9274 19417
rect 9218 19343 9220 19352
rect 9272 19343 9274 19352
rect 9220 19314 9272 19320
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9232 17882 9260 18226
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9324 17134 9352 31758
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9324 15706 9352 16118
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9416 14074 9444 14894
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9508 13705 9536 23598
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9600 20534 9628 23462
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9784 21010 9812 21286
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 10060 20874 10088 21490
rect 10048 20868 10100 20874
rect 10048 20810 10100 20816
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9876 19854 9904 20334
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9692 18426 9720 18634
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9784 17746 9812 18838
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16454 9720 16934
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9692 15570 9720 16390
rect 9784 16250 9812 17546
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9772 15496 9824 15502
rect 9876 15484 9904 16050
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9824 15456 9904 15484
rect 9772 15438 9824 15444
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9600 13938 9628 14282
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9494 13696 9550 13705
rect 9494 13631 9550 13640
rect 9692 13530 9720 15370
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9048 10606 9076 11154
rect 9232 11121 9260 13330
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 11150 9352 13126
rect 9508 12986 9536 13262
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9312 11144 9364 11150
rect 9218 11112 9274 11121
rect 9128 11076 9180 11082
rect 9312 11086 9364 11092
rect 9218 11047 9274 11056
rect 9128 11018 9180 11024
rect 9140 10810 9168 11018
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 9048 10130 9076 10542
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 6118 8800 8774
rect 8864 7546 8892 9658
rect 9048 9518 9076 10066
rect 9140 9926 9168 10610
rect 9218 10160 9274 10169
rect 9218 10095 9274 10104
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 9382 9076 9454
rect 9036 9376 9088 9382
rect 9232 9330 9260 10095
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9324 9382 9352 9998
rect 9036 9318 9088 9324
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8956 7206 8984 8910
rect 9048 8498 9076 9318
rect 9140 9302 9260 9330
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9140 8378 9168 9302
rect 9218 9208 9274 9217
rect 9416 9178 9444 9998
rect 9508 9353 9536 12242
rect 9600 12170 9628 12582
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9600 11694 9628 12106
rect 9692 12073 9720 12106
rect 9678 12064 9734 12073
rect 9678 11999 9734 12008
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9784 11014 9812 13874
rect 9876 12306 9904 15456
rect 9968 12442 9996 15846
rect 9956 12436 10008 12442
rect 10060 12434 10088 20810
rect 10152 20466 10180 33254
rect 10876 31816 10928 31822
rect 10876 31758 10928 31764
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10336 20466 10364 21830
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10520 21457 10548 21490
rect 10506 21448 10562 21457
rect 10506 21383 10562 21392
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10520 19310 10548 19994
rect 10612 19718 10640 20198
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10612 18970 10640 19314
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10140 17808 10192 17814
rect 10140 17750 10192 17756
rect 10152 13870 10180 17750
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10244 17338 10272 17546
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10230 16960 10286 16969
rect 10230 16895 10286 16904
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10152 13326 10180 13806
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10244 13258 10272 16895
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10428 15502 10456 16526
rect 10796 16250 10824 18702
rect 10888 17746 10916 31758
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10980 21010 11008 21830
rect 11164 21690 11192 21966
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 11256 20942 11284 21898
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11532 19854 11560 21966
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11624 20466 11652 21830
rect 11716 21554 11744 34886
rect 11992 34610 12020 37130
rect 14844 37126 14872 39200
rect 16132 39114 16160 39200
rect 16224 39114 16252 39222
rect 16132 39086 16252 39114
rect 14924 37256 14976 37262
rect 14924 37198 14976 37204
rect 12992 37120 13044 37126
rect 12992 37062 13044 37068
rect 14832 37120 14884 37126
rect 14832 37062 14884 37068
rect 13004 35086 13032 37062
rect 14936 35290 14964 37198
rect 16500 37108 16528 39222
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 20626 39200 20682 39800
rect 22558 39200 22614 39800
rect 23846 39200 23902 39800
rect 25778 39200 25834 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 31574 39200 31630 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 16580 37120 16632 37126
rect 16500 37080 16580 37108
rect 16580 37062 16632 37068
rect 16868 35290 16896 37198
rect 18064 37126 18092 39200
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 18156 35290 18184 37198
rect 19352 37126 19380 39200
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 20640 37210 20668 39200
rect 22572 37262 22600 39200
rect 20720 37256 20772 37262
rect 20640 37204 20720 37210
rect 20640 37198 20772 37204
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 22928 37256 22980 37262
rect 22928 37198 22980 37204
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 14924 35284 14976 35290
rect 14924 35226 14976 35232
rect 16856 35284 16908 35290
rect 16856 35226 16908 35232
rect 18144 35284 18196 35290
rect 18144 35226 18196 35232
rect 12992 35080 13044 35086
rect 12992 35022 13044 35028
rect 15660 35080 15712 35086
rect 15660 35022 15712 35028
rect 16672 35080 16724 35086
rect 16672 35022 16724 35028
rect 17592 35080 17644 35086
rect 17592 35022 17644 35028
rect 11980 34604 12032 34610
rect 11980 34546 12032 34552
rect 12164 34536 12216 34542
rect 12164 34478 12216 34484
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 12084 22642 12112 22918
rect 12072 22636 12124 22642
rect 12072 22578 12124 22584
rect 12176 21554 12204 34478
rect 15672 30326 15700 35022
rect 16684 30938 16712 35022
rect 16672 30932 16724 30938
rect 16672 30874 16724 30880
rect 17408 30728 17460 30734
rect 17408 30670 17460 30676
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 12900 23520 12952 23526
rect 12900 23462 12952 23468
rect 12912 23118 12940 23462
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 13188 23050 13216 23666
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23118 15240 23462
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12728 22098 12756 22918
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13280 22234 13308 22374
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 12084 21078 12112 21286
rect 12268 21146 12296 21966
rect 13372 21690 13400 23054
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15706 10732 15846
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10612 14074 10640 15438
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10704 14618 10732 14894
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10060 12406 10180 12434
rect 9956 12378 10008 12384
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9680 11008 9732 11014
rect 9678 10976 9680 10985
rect 9772 11008 9824 11014
rect 9732 10976 9734 10985
rect 9772 10950 9824 10956
rect 9678 10911 9734 10920
rect 9680 10464 9732 10470
rect 9784 10452 9812 10950
rect 9732 10424 9812 10452
rect 9680 10406 9732 10412
rect 9954 10024 10010 10033
rect 10152 9994 10180 12406
rect 10336 12238 10364 13670
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12782 10456 13262
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10520 12850 10548 13126
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10416 12776 10468 12782
rect 10468 12724 10548 12730
rect 10416 12718 10548 12724
rect 10428 12702 10548 12718
rect 10428 12653 10456 12702
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10428 12050 10456 12242
rect 10336 12022 10456 12050
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9954 9959 10010 9968
rect 10140 9988 10192 9994
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9494 9344 9550 9353
rect 9494 9279 9550 9288
rect 9218 9143 9220 9152
rect 9272 9143 9274 9152
rect 9404 9172 9456 9178
rect 9220 9114 9272 9120
rect 9404 9114 9456 9120
rect 9218 8936 9274 8945
rect 9218 8871 9274 8880
rect 9048 8350 9168 8378
rect 9232 8362 9260 8871
rect 9600 8838 9628 9590
rect 9678 9344 9734 9353
rect 9678 9279 9734 9288
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9692 8514 9720 9279
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9784 8566 9812 8910
rect 9876 8838 9904 8978
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9600 8486 9720 8514
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9600 8412 9628 8486
rect 9416 8384 9628 8412
rect 9220 8356 9272 8362
rect 9048 7750 9076 8350
rect 9220 8298 9272 8304
rect 9312 8288 9364 8294
rect 9416 8276 9444 8384
rect 9364 8248 9444 8276
rect 9588 8288 9640 8294
rect 9312 8230 9364 8236
rect 9588 8230 9640 8236
rect 9600 8129 9628 8230
rect 9126 8120 9182 8129
rect 9126 8055 9182 8064
rect 9586 8120 9642 8129
rect 9586 8055 9642 8064
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 9048 5302 9076 7482
rect 9140 5710 9168 8055
rect 9586 7984 9642 7993
rect 9312 7948 9364 7954
rect 9586 7919 9642 7928
rect 9312 7890 9364 7896
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9324 7834 9352 7890
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 9232 4978 9260 7822
rect 9324 7806 9444 7834
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 5914 9352 7686
rect 9416 6118 9444 7806
rect 9494 7032 9550 7041
rect 9494 6967 9550 6976
rect 9508 6662 9536 6967
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9600 5914 9628 7919
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9692 5574 9720 8486
rect 9784 7954 9812 8502
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9784 6866 9812 7890
rect 9968 7886 9996 9959
rect 10140 9930 10192 9936
rect 10152 8634 10180 9930
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10060 8129 10088 8502
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10046 8120 10102 8129
rect 10046 8055 10102 8064
rect 10152 7993 10180 8230
rect 10138 7984 10194 7993
rect 10138 7919 10194 7928
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9968 7410 9996 7822
rect 10244 7818 10272 11630
rect 10336 11558 10364 12022
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10336 9042 10364 11494
rect 10428 11218 10456 11494
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10428 10470 10456 11018
rect 10520 10577 10548 12702
rect 10506 10568 10562 10577
rect 10506 10503 10562 10512
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10428 8906 10456 9386
rect 10520 9353 10548 10503
rect 10612 9586 10640 13874
rect 10704 13190 10732 14350
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10704 12050 10732 12582
rect 10796 12434 10824 16186
rect 10888 16182 10916 17682
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10980 17202 11008 17614
rect 11072 17338 11100 19246
rect 11244 19236 11296 19242
rect 11244 19178 11296 19184
rect 11336 19236 11388 19242
rect 11336 19178 11388 19184
rect 11256 18222 11284 19178
rect 11348 18358 11376 19178
rect 11336 18352 11388 18358
rect 11336 18294 11388 18300
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 11428 17060 11480 17066
rect 11428 17002 11480 17008
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 10980 15014 11284 15042
rect 10980 14890 11008 15014
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 11072 14618 11100 14826
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10888 12714 10916 13330
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10796 12406 10916 12434
rect 10704 12022 10824 12050
rect 10796 11694 10824 12022
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10782 11520 10838 11529
rect 10782 11455 10838 11464
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10506 9344 10562 9353
rect 10506 9279 10562 9288
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10506 8800 10562 8809
rect 10506 8735 10562 8744
rect 10520 8634 10548 8735
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10612 8378 10640 9522
rect 10428 8350 10640 8378
rect 10322 7984 10378 7993
rect 10322 7919 10378 7928
rect 10336 7818 10364 7919
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 6458 9904 6734
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 10060 6254 10088 6938
rect 10336 6866 10364 7346
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10244 6633 10272 6666
rect 10230 6624 10286 6633
rect 10230 6559 10286 6568
rect 10336 6254 10364 6802
rect 10428 6746 10456 8350
rect 10506 8256 10562 8265
rect 10506 8191 10562 8200
rect 10520 7342 10548 8191
rect 10598 7576 10654 7585
rect 10598 7511 10600 7520
rect 10652 7511 10654 7520
rect 10600 7482 10652 7488
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10428 6730 10548 6746
rect 10428 6724 10560 6730
rect 10428 6718 10508 6724
rect 10508 6666 10560 6672
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10336 5778 10364 6190
rect 10520 6089 10548 6666
rect 10506 6080 10562 6089
rect 10506 6015 10562 6024
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9232 4950 9536 4978
rect 8942 4856 8998 4865
rect 8392 4820 8444 4826
rect 8942 4791 8998 4800
rect 9402 4856 9458 4865
rect 9402 4791 9404 4800
rect 8392 4762 8444 4768
rect 8298 4720 8354 4729
rect 8956 4690 8984 4791
rect 9456 4791 9458 4800
rect 9404 4762 9456 4768
rect 9402 4720 9458 4729
rect 8298 4655 8354 4664
rect 8944 4684 8996 4690
rect 8312 4622 8340 4655
rect 9402 4655 9404 4664
rect 8944 4626 8996 4632
rect 9456 4655 9458 4664
rect 9404 4626 9456 4632
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 9036 4616 9088 4622
rect 9312 4616 9364 4622
rect 9088 4576 9312 4604
rect 9036 4558 9088 4564
rect 9312 4558 9364 4564
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8036 3534 8064 4218
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7930 3224 7986 3233
rect 7930 3159 7986 3168
rect 8116 3120 8168 3126
rect 8168 3068 8340 3074
rect 8116 3062 8340 3068
rect 8128 3046 8340 3062
rect 7838 2544 7894 2553
rect 7838 2479 7894 2488
rect 8312 1834 8340 3046
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8496 2038 8524 2314
rect 8484 2032 8536 2038
rect 8484 1974 8536 1980
rect 8300 1828 8352 1834
rect 8300 1770 8352 1776
rect 8588 1426 8616 2314
rect 8576 1420 8628 1426
rect 8576 1362 8628 1368
rect 9048 800 9076 4422
rect 9310 4176 9366 4185
rect 9310 4111 9312 4120
rect 9364 4111 9366 4120
rect 9312 4082 9364 4088
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9324 2514 9352 3470
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9508 2145 9536 4950
rect 9600 4842 9628 5510
rect 10336 5370 10364 5714
rect 10704 5642 10732 10678
rect 10796 5914 10824 11455
rect 10888 6186 10916 12406
rect 10980 11218 11008 13874
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13394 11100 13670
rect 11164 13462 11192 14758
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 11072 10033 11100 13126
rect 11164 10538 11192 13126
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11058 10024 11114 10033
rect 11058 9959 11114 9968
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11072 8809 11100 9114
rect 11058 8800 11114 8809
rect 11058 8735 11114 8744
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10980 7410 11008 8366
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 8090 11100 8230
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11060 7472 11112 7478
rect 11058 7440 11060 7449
rect 11112 7440 11114 7449
rect 10968 7404 11020 7410
rect 11058 7375 11114 7384
rect 10968 7346 11020 7352
rect 11164 7274 11192 9318
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10782 5672 10838 5681
rect 10692 5636 10744 5642
rect 10782 5607 10784 5616
rect 10692 5578 10744 5584
rect 10836 5607 10838 5616
rect 10784 5578 10836 5584
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 9600 4814 9812 4842
rect 9678 4720 9734 4729
rect 9678 4655 9734 4664
rect 9588 4208 9640 4214
rect 9586 4176 9588 4185
rect 9640 4176 9642 4185
rect 9586 4111 9642 4120
rect 9692 4078 9720 4655
rect 9784 4214 9812 4814
rect 10336 4690 10364 5306
rect 10520 5030 10548 5510
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9968 4078 9996 4558
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 9680 4072 9732 4078
rect 9772 4072 9824 4078
rect 9680 4014 9732 4020
rect 9770 4040 9772 4049
rect 9956 4072 10008 4078
rect 9824 4040 9826 4049
rect 9956 4014 10008 4020
rect 9770 3975 9826 3984
rect 9770 3768 9826 3777
rect 9770 3703 9826 3712
rect 9784 3602 9812 3703
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9784 2650 9812 3402
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 9494 2136 9550 2145
rect 9494 2071 9550 2080
rect 9600 1698 9628 2314
rect 9968 2106 9996 2926
rect 10060 2378 10088 4422
rect 10152 3618 10180 4626
rect 10506 4448 10562 4457
rect 10506 4383 10562 4392
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10244 3738 10272 3946
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10336 3738 10364 3878
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10152 3590 10364 3618
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10152 2854 10180 2994
rect 10140 2848 10192 2854
rect 10244 2825 10272 3062
rect 10140 2790 10192 2796
rect 10230 2816 10286 2825
rect 10230 2751 10286 2760
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 9588 1692 9640 1698
rect 9588 1634 9640 1640
rect 10336 800 10364 3590
rect 10428 3398 10456 3878
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10520 2990 10548 4383
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10704 3126 10732 3334
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10796 2258 10824 5578
rect 10888 2378 10916 6122
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10980 5409 11008 5850
rect 10966 5400 11022 5409
rect 10966 5335 11022 5344
rect 10980 4554 11008 5335
rect 11072 5114 11100 6258
rect 11164 5953 11192 6666
rect 11150 5944 11206 5953
rect 11256 5914 11284 15014
rect 11348 13190 11376 15302
rect 11440 13802 11468 17002
rect 11532 15201 11560 19790
rect 11704 18624 11756 18630
rect 11808 18612 11836 19790
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12820 19242 12848 19722
rect 13004 19446 13032 19994
rect 13268 19984 13320 19990
rect 13268 19926 13320 19932
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12268 18970 12296 19110
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 11756 18584 11836 18612
rect 11704 18566 11756 18572
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11808 17270 11836 18226
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11612 17060 11664 17066
rect 11612 17002 11664 17008
rect 11624 16794 11652 17002
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11808 16454 11836 16526
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11518 15192 11574 15201
rect 11518 15127 11574 15136
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11348 12753 11376 12854
rect 11334 12744 11390 12753
rect 11334 12679 11390 12688
rect 11440 12434 11468 13262
rect 11532 13190 11560 14350
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11348 12406 11468 12434
rect 11348 11257 11376 12406
rect 11532 12322 11560 13126
rect 11624 12374 11652 15982
rect 11992 15688 12020 18838
rect 12532 18624 12584 18630
rect 12584 18572 12848 18578
rect 12532 18566 12848 18572
rect 12544 18550 12848 18566
rect 12254 18184 12310 18193
rect 12530 18184 12586 18193
rect 12254 18119 12256 18128
rect 12308 18119 12310 18128
rect 12348 18148 12400 18154
rect 12256 18090 12308 18096
rect 12530 18119 12532 18128
rect 12348 18090 12400 18096
rect 12584 18119 12586 18128
rect 12532 18090 12584 18096
rect 12360 17678 12388 18090
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12452 16794 12480 17138
rect 12728 16810 12756 17614
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12636 16782 12756 16810
rect 12636 16250 12664 16782
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 11808 15660 12020 15688
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11716 14618 11744 15030
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11716 13326 11744 13738
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11716 12850 11744 13262
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11440 12294 11560 12322
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11334 11248 11390 11257
rect 11334 11183 11390 11192
rect 11348 9194 11376 11183
rect 11440 9382 11468 12294
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11532 11286 11560 12174
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11702 11112 11758 11121
rect 11702 11047 11704 11056
rect 11756 11047 11758 11056
rect 11704 11018 11756 11024
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11518 9888 11574 9897
rect 11518 9823 11574 9832
rect 11532 9674 11560 9823
rect 11716 9722 11744 9930
rect 11704 9716 11756 9722
rect 11532 9646 11652 9674
rect 11704 9658 11756 9664
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11348 9166 11468 9194
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11348 6866 11376 8842
rect 11440 8514 11468 9166
rect 11624 9110 11652 9646
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11440 8486 11560 8514
rect 11428 8016 11480 8022
rect 11426 7984 11428 7993
rect 11480 7984 11482 7993
rect 11426 7919 11482 7928
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11440 7721 11468 7822
rect 11426 7712 11482 7721
rect 11426 7647 11482 7656
rect 11426 7168 11482 7177
rect 11426 7103 11482 7112
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11440 6746 11468 7103
rect 11532 7041 11560 8486
rect 11518 7032 11574 7041
rect 11518 6967 11574 6976
rect 11348 6718 11468 6746
rect 11150 5879 11206 5888
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11072 5086 11192 5114
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 11072 4146 11100 4966
rect 11164 4865 11192 5086
rect 11150 4856 11206 4865
rect 11150 4791 11206 4800
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 11072 3942 11100 3975
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11348 2774 11376 6718
rect 11624 6644 11652 9046
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11716 7206 11744 7822
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11440 6616 11652 6644
rect 11440 6322 11468 6616
rect 11808 6610 11836 15660
rect 12072 15496 12124 15502
rect 12124 15456 12204 15484
rect 12072 15438 12124 15444
rect 12176 14958 12204 15456
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 11900 13002 11928 14894
rect 12176 14822 12204 14894
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12360 14618 12388 16050
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12452 13870 12480 15914
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12544 15162 12572 15642
rect 12636 15570 12664 15846
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12728 15502 12756 16594
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11992 13190 12020 13262
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11900 12974 12020 13002
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11900 12306 11928 12786
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11992 11558 12020 12974
rect 12084 12889 12112 13738
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12176 13190 12204 13670
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12452 13190 12480 13330
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12532 12912 12584 12918
rect 12070 12880 12126 12889
rect 12532 12854 12584 12860
rect 12070 12815 12126 12824
rect 12440 12436 12492 12442
rect 12544 12434 12572 12854
rect 12492 12406 12572 12434
rect 12440 12378 12492 12384
rect 12636 12306 12664 13126
rect 12728 12628 12756 14418
rect 12820 12782 12848 18550
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13004 17746 13032 18226
rect 13096 18086 13124 19314
rect 13280 19174 13308 19926
rect 13372 19802 13400 21626
rect 13464 21554 13492 22918
rect 13728 22500 13780 22506
rect 13728 22442 13780 22448
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13740 21418 13768 22442
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 13832 21321 13860 22102
rect 13818 21312 13874 21321
rect 13818 21247 13874 21256
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13740 19922 13768 20198
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13832 19854 13860 20810
rect 14016 20466 14044 22986
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14384 22642 14412 22918
rect 14568 22778 14596 23054
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 15028 22778 15056 22918
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14464 22432 14516 22438
rect 14464 22374 14516 22380
rect 14476 21962 14504 22374
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 13820 19848 13872 19854
rect 13372 19774 13768 19802
rect 13820 19790 13872 19796
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13372 18902 13400 19110
rect 13464 18902 13492 19654
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13372 18222 13400 18362
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13004 16522 13032 17682
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12912 13530 12940 13806
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12728 12600 12940 12628
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12440 12232 12492 12238
rect 12492 12180 12572 12186
rect 12440 12174 12572 12180
rect 12256 12164 12308 12170
rect 12452 12158 12572 12174
rect 12256 12106 12308 12112
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11886 10976 11942 10985
rect 11886 10911 11942 10920
rect 11900 10198 11928 10911
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11992 10062 12020 11494
rect 12084 10266 12112 11698
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 12070 9888 12126 9897
rect 12070 9823 12126 9832
rect 12084 9654 12112 9823
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 11886 9208 11942 9217
rect 11886 9143 11942 9152
rect 11900 8974 11928 9143
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11978 8800 12034 8809
rect 11978 8735 12034 8744
rect 11992 8430 12020 8735
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12070 7984 12126 7993
rect 12070 7919 12072 7928
rect 12124 7919 12126 7928
rect 12072 7890 12124 7896
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11978 7576 12034 7585
rect 11978 7511 12034 7520
rect 11992 7478 12020 7511
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11716 6582 11836 6610
rect 11716 6474 11744 6582
rect 11532 6446 11744 6474
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11440 5574 11468 6258
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11440 3466 11468 4014
rect 11532 3602 11560 6446
rect 11900 6304 11928 6967
rect 12084 6934 12112 7686
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11992 6458 12020 6666
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11624 6276 11928 6304
rect 11624 6186 11652 6276
rect 11980 6248 12032 6254
rect 12084 6236 12112 6598
rect 12032 6208 12112 6236
rect 11980 6190 12032 6196
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11704 6112 11756 6118
rect 11992 6100 12020 6190
rect 11756 6072 12020 6100
rect 11704 6054 11756 6060
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11610 5536 11666 5545
rect 11610 5471 11666 5480
rect 11624 5098 11652 5471
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11716 5234 11744 5306
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11716 4146 11744 5170
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11716 3602 11744 4082
rect 11900 4060 11928 5850
rect 12084 5778 12112 5850
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 11992 4282 12020 5238
rect 12176 4457 12204 10950
rect 12268 9654 12296 12106
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11898 12480 12038
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12544 11234 12572 12158
rect 12636 11898 12664 12242
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12544 11206 12756 11234
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12346 10976 12402 10985
rect 12346 10911 12402 10920
rect 12360 10169 12388 10911
rect 12438 10840 12494 10849
rect 12438 10775 12494 10784
rect 12452 10742 12480 10775
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12544 10690 12572 11086
rect 12544 10662 12664 10690
rect 12346 10160 12402 10169
rect 12346 10095 12402 10104
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12254 8800 12310 8809
rect 12254 8735 12310 8744
rect 12268 8566 12296 8735
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12254 8256 12310 8265
rect 12254 8191 12310 8200
rect 12268 5302 12296 8191
rect 12360 5778 12388 9386
rect 12544 9217 12572 9454
rect 12530 9208 12586 9217
rect 12530 9143 12586 9152
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12452 7886 12480 8230
rect 12544 7993 12572 8230
rect 12530 7984 12586 7993
rect 12530 7919 12586 7928
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12346 5400 12402 5409
rect 12346 5335 12402 5344
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12360 4758 12388 5335
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12162 4448 12218 4457
rect 12162 4383 12218 4392
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11980 4072 12032 4078
rect 11900 4032 11980 4060
rect 11980 4014 12032 4020
rect 11978 3904 12034 3913
rect 12084 3890 12112 4218
rect 12268 4214 12296 4558
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12034 3862 12112 3890
rect 11978 3839 12034 3848
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11532 3126 11560 3538
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11716 3058 11744 3538
rect 12268 3466 12296 4150
rect 12636 4060 12664 10662
rect 12728 8090 12756 11206
rect 12820 10130 12848 12242
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12728 7818 12756 7890
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12728 6089 12756 6394
rect 12714 6080 12770 6089
rect 12714 6015 12770 6024
rect 12714 5672 12770 5681
rect 12714 5607 12770 5616
rect 12728 4554 12756 5607
rect 12820 5409 12848 9590
rect 12912 5545 12940 12600
rect 13004 12306 13032 16458
rect 13096 15484 13124 16526
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13188 15706 13216 15846
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13176 15496 13228 15502
rect 13096 15456 13176 15484
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 13096 11286 13124 15456
rect 13176 15438 13228 15444
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 11898 13216 15302
rect 13280 13802 13308 17138
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13372 16114 13400 16662
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13464 15638 13492 15982
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13280 13138 13308 13466
rect 13280 13110 13400 13138
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13280 12170 13308 12718
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13372 11778 13400 13110
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13188 11750 13400 11778
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13188 11014 13216 11750
rect 13464 11694 13492 12106
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13372 11354 13400 11630
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13176 10600 13228 10606
rect 13174 10568 13176 10577
rect 13228 10568 13230 10577
rect 13174 10503 13230 10512
rect 13280 10266 13308 11086
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13358 10568 13414 10577
rect 13358 10503 13414 10512
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12898 5536 12954 5545
rect 12898 5471 12954 5480
rect 12806 5400 12862 5409
rect 12806 5335 12862 5344
rect 13004 4690 13032 7482
rect 13096 6798 13124 10202
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13188 8265 13216 10066
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 9042 13308 9318
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13174 8256 13230 8265
rect 13174 8191 13230 8200
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13188 6866 13216 7822
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13084 6792 13136 6798
rect 13136 6740 13216 6746
rect 13084 6734 13216 6740
rect 13096 6718 13216 6734
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13096 5778 13124 6598
rect 13188 6089 13216 6718
rect 13174 6080 13230 6089
rect 13174 6015 13230 6024
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12452 4032 12664 4060
rect 12452 3942 12480 4032
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12176 3346 12204 3402
rect 12544 3369 12572 3878
rect 12530 3360 12586 3369
rect 12176 3318 12388 3346
rect 12360 3194 12388 3318
rect 12530 3295 12586 3304
rect 12990 3360 13046 3369
rect 12990 3295 13046 3304
rect 13004 3194 13032 3295
rect 13372 3194 13400 10503
rect 13464 9382 13492 10678
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13556 9110 13584 17682
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13648 15978 13676 16526
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13648 15366 13676 15914
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13648 14074 13676 14214
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13740 13954 13768 19774
rect 13924 19514 13952 20402
rect 14002 20360 14058 20369
rect 14002 20295 14058 20304
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13912 19304 13964 19310
rect 14016 19292 14044 20295
rect 14280 19780 14332 19786
rect 14280 19722 14332 19728
rect 13964 19264 14044 19292
rect 13912 19246 13964 19252
rect 13832 18630 13860 19246
rect 14016 18834 14044 19264
rect 14292 18834 14320 19722
rect 14384 19174 14412 20402
rect 14476 20058 14504 20878
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13832 17882 13860 18566
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14346 13860 14962
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13648 13926 13768 13954
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13648 13530 13676 13926
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12714 13676 13126
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 9897 13676 10406
rect 13634 9888 13690 9897
rect 13634 9823 13690 9832
rect 13740 9674 13768 13738
rect 13832 11830 13860 13942
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13924 11354 13952 14350
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14016 12102 14044 14282
rect 14108 14006 14136 18022
rect 14384 17270 14412 18226
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 14476 17134 14504 17750
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14292 14929 14320 17070
rect 14568 16266 14596 22714
rect 15488 22506 15516 23666
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15476 22500 15528 22506
rect 15476 22442 15528 22448
rect 15672 21554 15700 22918
rect 15752 22568 15804 22574
rect 15752 22510 15804 22516
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15108 20800 15160 20806
rect 15108 20742 15160 20748
rect 15120 20466 15148 20742
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 14936 19514 14964 20266
rect 15028 19854 15056 20402
rect 15212 20262 15240 21082
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15488 19854 15516 21422
rect 15580 20942 15608 21422
rect 15764 21418 15792 22510
rect 15856 21690 15884 23054
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 15292 19440 15344 19446
rect 15292 19382 15344 19388
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14936 19174 14964 19314
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 15304 18222 15332 19382
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14844 17678 14872 18022
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15304 17270 15332 18158
rect 15396 17746 15424 19722
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15488 17066 15516 17546
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15580 16946 15608 20878
rect 15948 20602 15976 20878
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15488 16918 15608 16946
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14384 16238 14596 16266
rect 14278 14920 14334 14929
rect 14278 14855 14334 14864
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 14096 13864 14148 13870
rect 14148 13824 14228 13852
rect 14096 13806 14148 13812
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14108 11914 14136 12718
rect 14016 11886 14136 11914
rect 14200 11898 14228 13824
rect 14292 12782 14320 14855
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14188 11892 14240 11898
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13832 10062 13860 10202
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13648 9646 13768 9674
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13450 8936 13506 8945
rect 13450 8871 13506 8880
rect 13464 8430 13492 8871
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 8430 13584 8774
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13648 8106 13676 9646
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13740 8265 13768 8502
rect 13726 8256 13782 8265
rect 13726 8191 13782 8200
rect 13556 8078 13676 8106
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13464 7342 13492 7482
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13464 7002 13492 7142
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13450 6624 13506 6633
rect 13450 6559 13506 6568
rect 13464 6186 13492 6559
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 13464 4457 13492 5238
rect 13556 5166 13584 8078
rect 13832 7886 13860 8774
rect 13820 7880 13872 7886
rect 13726 7848 13782 7857
rect 13820 7822 13872 7828
rect 13726 7783 13782 7792
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7002 13676 7686
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13634 5400 13690 5409
rect 13634 5335 13690 5344
rect 13648 5302 13676 5335
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13556 4729 13584 5102
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13542 4720 13598 4729
rect 13542 4655 13598 4664
rect 13648 4604 13676 4966
rect 13556 4576 13676 4604
rect 13740 4604 13768 7783
rect 13924 6390 13952 11154
rect 14016 8294 14044 11886
rect 14188 11834 14240 11840
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 9926 14136 11494
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 14016 7177 14044 7414
rect 14002 7168 14058 7177
rect 14002 7103 14058 7112
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5778 13860 6054
rect 13924 5778 13952 6190
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13832 4758 13860 5034
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13924 4690 13952 5510
rect 14108 5166 14136 9862
rect 14200 8242 14228 11562
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14292 10146 14320 11290
rect 14384 10577 14412 16238
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14568 15162 14596 15846
rect 14752 15434 14780 16390
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14740 15428 14792 15434
rect 14740 15370 14792 15376
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14922 14648 14978 14657
rect 14832 14612 14884 14618
rect 15028 14618 15056 15506
rect 14922 14583 14978 14592
rect 15016 14612 15068 14618
rect 14832 14554 14884 14560
rect 14844 13938 14872 14554
rect 14936 14414 14964 14583
rect 15016 14554 15068 14560
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15028 14006 15056 14214
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14556 13728 14608 13734
rect 15120 13705 15148 14554
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 14556 13670 14608 13676
rect 15106 13696 15162 13705
rect 14568 13530 14596 13670
rect 15106 13631 15162 13640
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 14476 11762 14504 13398
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14554 12744 14610 12753
rect 14554 12679 14610 12688
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14568 11694 14596 12679
rect 14936 12442 14964 13330
rect 15108 13320 15160 13326
rect 15028 13280 15108 13308
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 15028 12322 15056 13280
rect 15108 13262 15160 13268
rect 15304 12986 15332 13738
rect 15396 13530 15424 13806
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 14844 12294 15056 12322
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14462 10840 14518 10849
rect 14462 10775 14464 10784
rect 14516 10775 14518 10784
rect 14464 10746 14516 10752
rect 14370 10568 14426 10577
rect 14370 10503 14426 10512
rect 14476 10266 14596 10282
rect 14660 10266 14688 12174
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11762 14780 12038
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14464 10260 14596 10266
rect 14516 10254 14596 10260
rect 14464 10202 14516 10208
rect 14568 10146 14596 10254
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14752 10146 14780 11698
rect 14844 11626 14872 12294
rect 15016 11892 15068 11898
rect 14936 11852 15016 11880
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14844 11529 14872 11562
rect 14830 11520 14886 11529
rect 14830 11455 14886 11464
rect 14830 11248 14886 11257
rect 14830 11183 14886 11192
rect 14844 11150 14872 11183
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14292 10118 14504 10146
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14292 9722 14320 9998
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14384 9654 14412 9862
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 14292 8362 14320 8842
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14200 8214 14320 8242
rect 14292 6798 14320 8214
rect 14370 7848 14426 7857
rect 14370 7783 14426 7792
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14384 6730 14412 7783
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13740 4576 13860 4604
rect 13450 4448 13506 4457
rect 13450 4383 13506 4392
rect 13556 4298 13584 4576
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13464 4282 13584 4298
rect 13452 4276 13584 4282
rect 13504 4270 13584 4276
rect 13452 4218 13504 4224
rect 13648 4214 13676 4422
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13740 3670 13768 4014
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 12176 3097 12204 3130
rect 13268 3120 13320 3126
rect 12162 3088 12218 3097
rect 11704 3052 11756 3058
rect 13372 3097 13400 3130
rect 13268 3062 13320 3068
rect 13358 3088 13414 3097
rect 12162 3023 12218 3032
rect 13084 3052 13136 3058
rect 11704 2994 11756 3000
rect 13084 2994 13136 3000
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 11164 2746 11376 2774
rect 11164 2650 11192 2746
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10968 2304 11020 2310
rect 10796 2252 10968 2258
rect 10796 2246 11020 2252
rect 10796 2230 11008 2246
rect 11624 1902 11652 2858
rect 11716 2514 11744 2994
rect 13096 2961 13124 2994
rect 13082 2952 13138 2961
rect 13082 2887 13138 2896
rect 13280 2774 13308 3062
rect 13358 3023 13414 3032
rect 13280 2746 13400 2774
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 13268 2032 13320 2038
rect 13268 1974 13320 1980
rect 11612 1896 11664 1902
rect 11612 1838 11664 1844
rect 12256 1760 12308 1766
rect 12256 1702 12308 1708
rect 12268 800 12296 1702
rect 13280 1630 13308 1974
rect 13268 1624 13320 1630
rect 13268 1566 13320 1572
rect 13372 1578 13400 2746
rect 13464 2038 13492 3538
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13556 2689 13584 3402
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13648 2854 13676 3130
rect 13740 2990 13768 3402
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13832 2854 13860 4576
rect 14292 4128 14320 6326
rect 14476 5409 14504 10118
rect 14568 10118 14780 10146
rect 14568 6934 14596 10118
rect 14830 9752 14886 9761
rect 14830 9687 14886 9696
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14660 9178 14688 9590
rect 14844 9586 14872 9687
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14556 6928 14608 6934
rect 14556 6870 14608 6876
rect 14568 5642 14596 6870
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14462 5400 14518 5409
rect 14462 5335 14518 5344
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14292 4100 14412 4128
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14016 3534 14044 4014
rect 14384 3942 14412 4100
rect 14476 3942 14504 5034
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14016 2990 14044 3470
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13542 2680 13598 2689
rect 13542 2615 13598 2624
rect 14292 2514 14320 3470
rect 14476 3466 14504 3878
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 14384 2990 14412 3062
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14660 2650 14688 8910
rect 14936 7410 14964 11852
rect 15016 11834 15068 11840
rect 15120 11354 15148 12718
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15120 10266 15148 10610
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15028 8634 15056 9454
rect 15212 9382 15240 12106
rect 15304 9518 15332 12922
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15396 8974 15424 13466
rect 15488 9110 15516 16918
rect 15568 16516 15620 16522
rect 15672 16504 15700 18702
rect 16040 17746 16068 30194
rect 16764 29572 16816 29578
rect 16764 29514 16816 29520
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 16132 23866 16160 24142
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16224 21962 16252 22374
rect 16776 22098 16804 29514
rect 17132 24744 17184 24750
rect 17132 24686 17184 24692
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16960 23730 16988 24142
rect 17144 23798 17172 24686
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17236 23798 17264 24006
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 17224 23792 17276 23798
rect 17224 23734 17276 23740
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 17420 23662 17448 30670
rect 17604 29850 17632 35022
rect 19444 34746 19472 37198
rect 20640 37182 20760 37198
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 21732 37120 21784 37126
rect 21732 37062 21784 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19984 35080 20036 35086
rect 19984 35022 20036 35028
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19432 34740 19484 34746
rect 19432 34682 19484 34688
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 18420 31952 18472 31958
rect 18420 31894 18472 31900
rect 17592 29844 17644 29850
rect 17592 29786 17644 29792
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 17420 23254 17448 23598
rect 17408 23248 17460 23254
rect 17408 23190 17460 23196
rect 17512 23050 17540 24006
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17604 22710 17632 29582
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 17592 22704 17644 22710
rect 17592 22646 17644 22652
rect 17604 22506 17632 22646
rect 17592 22500 17644 22506
rect 17592 22442 17644 22448
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 16120 21956 16172 21962
rect 16120 21898 16172 21904
rect 16212 21956 16264 21962
rect 16212 21898 16264 21904
rect 16132 21146 16160 21898
rect 17696 21622 17724 21966
rect 17684 21616 17736 21622
rect 17684 21558 17736 21564
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16132 20058 16160 21082
rect 16856 20936 16908 20942
rect 16960 20924 16988 21422
rect 17040 21412 17092 21418
rect 17040 21354 17092 21360
rect 16908 20896 16988 20924
rect 16856 20878 16908 20884
rect 16960 20534 16988 20896
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16120 17808 16172 17814
rect 16304 17808 16356 17814
rect 16172 17768 16304 17796
rect 16120 17750 16172 17756
rect 16304 17750 16356 17756
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16040 16726 16068 17682
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16500 17338 16528 17614
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 15752 16516 15804 16522
rect 15672 16476 15752 16504
rect 15568 16458 15620 16464
rect 15752 16458 15804 16464
rect 15580 15706 15608 16458
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15672 15026 15700 16050
rect 16592 15586 16620 20198
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16684 19514 16712 19722
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16776 19378 16804 19654
rect 16868 19514 16896 19654
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16960 18850 16988 20470
rect 17052 20398 17080 21354
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17144 20466 17172 21286
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17040 20392 17092 20398
rect 17040 20334 17092 20340
rect 17224 20324 17276 20330
rect 17224 20266 17276 20272
rect 17236 19786 17264 20266
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17144 18970 17172 19314
rect 17328 18970 17356 21490
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17880 21078 17908 21286
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 17500 20324 17552 20330
rect 17500 20266 17552 20272
rect 17512 19514 17540 20266
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 16960 18822 17172 18850
rect 17144 18766 17172 18822
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16960 17882 16988 18158
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16776 16794 16804 17138
rect 16868 16998 16896 17546
rect 16960 17338 16988 17818
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16764 16516 16816 16522
rect 16764 16458 16816 16464
rect 16670 16008 16726 16017
rect 16670 15943 16672 15952
rect 16724 15943 16726 15952
rect 16672 15914 16724 15920
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16316 15558 16620 15586
rect 16224 15162 16252 15506
rect 16316 15502 16344 15558
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 15660 13456 15712 13462
rect 15660 13398 15712 13404
rect 15672 13326 15700 13398
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15750 12880 15806 12889
rect 15750 12815 15752 12824
rect 15804 12815 15806 12824
rect 15752 12786 15804 12792
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11098 15608 12038
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15580 11070 15700 11098
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10266 15608 10950
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 15028 6662 15056 7822
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15014 5536 15070 5545
rect 15014 5471 15070 5480
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14752 4554 14780 5034
rect 15028 4622 15056 5471
rect 15212 5370 15240 7414
rect 15290 6896 15346 6905
rect 15290 6831 15346 6840
rect 15384 6860 15436 6866
rect 15304 6322 15332 6831
rect 15384 6802 15436 6808
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15304 6089 15332 6122
rect 15290 6080 15346 6089
rect 15290 6015 15346 6024
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15396 4758 15424 6802
rect 15488 5234 15516 8910
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 15488 4486 15516 4966
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 14832 3460 14884 3466
rect 14884 3420 15240 3448
rect 14832 3402 14884 3408
rect 15212 2961 15240 3420
rect 15198 2952 15254 2961
rect 15198 2887 15254 2896
rect 15580 2774 15608 10202
rect 15672 7818 15700 11070
rect 15764 10810 15792 11630
rect 15856 11218 15884 13262
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15948 11286 15976 12922
rect 16316 12866 16344 14962
rect 16408 13802 16436 15098
rect 16500 14482 16528 15438
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 16592 14482 16620 14826
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16500 12986 16528 13806
rect 16592 13734 16620 14282
rect 16684 13938 16712 15438
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16316 12838 16528 12866
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 12322 16160 12718
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16302 12336 16358 12345
rect 16132 12294 16302 12322
rect 16302 12271 16304 12280
rect 16356 12271 16358 12280
rect 16304 12242 16356 12248
rect 16120 12232 16172 12238
rect 16408 12186 16436 12582
rect 16120 12174 16172 12180
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 16040 10674 16068 11086
rect 16132 10810 16160 12174
rect 16316 12158 16436 12186
rect 16316 12102 16344 12158
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16500 11354 16528 12838
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16684 12374 16712 12718
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16592 12170 16620 12242
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16592 11898 16620 12106
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 15844 10464 15896 10470
rect 16316 10441 16344 11290
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 15844 10406 15896 10412
rect 16302 10432 16358 10441
rect 15856 10180 15884 10406
rect 16302 10367 16358 10376
rect 15936 10192 15988 10198
rect 15856 10152 15936 10180
rect 15936 10134 15988 10140
rect 16212 10192 16264 10198
rect 16264 10140 16344 10146
rect 16212 10134 16344 10140
rect 16224 10118 16344 10134
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15764 8430 15792 9114
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15672 3942 15700 5170
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15304 2746 15608 2774
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 14476 2106 14504 2314
rect 14464 2100 14516 2106
rect 14464 2042 14516 2048
rect 13452 2032 13504 2038
rect 13452 1974 13504 1980
rect 13372 1550 13584 1578
rect 13556 800 13584 1550
rect 14568 1426 14596 2314
rect 15304 2310 15332 2746
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15580 2310 15608 2450
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15672 1698 15700 3878
rect 15750 2952 15806 2961
rect 15856 2922 15884 7346
rect 16040 6118 16068 8298
rect 16132 8294 16160 9862
rect 16316 9674 16344 10118
rect 16408 9738 16436 10610
rect 16500 10130 16528 11086
rect 16684 10266 16712 11086
rect 16776 11014 16804 16458
rect 16868 14618 16896 16526
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16960 15502 16988 15982
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16960 14498 16988 15438
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16868 14470 16988 14498
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16868 10742 16896 14470
rect 17052 13394 17080 15302
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 17052 12782 17080 12854
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17144 10985 17172 18702
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17236 16980 17264 17138
rect 17316 16992 17368 16998
rect 17236 16969 17316 16980
rect 17222 16960 17316 16969
rect 17278 16952 17316 16960
rect 17316 16934 17368 16940
rect 17222 16895 17278 16904
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17236 15706 17264 15846
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17236 14958 17264 15642
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17236 11898 17264 13262
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17224 11008 17276 11014
rect 17130 10976 17186 10985
rect 17224 10950 17276 10956
rect 17130 10911 17186 10920
rect 16946 10840 17002 10849
rect 16946 10775 17002 10784
rect 16960 10742 16988 10775
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16868 10606 16896 10678
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 17236 10538 17264 10950
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 17236 10146 17264 10474
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 17052 10118 17264 10146
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 16486 9752 16542 9761
rect 16408 9710 16486 9738
rect 16486 9687 16542 9696
rect 16316 9646 16436 9674
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16224 7546 16252 8978
rect 16316 8809 16344 8978
rect 16302 8800 16358 8809
rect 16302 8735 16358 8744
rect 16408 8430 16436 9646
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16302 7984 16358 7993
rect 16302 7919 16304 7928
rect 16356 7919 16358 7928
rect 16396 7948 16448 7954
rect 16304 7890 16356 7896
rect 16396 7890 16448 7896
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 16040 5409 16068 5714
rect 16026 5400 16082 5409
rect 16026 5335 16082 5344
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 4826 15976 4966
rect 16132 4826 16160 5170
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16224 4622 16252 6938
rect 16302 6760 16358 6769
rect 16302 6695 16358 6704
rect 16316 6322 16344 6695
rect 16408 6458 16436 7890
rect 16500 7274 16528 9687
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16316 5710 16344 6258
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16500 5778 16528 6190
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16592 5234 16620 7686
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16026 3768 16082 3777
rect 16026 3703 16082 3712
rect 16210 3768 16266 3777
rect 16210 3703 16266 3712
rect 16040 3670 16068 3703
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 15750 2887 15752 2896
rect 15804 2887 15806 2896
rect 15844 2916 15896 2922
rect 15752 2858 15804 2864
rect 15844 2858 15896 2864
rect 16040 2774 16068 3606
rect 16224 3097 16252 3703
rect 16210 3088 16266 3097
rect 16684 3058 16712 8774
rect 16776 7410 16804 9930
rect 17052 9518 17080 10118
rect 17132 9988 17184 9994
rect 17132 9930 17184 9936
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16868 7750 16896 9114
rect 17144 8090 17172 9930
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17236 9217 17264 9454
rect 17222 9208 17278 9217
rect 17420 9178 17448 16594
rect 17604 16590 17632 18226
rect 17880 17678 17908 18566
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17498 16008 17554 16017
rect 17498 15943 17500 15952
rect 17552 15943 17554 15952
rect 17500 15914 17552 15920
rect 17500 15088 17552 15094
rect 17500 15030 17552 15036
rect 17512 14657 17540 15030
rect 17880 15026 17908 16050
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17498 14648 17554 14657
rect 17498 14583 17554 14592
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17604 14414 17632 14554
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17696 14006 17724 14826
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17788 13530 17816 14214
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17788 13274 17816 13466
rect 17696 13246 17816 13274
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17498 9616 17554 9625
rect 17604 9586 17632 11494
rect 17696 11150 17724 13246
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17788 11762 17816 13126
rect 17880 12918 17908 14758
rect 17972 14634 18000 29106
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 18156 24410 18184 24686
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18064 23322 18092 24142
rect 18340 23866 18368 24142
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18236 22568 18288 22574
rect 18236 22510 18288 22516
rect 18156 22234 18184 22510
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18248 22098 18276 22510
rect 18236 22092 18288 22098
rect 18236 22034 18288 22040
rect 18432 20942 18460 31894
rect 18524 29306 18552 34546
rect 19064 34536 19116 34542
rect 19064 34478 19116 34484
rect 18788 32224 18840 32230
rect 18788 32166 18840 32172
rect 18512 29300 18564 29306
rect 18512 29242 18564 29248
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18524 23633 18552 23666
rect 18510 23624 18566 23633
rect 18510 23559 18566 23568
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18524 22098 18552 22374
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18512 22092 18564 22098
rect 18512 22034 18564 22040
rect 18616 21690 18644 22170
rect 18708 21894 18736 22578
rect 18800 21962 18828 32166
rect 19076 24818 19104 34478
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19340 33652 19392 33658
rect 19340 33594 19392 33600
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 18788 21956 18840 21962
rect 18788 21898 18840 21904
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 18696 21480 18748 21486
rect 18696 21422 18748 21428
rect 18708 21146 18736 21422
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 18064 20602 18092 20810
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 18144 19780 18196 19786
rect 18144 19722 18196 19728
rect 18156 19514 18184 19722
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 18248 18766 18276 20878
rect 18800 19378 18828 21898
rect 19352 21010 19380 33594
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19996 29850 20024 35022
rect 20732 34610 20760 37062
rect 20720 34604 20772 34610
rect 20720 34546 20772 34552
rect 21744 33998 21772 37062
rect 22940 35290 22968 37198
rect 23860 37126 23888 39200
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 24688 35290 24716 37198
rect 25792 37126 25820 39200
rect 27080 37262 27108 39200
rect 27068 37256 27120 37262
rect 27068 37198 27120 37204
rect 27804 37256 27856 37262
rect 27804 37198 27856 37204
rect 25780 37120 25832 37126
rect 25780 37062 25832 37068
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 22928 35284 22980 35290
rect 22928 35226 22980 35232
rect 24676 35284 24728 35290
rect 24676 35226 24728 35232
rect 22008 35080 22060 35086
rect 22008 35022 22060 35028
rect 21732 33992 21784 33998
rect 21732 33934 21784 33940
rect 21824 33856 21876 33862
rect 21824 33798 21876 33804
rect 20168 32428 20220 32434
rect 20168 32370 20220 32376
rect 20180 31754 20208 32370
rect 20180 31726 20392 31754
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19444 23662 19472 24550
rect 19996 24274 20024 24686
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19444 23322 19472 23598
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19812 22166 19840 22578
rect 19800 22160 19852 22166
rect 19800 22102 19852 22108
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19444 21554 19472 21830
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19800 21412 19852 21418
rect 19800 21354 19852 21360
rect 19812 21146 19840 21354
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18892 20602 18920 20878
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 19352 19854 19380 20810
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20398 20024 21422
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20088 19446 20116 19654
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 17972 14606 18092 14634
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17972 11898 18000 14418
rect 18064 14414 18092 14606
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18052 12844 18104 12850
rect 18156 12832 18184 18022
rect 18248 17882 18276 18702
rect 18984 18426 19012 19246
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 19076 17882 19104 18158
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 14074 18276 17478
rect 19444 17338 19472 19314
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18420 14952 18472 14958
rect 18418 14920 18420 14929
rect 18472 14920 18474 14929
rect 18418 14855 18474 14864
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18248 13462 18276 14010
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18104 12804 18184 12832
rect 18052 12786 18104 12792
rect 18248 12306 18276 13262
rect 18340 12442 18368 13262
rect 18432 12986 18460 13806
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 18432 11354 18460 12174
rect 18524 12170 18552 16594
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 18616 13530 18644 14282
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17682 9888 17738 9897
rect 17682 9823 17738 9832
rect 17498 9551 17554 9560
rect 17592 9580 17644 9586
rect 17222 9143 17278 9152
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17328 8566 17356 8774
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17420 8090 17448 8502
rect 17512 8090 17540 9551
rect 17592 9522 17644 9528
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 17590 7848 17646 7857
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16960 7546 16988 7822
rect 17500 7812 17552 7818
rect 17696 7818 17724 9823
rect 17590 7783 17646 7792
rect 17684 7812 17736 7818
rect 17500 7754 17552 7760
rect 17314 7712 17370 7721
rect 17314 7647 17370 7656
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 17052 7342 17080 7482
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 16948 7268 17000 7274
rect 16948 7210 17000 7216
rect 16960 6798 16988 7210
rect 17130 7168 17186 7177
rect 17130 7103 17186 7112
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16868 6474 16896 6734
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17052 6474 17080 6598
rect 16868 6446 17080 6474
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 17052 5370 17080 6326
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16210 3023 16266 3032
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 15856 2746 16068 2774
rect 15856 2281 15884 2746
rect 16776 2650 16804 4558
rect 16960 4321 16988 4558
rect 16946 4312 17002 4321
rect 16946 4247 17002 4256
rect 17144 4214 17172 7103
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17236 5778 17264 6190
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17236 5545 17264 5714
rect 17222 5536 17278 5545
rect 17222 5471 17278 5480
rect 17328 5370 17356 7647
rect 17512 7002 17540 7754
rect 17604 7750 17632 7783
rect 17684 7754 17736 7760
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17682 7304 17738 7313
rect 17592 7268 17644 7274
rect 17682 7239 17738 7248
rect 17592 7210 17644 7216
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17406 5808 17462 5817
rect 17406 5743 17462 5752
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16868 3670 16896 3946
rect 17420 3738 17448 5743
rect 17604 5681 17632 7210
rect 17696 6322 17724 7239
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17590 5672 17646 5681
rect 17590 5607 17646 5616
rect 17498 4856 17554 4865
rect 17498 4791 17500 4800
rect 17552 4791 17554 4800
rect 17500 4762 17552 4768
rect 17788 4162 17816 11018
rect 18524 10062 18552 11086
rect 18616 10810 18644 13466
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18708 11762 18736 12650
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18616 10266 18644 10542
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18512 10056 18564 10062
rect 18510 10024 18512 10033
rect 18564 10024 18566 10033
rect 18510 9959 18566 9968
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18064 9178 18092 9590
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17866 8664 17922 8673
rect 17866 8599 17922 8608
rect 17880 7834 17908 8599
rect 17972 8129 18000 8774
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 18064 8265 18092 8298
rect 18050 8256 18106 8265
rect 18050 8191 18106 8200
rect 17958 8120 18014 8129
rect 17958 8055 18014 8064
rect 17880 7806 18184 7834
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17880 7206 17908 7346
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17880 6798 17908 7142
rect 18050 7032 18106 7041
rect 18050 6967 18106 6976
rect 18064 6798 18092 6967
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17868 5296 17920 5302
rect 17868 5238 17920 5244
rect 17696 4146 17816 4162
rect 17684 4140 17816 4146
rect 17736 4134 17816 4140
rect 17684 4082 17736 4088
rect 17880 4078 17908 5238
rect 17972 4622 18000 5646
rect 18064 5166 18092 6054
rect 18156 5352 18184 7806
rect 18248 7546 18276 8570
rect 18340 8022 18368 9658
rect 18512 8560 18564 8566
rect 18510 8528 18512 8537
rect 18564 8528 18566 8537
rect 18420 8492 18472 8498
rect 18510 8463 18566 8472
rect 18420 8434 18472 8440
rect 18328 8016 18380 8022
rect 18328 7958 18380 7964
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18340 7478 18368 7686
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 18432 5710 18460 8434
rect 18708 8412 18736 11698
rect 18800 10198 18828 12718
rect 18984 12345 19012 17138
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19352 16590 19380 17070
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19444 16454 19472 17070
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 19628 15570 19656 15914
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19352 14414 19380 15098
rect 19996 15042 20024 17274
rect 20088 17270 20116 19246
rect 20272 18902 20300 20198
rect 20260 18896 20312 18902
rect 20260 18838 20312 18844
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19904 15014 20024 15042
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19444 14414 19472 14826
rect 19904 14482 19932 15014
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19352 12986 19380 14214
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 18970 12336 19026 12345
rect 18970 12271 19026 12280
rect 19062 12200 19118 12209
rect 19062 12135 19118 12144
rect 18788 10192 18840 10198
rect 18788 10134 18840 10140
rect 19076 9722 19104 12135
rect 19352 11354 19380 12718
rect 19444 12442 19472 14214
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14074 20024 14894
rect 20088 14618 20116 16390
rect 20180 14890 20208 18770
rect 20272 18204 20300 18838
rect 20364 18306 20392 31726
rect 20444 31136 20496 31142
rect 20444 31078 20496 31084
rect 20456 22642 20484 31078
rect 20628 29640 20680 29646
rect 20628 29582 20680 29588
rect 20640 24274 20668 29582
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20640 23798 20668 24210
rect 20628 23792 20680 23798
rect 20628 23734 20680 23740
rect 20732 23186 20760 27270
rect 21088 23248 21140 23254
rect 21088 23190 21140 23196
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20916 22778 20944 23054
rect 21100 22778 21128 23190
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21192 22778 21220 22986
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20456 21486 20484 22578
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20640 22234 20668 22510
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 20456 18902 20484 19178
rect 20444 18896 20496 18902
rect 20444 18838 20496 18844
rect 20640 18698 20668 20742
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20364 18278 20668 18306
rect 20272 18176 20484 18204
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20260 17264 20312 17270
rect 20260 17206 20312 17212
rect 20272 15366 20300 17206
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19996 13530 20024 13874
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 20088 13462 20116 14418
rect 20076 13456 20128 13462
rect 20128 13416 20208 13444
rect 20076 13398 20128 13404
rect 19984 13252 20036 13258
rect 20036 13212 20116 13240
rect 19984 13194 20036 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19996 12238 20024 12582
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20088 11898 20116 13212
rect 20180 12442 20208 13416
rect 20272 12986 20300 14962
rect 20364 13394 20392 18022
rect 20456 17660 20484 18176
rect 20456 17632 20576 17660
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20456 16726 20484 17478
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20456 15162 20484 15846
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20456 12866 20484 13806
rect 20272 12838 20484 12866
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18524 8384 18736 8412
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18156 5324 18276 5352
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18156 4690 18184 5170
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17592 4072 17644 4078
rect 17590 4040 17592 4049
rect 17868 4072 17920 4078
rect 17644 4040 17646 4049
rect 17868 4014 17920 4020
rect 17590 3975 17646 3984
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 18248 3602 18276 5324
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18326 4448 18382 4457
rect 18326 4383 18382 4392
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 16868 3369 16896 3470
rect 16854 3360 16910 3369
rect 16854 3295 16910 3304
rect 17880 3058 17908 3470
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17972 3126 18000 3334
rect 18340 3194 18368 4383
rect 18432 4146 18460 4558
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18432 3534 18460 4082
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 15842 2272 15898 2281
rect 15842 2207 15898 2216
rect 15660 1692 15712 1698
rect 15660 1634 15712 1640
rect 16132 1426 16160 2314
rect 14556 1420 14608 1426
rect 14556 1362 14608 1368
rect 15476 1420 15528 1426
rect 15476 1362 15528 1368
rect 16120 1420 16172 1426
rect 16120 1362 16172 1368
rect 15488 800 15516 1362
rect 16776 800 16804 2382
rect 17236 2106 17264 2518
rect 18524 2310 18552 8384
rect 18602 7576 18658 7585
rect 18602 7511 18658 7520
rect 18616 7478 18644 7511
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18616 5846 18644 6734
rect 18694 6488 18750 6497
rect 18694 6423 18696 6432
rect 18748 6423 18750 6432
rect 18696 6394 18748 6400
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 18800 4622 18828 9318
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18892 7546 18920 8230
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 19168 6254 19196 10474
rect 19352 10130 19380 11154
rect 19444 10810 19472 11698
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19536 11218 19564 11494
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19982 11112 20038 11121
rect 19982 11047 20038 11056
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19246 7440 19302 7449
rect 19246 7375 19302 7384
rect 19260 6458 19288 7375
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19248 6452 19300 6458
rect 19352 6440 19380 7278
rect 19444 6934 19472 8026
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19432 6928 19484 6934
rect 19432 6870 19484 6876
rect 19904 6644 19932 7346
rect 19996 6798 20024 11047
rect 20180 10810 20208 11630
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20272 10198 20300 12838
rect 20352 12368 20404 12374
rect 20352 12310 20404 12316
rect 20364 11626 20392 12310
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20456 11558 20484 12038
rect 20548 11762 20576 17632
rect 20640 16182 20668 18278
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20732 17882 20760 18158
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20824 17338 20852 20470
rect 20916 19514 20944 21286
rect 21560 19854 21588 22714
rect 21836 20602 21864 33798
rect 22020 29850 22048 35022
rect 23204 33992 23256 33998
rect 23204 33934 23256 33940
rect 22008 29844 22060 29850
rect 22008 29786 22060 29792
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22572 21010 22600 21422
rect 23216 21010 23244 33934
rect 27172 32434 27200 37062
rect 27816 34746 27844 37198
rect 29012 37126 29040 39200
rect 30300 37210 30328 39200
rect 30380 37256 30432 37262
rect 30300 37204 30380 37210
rect 30300 37198 30432 37204
rect 31588 37210 31616 39200
rect 33520 37262 33548 39200
rect 34808 37262 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 36740 37262 36768 39200
rect 31760 37256 31812 37262
rect 31588 37204 31760 37210
rect 31588 37198 31812 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 36728 37256 36780 37262
rect 36728 37198 36780 37204
rect 30300 37182 30420 37198
rect 31588 37182 31800 37198
rect 31852 37188 31904 37194
rect 31852 37130 31904 37136
rect 35532 37188 35584 37194
rect 35532 37130 35584 37136
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 30012 37120 30064 37126
rect 30012 37062 30064 37068
rect 29736 36916 29788 36922
rect 29736 36858 29788 36864
rect 27804 34740 27856 34746
rect 27804 34682 27856 34688
rect 27344 34604 27396 34610
rect 27344 34546 27396 34552
rect 27356 34202 27384 34546
rect 27344 34196 27396 34202
rect 27344 34138 27396 34144
rect 29748 33998 29776 36858
rect 29736 33992 29788 33998
rect 29736 33934 29788 33940
rect 29828 33856 29880 33862
rect 29828 33798 29880 33804
rect 29840 33658 29868 33798
rect 29828 33652 29880 33658
rect 29828 33594 29880 33600
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 29000 32360 29052 32366
rect 29000 32302 29052 32308
rect 29012 31890 29040 32302
rect 29000 31884 29052 31890
rect 29000 31826 29052 31832
rect 29828 31884 29880 31890
rect 29828 31826 29880 31832
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 23204 21004 23256 21010
rect 23204 20946 23256 20952
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22388 20602 22416 20878
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 21824 20392 21876 20398
rect 21824 20334 21876 20340
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20916 16726 20944 19450
rect 21364 19440 21416 19446
rect 21364 19382 21416 19388
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21192 18834 21220 19110
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21192 18426 21220 18566
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 20916 16538 20944 16662
rect 20916 16510 21036 16538
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20640 15366 20668 16118
rect 20916 16114 20944 16390
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20812 16040 20864 16046
rect 20812 15982 20864 15988
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20732 14414 20760 15030
rect 20824 14618 20852 15982
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 21008 14482 21036 16510
rect 21192 16250 21220 17682
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21284 15162 21312 16594
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20640 12730 20668 13330
rect 20732 13326 20760 14350
rect 21376 13705 21404 19382
rect 21560 18290 21588 19790
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21652 17882 21680 18022
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21744 17678 21772 19314
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21744 16182 21772 17614
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21468 14890 21496 15574
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21362 13696 21418 13705
rect 21362 13631 21418 13640
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20640 12702 20760 12730
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20640 12374 20668 12582
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20732 11694 20760 12702
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20720 11688 20772 11694
rect 20534 11656 20590 11665
rect 20720 11630 20772 11636
rect 20534 11591 20590 11600
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 20364 10062 20392 10610
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20088 8498 20116 8978
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20088 7410 20116 8434
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19904 6616 20024 6644
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19352 6412 19564 6440
rect 19248 6394 19300 6400
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19352 5794 19380 6258
rect 19430 6080 19486 6089
rect 19430 6015 19486 6024
rect 19444 5914 19472 6015
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19352 5766 19472 5794
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 19076 4554 19104 5170
rect 19352 5166 19380 5646
rect 19444 5574 19472 5766
rect 19536 5710 19564 6412
rect 19996 6322 20024 6616
rect 20076 6384 20128 6390
rect 20074 6352 20076 6361
rect 20128 6352 20130 6361
rect 19984 6316 20036 6322
rect 20074 6287 20130 6296
rect 19984 6258 20036 6264
rect 19996 5710 20024 6258
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19984 5704 20036 5710
rect 20168 5704 20220 5710
rect 20036 5664 20116 5692
rect 19984 5646 20036 5652
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19352 5001 19380 5102
rect 19338 4992 19394 5001
rect 19338 4927 19394 4936
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 19076 4146 19104 4490
rect 19444 4486 19472 5510
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19524 5296 19576 5302
rect 19522 5264 19524 5273
rect 19576 5264 19578 5273
rect 19522 5199 19578 5208
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19628 4486 19656 5170
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19444 4214 19472 4422
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19522 4176 19578 4185
rect 19064 4140 19116 4146
rect 19522 4111 19578 4120
rect 19064 4082 19116 4088
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18616 2446 18644 2858
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 17224 2100 17276 2106
rect 17224 2042 17276 2048
rect 18708 800 18736 2246
rect 18800 1766 18828 2382
rect 18788 1760 18840 1766
rect 18788 1702 18840 1708
rect 18892 1290 18920 2790
rect 18984 2514 19012 2790
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 18880 1284 18932 1290
rect 18880 1226 18932 1232
rect 19168 1086 19196 3878
rect 19260 3738 19288 3878
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19352 3534 19380 4014
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19352 3058 19380 3470
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19352 1834 19380 2586
rect 19444 2514 19472 3946
rect 19536 3738 19564 4111
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19812 3670 19840 4014
rect 19800 3664 19852 3670
rect 19800 3606 19852 3612
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19996 2394 20024 5510
rect 20088 5370 20116 5664
rect 20168 5646 20220 5652
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 20076 5228 20128 5234
rect 20180 5216 20208 5646
rect 20128 5188 20208 5216
rect 20076 5170 20128 5176
rect 20088 4622 20116 5170
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 20088 3913 20116 4422
rect 20074 3904 20130 3913
rect 20074 3839 20130 3848
rect 20088 3534 20116 3839
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 20088 2530 20116 3334
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 20180 2650 20208 2790
rect 20272 2650 20300 9998
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20364 4826 20392 8774
rect 20456 7426 20484 10678
rect 20548 7818 20576 11591
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20732 11014 20760 11494
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20824 10810 20852 11086
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20916 10146 20944 11698
rect 21008 10810 21036 12854
rect 21560 12238 21588 16050
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21652 13530 21680 14350
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21192 11830 21220 12038
rect 21180 11824 21232 11830
rect 21086 11792 21142 11801
rect 21180 11766 21232 11772
rect 21560 11762 21588 12174
rect 21086 11727 21142 11736
rect 21548 11756 21600 11762
rect 21100 11098 21128 11727
rect 21548 11698 21600 11704
rect 21100 11070 21220 11098
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21100 10674 21128 10950
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21008 10266 21036 10610
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 20916 10118 21036 10146
rect 20810 9480 20866 9489
rect 20810 9415 20866 9424
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 7886 20668 8230
rect 20732 8090 20760 8366
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20824 7886 20852 9415
rect 21008 8974 21036 10118
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 20902 8392 20958 8401
rect 20902 8327 20958 8336
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20456 7398 20852 7426
rect 20444 6928 20496 6934
rect 20444 6870 20496 6876
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20456 4690 20484 6870
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20640 5710 20668 6258
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20732 5234 20760 6666
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20088 2502 20300 2530
rect 19996 2366 20116 2394
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19444 2145 19472 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19430 2136 19486 2145
rect 19574 2139 19882 2148
rect 19430 2071 19486 2080
rect 19340 1828 19392 1834
rect 19340 1770 19392 1776
rect 19156 1080 19208 1086
rect 19156 1022 19208 1028
rect 19996 800 20024 2246
rect 20088 1358 20116 2366
rect 20076 1352 20128 1358
rect 20076 1294 20128 1300
rect 20272 1018 20300 2502
rect 20364 2038 20392 3334
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20352 2032 20404 2038
rect 20352 1974 20404 1980
rect 20456 1970 20484 2246
rect 20444 1964 20496 1970
rect 20444 1906 20496 1912
rect 20548 1494 20576 3878
rect 20536 1488 20588 1494
rect 20536 1430 20588 1436
rect 20640 1222 20668 4966
rect 20732 4146 20760 5170
rect 20824 4298 20852 7398
rect 20916 5914 20944 8327
rect 21008 7478 21036 8910
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21008 6866 21036 7142
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 21100 4826 21128 8298
rect 21192 5370 21220 11070
rect 21270 10704 21326 10713
rect 21270 10639 21326 10648
rect 21284 5914 21312 10639
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21468 6254 21496 6598
rect 21456 6248 21508 6254
rect 21362 6216 21418 6225
rect 21456 6190 21508 6196
rect 21362 6151 21364 6160
rect 21416 6151 21418 6160
rect 21364 6122 21416 6128
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21560 4826 21588 9658
rect 21652 6458 21680 13126
rect 21744 12918 21772 13262
rect 21732 12912 21784 12918
rect 21732 12854 21784 12860
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21744 11898 21772 12174
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21836 9178 21864 20334
rect 22020 19446 22048 20334
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22848 20058 22876 20198
rect 22836 20052 22888 20058
rect 22888 20012 22968 20040
rect 22836 19994 22888 20000
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22836 19780 22888 19786
rect 22836 19722 22888 19728
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22664 17882 22692 18158
rect 22756 18086 22784 19722
rect 22848 19514 22876 19722
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22940 19446 22968 20012
rect 23216 19922 23244 20946
rect 24584 20392 24636 20398
rect 24584 20334 24636 20340
rect 24596 20058 24624 20334
rect 24584 20052 24636 20058
rect 24584 19994 24636 20000
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 22928 19440 22980 19446
rect 22928 19382 22980 19388
rect 23664 19304 23716 19310
rect 23570 19272 23626 19281
rect 23664 19246 23716 19252
rect 23570 19207 23626 19216
rect 23020 18692 23072 18698
rect 23020 18634 23072 18640
rect 23112 18692 23164 18698
rect 23112 18634 23164 18640
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22756 17814 22784 18022
rect 22744 17808 22796 17814
rect 22744 17750 22796 17756
rect 22284 17740 22336 17746
rect 22284 17682 22336 17688
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 22020 16998 22048 17070
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 21824 9172 21876 9178
rect 21824 9114 21876 9120
rect 22020 8498 22048 16934
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22204 12986 22232 13806
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 22112 11898 22140 12854
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22204 9518 22232 12650
rect 22296 12646 22324 17682
rect 23032 17338 23060 18634
rect 23124 18426 23152 18634
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23584 18290 23612 19207
rect 23676 18834 23704 19246
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23860 18630 23888 19790
rect 24676 19372 24728 19378
rect 24676 19314 24728 19320
rect 24688 19281 24716 19314
rect 24674 19272 24730 19281
rect 24674 19207 24730 19216
rect 24780 18970 24808 19790
rect 24872 19718 24900 21966
rect 25240 20330 25268 31758
rect 29092 29164 29144 29170
rect 29092 29106 29144 29112
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 25228 20324 25280 20330
rect 25228 20266 25280 20272
rect 25412 19848 25464 19854
rect 25412 19790 25464 19796
rect 24860 19712 24912 19718
rect 24860 19654 24912 19660
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25240 19446 25268 19654
rect 25424 19514 25452 19790
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 25228 19440 25280 19446
rect 25228 19382 25280 19388
rect 28736 19242 28764 25230
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28724 19236 28776 19242
rect 28724 19178 28776 19184
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22848 16794 22876 17070
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 23032 16250 23060 17274
rect 23308 17241 23336 17614
rect 23294 17232 23350 17241
rect 23112 17196 23164 17202
rect 23860 17202 23888 18566
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24228 17746 24256 18022
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24412 17338 24440 18226
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 23294 17167 23296 17176
rect 23112 17138 23164 17144
rect 23348 17167 23350 17176
rect 23848 17196 23900 17202
rect 23296 17138 23348 17144
rect 23848 17138 23900 17144
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 23124 16250 23152 17138
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23492 16590 23520 16934
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23124 15570 23152 15846
rect 23676 15706 23704 16526
rect 23860 16114 23888 17138
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23664 15700 23716 15706
rect 23664 15642 23716 15648
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 22572 15094 22600 15506
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22940 15162 22968 15438
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 22560 15088 22612 15094
rect 22560 15030 22612 15036
rect 22572 14414 22600 15030
rect 23492 15026 23520 15302
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22664 14618 22692 14894
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 23860 14521 23888 16050
rect 24596 15434 24624 17138
rect 24584 15428 24636 15434
rect 24584 15370 24636 15376
rect 23846 14512 23902 14521
rect 23756 14476 23808 14482
rect 23846 14447 23902 14456
rect 23756 14418 23808 14424
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22388 13802 22416 14214
rect 22480 13938 22508 14214
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22572 13818 22600 14350
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 22376 13796 22428 13802
rect 22376 13738 22428 13744
rect 22480 13790 22600 13818
rect 22388 13462 22416 13738
rect 22376 13456 22428 13462
rect 22376 13398 22428 13404
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22480 10305 22508 13790
rect 22560 13252 22612 13258
rect 22560 13194 22612 13200
rect 22572 11898 22600 13194
rect 23216 12782 23244 13942
rect 23492 13394 23520 14350
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23768 13326 23796 14418
rect 28828 14074 28856 20878
rect 29104 17610 29132 29106
rect 29736 28552 29788 28558
rect 29736 28494 29788 28500
rect 29644 26376 29696 26382
rect 29644 26318 29696 26324
rect 29656 18154 29684 26318
rect 29748 19310 29776 28494
rect 29840 22778 29868 31826
rect 29932 28762 29960 32370
rect 30024 32366 30052 37062
rect 31864 35086 31892 37130
rect 32312 37120 32364 37126
rect 32312 37062 32364 37068
rect 33600 37120 33652 37126
rect 33600 37062 33652 37068
rect 31852 35080 31904 35086
rect 31852 35022 31904 35028
rect 30564 34944 30616 34950
rect 30564 34886 30616 34892
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30012 32360 30064 32366
rect 30012 32302 30064 32308
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 29920 28756 29972 28762
rect 29920 28698 29972 28704
rect 30024 26586 30052 30670
rect 30116 29306 30144 33934
rect 30104 29300 30156 29306
rect 30104 29242 30156 29248
rect 30012 26580 30064 26586
rect 30012 26522 30064 26528
rect 29828 22772 29880 22778
rect 29828 22714 29880 22720
rect 29736 19304 29788 19310
rect 29736 19246 29788 19252
rect 30576 18902 30604 34886
rect 32324 32026 32352 37062
rect 33612 36922 33640 37062
rect 33600 36916 33652 36922
rect 33600 36858 33652 36864
rect 35348 36712 35400 36718
rect 35348 36654 35400 36660
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34520 36032 34572 36038
rect 34520 35974 34572 35980
rect 34532 34610 34560 35974
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34520 34604 34572 34610
rect 34520 34546 34572 34552
rect 33324 34536 33376 34542
rect 33324 34478 33376 34484
rect 32312 32020 32364 32026
rect 32312 31962 32364 31968
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 32036 24812 32088 24818
rect 32036 24754 32088 24760
rect 31760 23724 31812 23730
rect 31760 23666 31812 23672
rect 31772 22098 31800 23666
rect 31760 22092 31812 22098
rect 31760 22034 31812 22040
rect 32048 21146 32076 24754
rect 32036 21140 32088 21146
rect 32036 21082 32088 21088
rect 30564 18896 30616 18902
rect 30564 18838 30616 18844
rect 29644 18148 29696 18154
rect 29644 18090 29696 18096
rect 29092 17604 29144 17610
rect 29092 17546 29144 17552
rect 31576 17536 31628 17542
rect 31576 17478 31628 17484
rect 31588 17270 31616 17478
rect 31576 17264 31628 17270
rect 31576 17206 31628 17212
rect 32416 15638 32444 27814
rect 33140 18624 33192 18630
rect 33140 18566 33192 18572
rect 32404 15632 32456 15638
rect 32404 15574 32456 15580
rect 33152 15570 33180 18566
rect 33336 18222 33364 34478
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35360 34202 35388 36654
rect 35440 35080 35492 35086
rect 35440 35022 35492 35028
rect 35348 34196 35400 34202
rect 35348 34138 35400 34144
rect 35348 33516 35400 33522
rect 35348 33458 35400 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34152 30048 34204 30054
rect 34152 29990 34204 29996
rect 34164 27470 34192 29990
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29850 35388 33458
rect 35452 30938 35480 35022
rect 35544 32570 35572 37130
rect 35900 37120 35952 37126
rect 35900 37062 35952 37068
rect 35532 32564 35584 32570
rect 35532 32506 35584 32512
rect 35912 31822 35940 37062
rect 36728 36576 36780 36582
rect 36728 36518 36780 36524
rect 35900 31816 35952 31822
rect 35900 31758 35952 31764
rect 36740 31346 36768 36518
rect 38028 36174 38056 39200
rect 38290 38176 38346 38185
rect 38290 38111 38346 38120
rect 38200 37120 38252 37126
rect 38200 37062 38252 37068
rect 38212 36825 38240 37062
rect 38304 36922 38332 38111
rect 38292 36916 38344 36922
rect 38292 36858 38344 36864
rect 39316 36854 39344 39200
rect 39304 36848 39356 36854
rect 38198 36816 38254 36825
rect 39304 36790 39356 36796
rect 38198 36751 38254 36760
rect 38016 36168 38068 36174
rect 38016 36110 38068 36116
rect 38200 34944 38252 34950
rect 38200 34886 38252 34892
rect 38212 34785 38240 34886
rect 38198 34776 38254 34785
rect 38198 34711 38254 34720
rect 38198 33416 38254 33425
rect 38198 33351 38200 33360
rect 38252 33351 38254 33360
rect 38200 33322 38252 33328
rect 37004 31952 37056 31958
rect 37004 31894 37056 31900
rect 36728 31340 36780 31346
rect 36728 31282 36780 31288
rect 35440 30932 35492 30938
rect 35440 30874 35492 30880
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34152 27464 34204 27470
rect 34152 27406 34204 27412
rect 34716 25498 34744 29582
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 37016 28082 37044 31894
rect 38292 31816 38344 31822
rect 38292 31758 38344 31764
rect 38304 31385 38332 31758
rect 38290 31376 38346 31385
rect 38290 31311 38346 31320
rect 38292 30252 38344 30258
rect 38292 30194 38344 30200
rect 38304 30025 38332 30194
rect 38290 30016 38346 30025
rect 38290 29951 38346 29960
rect 38016 29164 38068 29170
rect 38016 29106 38068 29112
rect 37004 28076 37056 28082
rect 37004 28018 37056 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 26988 34848 26994
rect 34796 26930 34848 26936
rect 34704 25492 34756 25498
rect 34704 25434 34756 25440
rect 34612 25152 34664 25158
rect 34612 25094 34664 25100
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34532 21554 34560 23462
rect 34624 21554 34652 25094
rect 34808 23866 34836 26930
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 38028 24682 38056 29106
rect 38200 29028 38252 29034
rect 38200 28970 38252 28976
rect 38212 28665 38240 28970
rect 38198 28656 38254 28665
rect 38198 28591 38254 28600
rect 38200 26784 38252 26790
rect 38200 26726 38252 26732
rect 38212 26625 38240 26726
rect 38198 26616 38254 26625
rect 38198 26551 38254 26560
rect 38292 25288 38344 25294
rect 38290 25256 38292 25265
rect 38344 25256 38346 25265
rect 38290 25191 38346 25200
rect 38016 24676 38068 24682
rect 38016 24618 38068 24624
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 38304 23225 38332 23666
rect 38290 23216 38346 23225
rect 38290 23151 38346 23160
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38108 21888 38160 21894
rect 38304 21865 38332 21966
rect 38108 21830 38160 21836
rect 38290 21856 38346 21865
rect 34520 21548 34572 21554
rect 34520 21490 34572 21496
rect 34612 21548 34664 21554
rect 34612 21490 34664 21496
rect 34704 21344 34756 21350
rect 34704 21286 34756 21292
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 33324 18216 33376 18222
rect 33324 18158 33376 18164
rect 34532 17678 34560 18566
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 33232 17536 33284 17542
rect 33232 17478 33284 17484
rect 33244 16658 33272 17478
rect 33232 16652 33284 16658
rect 33232 16594 33284 16600
rect 33140 15564 33192 15570
rect 33140 15506 33192 15512
rect 31944 15496 31996 15502
rect 31944 15438 31996 15444
rect 31956 14618 31984 15438
rect 33416 14952 33468 14958
rect 33416 14894 33468 14900
rect 31944 14612 31996 14618
rect 31944 14554 31996 14560
rect 28816 14068 28868 14074
rect 28816 14010 28868 14016
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24412 13530 24440 13874
rect 33428 13530 33456 14894
rect 34244 13932 34296 13938
rect 34244 13874 34296 13880
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 33416 13524 33468 13530
rect 33416 13466 33468 13472
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23388 12912 23440 12918
rect 23388 12854 23440 12860
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 23400 12714 23428 12854
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23572 12640 23624 12646
rect 23572 12582 23624 12588
rect 23480 12368 23532 12374
rect 23480 12310 23532 12316
rect 22560 11892 22612 11898
rect 22560 11834 22612 11840
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22848 11150 22876 11698
rect 22836 11144 22888 11150
rect 22836 11086 22888 11092
rect 22466 10296 22522 10305
rect 22466 10231 22522 10240
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 22848 9081 22876 11086
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 22834 9072 22890 9081
rect 22834 9007 22890 9016
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22112 7342 22140 8298
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22204 7478 22232 7686
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22112 6866 22140 7278
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 22098 5944 22154 5953
rect 22098 5879 22100 5888
rect 22152 5879 22154 5888
rect 22100 5850 22152 5856
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 22098 5128 22154 5137
rect 22098 5063 22100 5072
rect 22152 5063 22154 5072
rect 22100 5034 22152 5040
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 21916 4752 21968 4758
rect 21916 4694 21968 4700
rect 20824 4270 20944 4298
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20732 1630 20760 2790
rect 20824 2689 20852 3946
rect 20916 3942 20944 4270
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 21454 3768 21510 3777
rect 21454 3703 21456 3712
rect 21508 3703 21510 3712
rect 21456 3674 21508 3680
rect 20810 2680 20866 2689
rect 20810 2615 20866 2624
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20824 1902 20852 2246
rect 20812 1896 20864 1902
rect 20812 1838 20864 1844
rect 20720 1624 20772 1630
rect 20720 1566 20772 1572
rect 20628 1216 20680 1222
rect 20628 1158 20680 1164
rect 20260 1012 20312 1018
rect 20260 954 20312 960
rect 21284 800 21312 2382
rect 21928 2378 21956 4694
rect 22204 4622 22232 5578
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22192 4616 22244 4622
rect 22098 4584 22154 4593
rect 22192 4558 22244 4564
rect 22098 4519 22100 4528
rect 22152 4519 22154 4528
rect 22100 4490 22152 4496
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22020 4146 22048 4422
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22098 3632 22154 3641
rect 22098 3567 22100 3576
rect 22152 3567 22154 3576
rect 22100 3538 22152 3544
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 22100 2848 22152 2854
rect 22098 2816 22100 2825
rect 22152 2816 22154 2825
rect 22098 2751 22154 2760
rect 22204 2417 22232 2858
rect 22190 2408 22246 2417
rect 21916 2372 21968 2378
rect 22190 2343 22246 2352
rect 21916 2314 21968 2320
rect 22296 1329 22324 3878
rect 22282 1320 22338 1329
rect 22282 1255 22338 1264
rect 22388 1154 22416 4966
rect 22480 3738 22508 7754
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 6798 22692 7686
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22664 4146 22692 5170
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 22756 4282 22784 4422
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 2582 22876 3334
rect 23124 3058 23152 4558
rect 23216 3738 23244 10746
rect 23492 10266 23520 12310
rect 23584 10674 23612 12582
rect 23768 11626 23796 12718
rect 24044 12306 24072 13330
rect 31392 12844 31444 12850
rect 31392 12786 31444 12792
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23664 11620 23716 11626
rect 23664 11562 23716 11568
rect 23756 11620 23808 11626
rect 23756 11562 23808 11568
rect 23676 10674 23704 11562
rect 23860 10810 23888 12038
rect 24136 11218 24164 12174
rect 24676 12164 24728 12170
rect 24676 12106 24728 12112
rect 24688 11898 24716 12106
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24228 11354 24256 11698
rect 24308 11620 24360 11626
rect 24308 11562 24360 11568
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 24320 11218 24348 11562
rect 24596 11354 24624 11766
rect 30380 11756 30432 11762
rect 30380 11698 30432 11704
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24308 11212 24360 11218
rect 24308 11154 24360 11160
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24780 10810 24808 11086
rect 30392 10810 30420 11698
rect 30840 11076 30892 11082
rect 30840 11018 30892 11024
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 30380 10804 30432 10810
rect 30380 10746 30432 10752
rect 30852 10674 30880 11018
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 30840 10668 30892 10674
rect 30840 10610 30892 10616
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23308 9722 23336 9998
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23308 7478 23336 7686
rect 23296 7472 23348 7478
rect 23296 7414 23348 7420
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23400 7002 23428 7414
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 23388 5772 23440 5778
rect 23388 5714 23440 5720
rect 23400 5302 23428 5714
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 23480 3528 23532 3534
rect 23478 3496 23480 3505
rect 23532 3496 23534 3505
rect 23478 3431 23534 3440
rect 23940 3188 23992 3194
rect 23940 3130 23992 3136
rect 23952 3097 23980 3130
rect 23938 3088 23994 3097
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23572 3052 23624 3058
rect 23938 3023 23994 3032
rect 23572 2994 23624 3000
rect 22836 2576 22888 2582
rect 22742 2544 22798 2553
rect 22836 2518 22888 2524
rect 22742 2479 22744 2488
rect 22796 2479 22798 2488
rect 22744 2450 22796 2456
rect 23124 2446 23152 2994
rect 23112 2440 23164 2446
rect 23112 2382 23164 2388
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 22376 1148 22428 1154
rect 22376 1090 22428 1096
rect 23216 800 23244 2246
rect 23584 1465 23612 2994
rect 24228 2650 24256 6258
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24596 2582 24624 6802
rect 24780 5710 24808 10474
rect 24872 8634 24900 10610
rect 29552 9988 29604 9994
rect 29552 9930 29604 9936
rect 28264 9444 28316 9450
rect 28264 9386 28316 9392
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 28276 8498 28304 9386
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 25688 5568 25740 5574
rect 25688 5510 25740 5516
rect 24584 2576 24636 2582
rect 24584 2518 24636 2524
rect 25700 2514 25728 5510
rect 26700 4140 26752 4146
rect 26700 4082 26752 4088
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 26620 3534 26648 4014
rect 26712 3738 26740 4082
rect 26700 3732 26752 3738
rect 26700 3674 26752 3680
rect 26608 3528 26660 3534
rect 26608 3470 26660 3476
rect 28460 2650 28488 8910
rect 29564 7546 29592 9930
rect 30012 8356 30064 8362
rect 30012 8298 30064 8304
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 29552 7336 29604 7342
rect 29552 7278 29604 7284
rect 29564 6322 29592 7278
rect 29552 6316 29604 6322
rect 29552 6258 29604 6264
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29656 5710 29684 6054
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 30024 5166 30052 8298
rect 30196 7880 30248 7886
rect 30196 7822 30248 7828
rect 30012 5160 30064 5166
rect 30012 5102 30064 5108
rect 28908 3936 28960 3942
rect 28908 3878 28960 3884
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 28920 2514 28948 3878
rect 30208 2650 30236 7822
rect 31208 6724 31260 6730
rect 31208 6666 31260 6672
rect 31220 5234 31248 6666
rect 31116 5228 31168 5234
rect 31116 5170 31168 5176
rect 31208 5228 31260 5234
rect 31208 5170 31260 5176
rect 31128 5098 31156 5170
rect 31116 5092 31168 5098
rect 31116 5034 31168 5040
rect 31404 3738 31432 12786
rect 34256 11898 34284 13874
rect 34716 13870 34744 21286
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 37004 19712 37056 19718
rect 37004 19654 37056 19660
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 37016 18766 37044 19654
rect 37004 18760 37056 18766
rect 37004 18702 37056 18708
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 38120 17746 38148 21830
rect 38290 21791 38346 21800
rect 38292 19848 38344 19854
rect 38290 19816 38292 19825
rect 38344 19816 38346 19825
rect 38290 19751 38346 19760
rect 38292 18760 38344 18766
rect 38292 18702 38344 18708
rect 38304 18465 38332 18702
rect 38290 18456 38346 18465
rect 38290 18391 38346 18400
rect 38108 17740 38160 17746
rect 38108 17682 38160 17688
rect 35900 17196 35952 17202
rect 35900 17138 35952 17144
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35912 15706 35940 17138
rect 38198 17096 38254 17105
rect 38198 17031 38200 17040
rect 38252 17031 38254 17040
rect 38200 17002 38252 17008
rect 38108 16108 38160 16114
rect 38108 16050 38160 16056
rect 38120 15706 38148 16050
rect 35900 15700 35952 15706
rect 35900 15642 35952 15648
rect 38108 15700 38160 15706
rect 38108 15642 38160 15648
rect 38292 15496 38344 15502
rect 38292 15438 38344 15444
rect 38304 15065 38332 15438
rect 38290 15056 38346 15065
rect 38290 14991 38346 15000
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34704 13864 34756 13870
rect 34704 13806 34756 13812
rect 38200 13728 38252 13734
rect 38198 13696 38200 13705
rect 38252 13696 38254 13705
rect 34934 13628 35242 13637
rect 38198 13631 38254 13640
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34612 13320 34664 13326
rect 34612 13262 34664 13268
rect 34624 11898 34652 13262
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 34244 11892 34296 11898
rect 34244 11834 34296 11840
rect 34612 11892 34664 11898
rect 34612 11834 34664 11840
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 36464 10674 36492 12038
rect 38292 11756 38344 11762
rect 38292 11698 38344 11704
rect 38304 11665 38332 11698
rect 38290 11656 38346 11665
rect 38290 11591 38346 11600
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 38016 10464 38068 10470
rect 38016 10406 38068 10412
rect 38200 10464 38252 10470
rect 38200 10406 38252 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 36912 10056 36964 10062
rect 36912 9998 36964 10004
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 33874 7984 33930 7993
rect 33874 7919 33930 7928
rect 33888 7546 33916 7919
rect 36924 7546 36952 9998
rect 38028 8974 38056 10406
rect 38212 10305 38240 10406
rect 38198 10296 38254 10305
rect 38198 10231 38254 10240
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 33876 7540 33928 7546
rect 33876 7482 33928 7488
rect 36912 7540 36964 7546
rect 36912 7482 36964 7488
rect 35716 7404 35768 7410
rect 35716 7346 35768 7352
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 34704 7336 34756 7342
rect 34704 7278 34756 7284
rect 33876 6792 33928 6798
rect 33876 6734 33928 6740
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 30196 2644 30248 2650
rect 30196 2586 30248 2592
rect 25688 2508 25740 2514
rect 25688 2450 25740 2456
rect 28908 2508 28960 2514
rect 28908 2450 28960 2456
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 23570 1456 23626 1465
rect 23570 1391 23626 1400
rect 24504 800 24532 2382
rect 26436 800 26464 2382
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27724 800 27752 2246
rect 29012 800 29040 2382
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 30944 800 30972 2246
rect 32232 800 32260 2382
rect 33888 2378 33916 6734
rect 34428 5092 34480 5098
rect 34428 5034 34480 5040
rect 34440 2582 34468 5034
rect 34716 2650 34744 7278
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35728 3194 35756 7346
rect 38304 6905 38332 7346
rect 38290 6896 38346 6905
rect 38290 6831 38346 6840
rect 38200 5568 38252 5574
rect 38198 5536 38200 5545
rect 38252 5536 38254 5545
rect 38198 5471 38254 5480
rect 35808 5024 35860 5030
rect 35808 4966 35860 4972
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 35716 3188 35768 3194
rect 35716 3130 35768 3136
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34704 2644 34756 2650
rect 34704 2586 34756 2592
rect 34428 2576 34480 2582
rect 34428 2518 34480 2524
rect 35624 2576 35676 2582
rect 35624 2518 35676 2524
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 33876 2372 33928 2378
rect 33876 2314 33928 2320
rect 34164 800 34192 2382
rect 35452 800 35480 2382
rect 35636 2378 35664 2518
rect 35820 2514 35848 4966
rect 38028 3058 38056 4966
rect 38292 3528 38344 3534
rect 38290 3496 38292 3505
rect 38344 3496 38346 3505
rect 38290 3431 38346 3440
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 38016 3052 38068 3058
rect 38016 2994 38068 3000
rect 35808 2508 35860 2514
rect 35808 2450 35860 2456
rect 35624 2372 35676 2378
rect 35624 2314 35676 2320
rect 18 200 74 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 7746 200 7802 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 12254 200 12310 800
rect 13542 200 13598 800
rect 15474 200 15530 800
rect 16762 200 16818 800
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 26422 200 26478 800
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 37292 105 37320 2994
rect 38200 2848 38252 2854
rect 38200 2790 38252 2796
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 37384 800 37412 2246
rect 38212 2145 38240 2790
rect 38660 2372 38712 2378
rect 38660 2314 38712 2320
rect 38198 2136 38254 2145
rect 38198 2071 38254 2080
rect 38672 800 38700 2314
rect 37370 200 37426 800
rect 38658 200 38714 800
rect 37278 96 37334 105
rect 37278 31 37334 40
<< via2 >>
rect 2778 39480 2834 39536
rect 3146 37440 3202 37496
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1766 36116 1768 36136
rect 1768 36116 1820 36136
rect 1820 36116 1822 36136
rect 1766 36080 1822 36116
rect 1766 34040 1822 34096
rect 1766 32680 1822 32736
rect 1766 30676 1768 30696
rect 1768 30676 1820 30696
rect 1820 30676 1822 30696
rect 1766 30640 1822 30676
rect 1766 29280 1822 29336
rect 1766 27920 1822 27976
rect 1766 25880 1822 25936
rect 1766 24556 1768 24576
rect 1768 24556 1820 24576
rect 1820 24556 1822 24576
rect 1766 24520 1822 24556
rect 1766 22480 1822 22536
rect 1766 21120 1822 21176
rect 2410 20304 2466 20360
rect 1766 19796 1768 19816
rect 1768 19796 1820 19816
rect 1820 19796 1822 19816
rect 1766 19760 1822 19796
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4066 29008 4122 29064
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 7470 36488 7526 36544
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 1766 17720 1822 17776
rect 1766 16396 1768 16416
rect 1768 16396 1820 16416
rect 1820 16396 1822 16416
rect 1766 16360 1822 16396
rect 1766 14320 1822 14376
rect 1766 12960 1822 13016
rect 1950 12688 2006 12744
rect 1858 9460 1860 9480
rect 1860 9460 1912 9480
rect 1912 9460 1914 9480
rect 1858 9424 1914 9460
rect 2686 16768 2742 16824
rect 2686 15408 2742 15464
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 3330 17060 3386 17096
rect 3330 17040 3332 17060
rect 3332 17040 3384 17060
rect 3384 17040 3386 17060
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 3238 15272 3294 15328
rect 2778 12144 2834 12200
rect 2686 11600 2742 11656
rect 2686 11056 2742 11112
rect 3054 12008 3110 12064
rect 3238 12144 3294 12200
rect 3606 11076 3662 11112
rect 3606 11056 3608 11076
rect 3608 11056 3660 11076
rect 3660 11056 3662 11076
rect 1766 5752 1822 5808
rect 1766 4800 1822 4856
rect 3054 9696 3110 9752
rect 3606 10920 3662 10976
rect 3330 9052 3332 9072
rect 3332 9052 3384 9072
rect 3384 9052 3386 9072
rect 3330 9016 3386 9052
rect 3330 8492 3386 8528
rect 3330 8472 3332 8492
rect 3332 8472 3384 8492
rect 3384 8472 3386 8492
rect 3054 6160 3110 6216
rect 3422 6296 3478 6352
rect 4434 15952 4490 16008
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4158 13232 4214 13288
rect 4434 13132 4436 13152
rect 4436 13132 4488 13152
rect 4488 13132 4490 13152
rect 4434 13096 4490 13132
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4066 12164 4122 12200
rect 4066 12144 4068 12164
rect 4068 12144 4120 12164
rect 4120 12144 4122 12164
rect 4066 11772 4068 11792
rect 4068 11772 4120 11792
rect 4120 11772 4122 11792
rect 4066 11736 4122 11772
rect 4250 11872 4306 11928
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4526 10104 4582 10160
rect 3882 9560 3938 9616
rect 3698 8236 3700 8256
rect 3700 8236 3752 8256
rect 3752 8236 3754 8256
rect 3698 8200 3754 8236
rect 3882 7928 3938 7984
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4526 9016 4582 9072
rect 4894 11600 4950 11656
rect 5446 13232 5502 13288
rect 5262 12960 5318 13016
rect 5262 12552 5318 12608
rect 4802 9424 4858 9480
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3514 6160 3570 6216
rect 4618 7112 4674 7168
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4066 6432 4122 6488
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4158 5752 4214 5808
rect 1950 2216 2006 2272
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4618 3576 4674 3632
rect 4158 3304 4214 3360
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5446 12280 5502 12336
rect 5446 10684 5448 10704
rect 5448 10684 5500 10704
rect 5500 10684 5502 10704
rect 5446 10648 5502 10684
rect 5078 4936 5134 4992
rect 5170 1264 5226 1320
rect 5814 11600 5870 11656
rect 5998 10376 6054 10432
rect 5722 9172 5778 9208
rect 5722 9152 5724 9172
rect 5724 9152 5776 9172
rect 5776 9152 5778 9172
rect 5354 5208 5410 5264
rect 5630 4256 5686 4312
rect 6274 11872 6330 11928
rect 6182 11464 6238 11520
rect 6274 8744 6330 8800
rect 6642 11872 6698 11928
rect 7562 13096 7618 13152
rect 6458 9832 6514 9888
rect 6458 7948 6514 7984
rect 6458 7928 6460 7948
rect 6460 7928 6512 7948
rect 6512 7928 6514 7948
rect 6458 4548 6514 4584
rect 6458 4528 6460 4548
rect 6460 4528 6512 4548
rect 6512 4528 6514 4548
rect 6274 4120 6330 4176
rect 5906 3984 5962 4040
rect 6918 5344 6974 5400
rect 7378 12688 7434 12744
rect 7286 8064 7342 8120
rect 7286 7268 7342 7304
rect 7286 7248 7288 7268
rect 7288 7248 7340 7268
rect 7340 7248 7342 7268
rect 6826 3304 6882 3360
rect 6826 2372 6882 2408
rect 6826 2352 6828 2372
rect 6828 2352 6880 2372
rect 6880 2352 6882 2372
rect 8206 15136 8262 15192
rect 7838 10240 7894 10296
rect 7654 6840 7710 6896
rect 7654 3848 7710 3904
rect 7654 2796 7656 2816
rect 7656 2796 7708 2816
rect 7708 2796 7710 2816
rect 7654 2760 7710 2796
rect 8114 11464 8170 11520
rect 8206 9596 8208 9616
rect 8208 9596 8260 9616
rect 8260 9596 8262 9616
rect 8206 9560 8262 9596
rect 8206 8608 8262 8664
rect 9034 13504 9090 13560
rect 8390 8336 8446 8392
rect 8574 8064 8630 8120
rect 8298 6704 8354 6760
rect 8206 5752 8262 5808
rect 9218 19372 9274 19408
rect 9218 19352 9220 19372
rect 9220 19352 9272 19372
rect 9272 19352 9274 19372
rect 9494 13640 9550 13696
rect 9218 11056 9274 11112
rect 9218 10104 9274 10160
rect 9218 9172 9274 9208
rect 9678 12008 9734 12064
rect 10506 21392 10562 21448
rect 10230 16904 10286 16960
rect 9678 10956 9680 10976
rect 9680 10956 9732 10976
rect 9732 10956 9734 10976
rect 9678 10920 9734 10956
rect 9954 9968 10010 10024
rect 9494 9288 9550 9344
rect 9218 9152 9220 9172
rect 9220 9152 9272 9172
rect 9272 9152 9274 9172
rect 9218 8880 9274 8936
rect 9678 9288 9734 9344
rect 9126 8064 9182 8120
rect 9586 8064 9642 8120
rect 9586 7928 9642 7984
rect 9494 6976 9550 7032
rect 10046 8064 10102 8120
rect 10138 7928 10194 7984
rect 10506 10512 10562 10568
rect 10782 11464 10838 11520
rect 10506 9288 10562 9344
rect 10506 8744 10562 8800
rect 10322 7928 10378 7984
rect 10230 6568 10286 6624
rect 10506 8200 10562 8256
rect 10598 7540 10654 7576
rect 10598 7520 10600 7540
rect 10600 7520 10652 7540
rect 10652 7520 10654 7540
rect 10506 6024 10562 6080
rect 8942 4800 8998 4856
rect 9402 4820 9458 4856
rect 9402 4800 9404 4820
rect 9404 4800 9456 4820
rect 9456 4800 9458 4820
rect 8298 4664 8354 4720
rect 9402 4684 9458 4720
rect 9402 4664 9404 4684
rect 9404 4664 9456 4684
rect 9456 4664 9458 4684
rect 7930 3168 7986 3224
rect 7838 2488 7894 2544
rect 9310 4140 9366 4176
rect 9310 4120 9312 4140
rect 9312 4120 9364 4140
rect 9364 4120 9366 4140
rect 11058 9968 11114 10024
rect 11058 8744 11114 8800
rect 11058 7420 11060 7440
rect 11060 7420 11112 7440
rect 11112 7420 11114 7440
rect 11058 7384 11114 7420
rect 10782 5636 10838 5672
rect 10782 5616 10784 5636
rect 10784 5616 10836 5636
rect 10836 5616 10838 5636
rect 9678 4664 9734 4720
rect 9586 4156 9588 4176
rect 9588 4156 9640 4176
rect 9640 4156 9642 4176
rect 9586 4120 9642 4156
rect 9770 4020 9772 4040
rect 9772 4020 9824 4040
rect 9824 4020 9826 4040
rect 9770 3984 9826 4020
rect 9770 3712 9826 3768
rect 9494 2080 9550 2136
rect 10506 4392 10562 4448
rect 10230 2760 10286 2816
rect 10966 5344 11022 5400
rect 11150 5888 11206 5944
rect 11518 15136 11574 15192
rect 11334 12688 11390 12744
rect 12254 18148 12310 18184
rect 12254 18128 12256 18148
rect 12256 18128 12308 18148
rect 12308 18128 12310 18148
rect 12530 18148 12586 18184
rect 12530 18128 12532 18148
rect 12532 18128 12584 18148
rect 12584 18128 12586 18148
rect 11334 11192 11390 11248
rect 11702 11076 11758 11112
rect 11702 11056 11704 11076
rect 11704 11056 11756 11076
rect 11756 11056 11758 11076
rect 11518 9832 11574 9888
rect 11426 7964 11428 7984
rect 11428 7964 11480 7984
rect 11480 7964 11482 7984
rect 11426 7928 11482 7964
rect 11426 7656 11482 7712
rect 11426 7112 11482 7168
rect 11518 6976 11574 7032
rect 11150 4800 11206 4856
rect 11058 3984 11114 4040
rect 12070 12824 12126 12880
rect 13818 21256 13874 21312
rect 11886 10920 11942 10976
rect 12070 9832 12126 9888
rect 11886 9152 11942 9208
rect 11978 8744 12034 8800
rect 12070 7948 12126 7984
rect 12070 7928 12072 7948
rect 12072 7928 12124 7948
rect 12124 7928 12126 7948
rect 11978 7520 12034 7576
rect 11886 6976 11942 7032
rect 11610 5480 11666 5536
rect 12346 10920 12402 10976
rect 12438 10784 12494 10840
rect 12346 10104 12402 10160
rect 12254 8744 12310 8800
rect 12254 8200 12310 8256
rect 12530 9152 12586 9208
rect 12530 7928 12586 7984
rect 12346 5344 12402 5400
rect 12162 4392 12218 4448
rect 11978 3848 12034 3904
rect 12714 6024 12770 6080
rect 12714 5616 12770 5672
rect 13174 10548 13176 10568
rect 13176 10548 13228 10568
rect 13228 10548 13230 10568
rect 13174 10512 13230 10548
rect 13358 10512 13414 10568
rect 12898 5480 12954 5536
rect 12806 5344 12862 5400
rect 13174 8200 13230 8256
rect 13174 6024 13230 6080
rect 12530 3304 12586 3360
rect 12990 3304 13046 3360
rect 14002 20304 14058 20360
rect 13634 9832 13690 9888
rect 14278 14864 14334 14920
rect 13450 8880 13506 8936
rect 13726 8200 13782 8256
rect 13450 6568 13506 6624
rect 13726 7792 13782 7848
rect 13634 5344 13690 5400
rect 13542 4664 13598 4720
rect 14002 7112 14058 7168
rect 14922 14592 14978 14648
rect 15106 13640 15162 13696
rect 14554 12688 14610 12744
rect 14462 10804 14518 10840
rect 14462 10784 14464 10804
rect 14464 10784 14516 10804
rect 14516 10784 14518 10804
rect 14370 10512 14426 10568
rect 14830 11464 14886 11520
rect 14830 11192 14886 11248
rect 14370 7792 14426 7848
rect 13450 4392 13506 4448
rect 12162 3032 12218 3088
rect 13082 2896 13138 2952
rect 13358 3032 13414 3088
rect 14830 9696 14886 9752
rect 14462 5344 14518 5400
rect 13542 2624 13598 2680
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 16670 15972 16726 16008
rect 16670 15952 16672 15972
rect 16672 15952 16724 15972
rect 16724 15952 16726 15972
rect 15750 12844 15806 12880
rect 15750 12824 15752 12844
rect 15752 12824 15804 12844
rect 15804 12824 15806 12844
rect 15014 5480 15070 5536
rect 15290 6840 15346 6896
rect 15290 6024 15346 6080
rect 15198 2896 15254 2952
rect 16302 12300 16358 12336
rect 16302 12280 16304 12300
rect 16304 12280 16356 12300
rect 16356 12280 16358 12300
rect 16302 10376 16358 10432
rect 15750 2916 15806 2952
rect 17222 16904 17278 16960
rect 17130 10920 17186 10976
rect 16946 10784 17002 10840
rect 16486 9696 16542 9752
rect 16302 8744 16358 8800
rect 16302 7948 16358 7984
rect 16302 7928 16304 7948
rect 16304 7928 16356 7948
rect 16356 7928 16358 7948
rect 16026 5344 16082 5400
rect 16302 6704 16358 6760
rect 16026 3712 16082 3768
rect 16210 3712 16266 3768
rect 15750 2896 15752 2916
rect 15752 2896 15804 2916
rect 15804 2896 15806 2916
rect 16210 3032 16266 3088
rect 17222 9152 17278 9208
rect 17498 15972 17554 16008
rect 17498 15952 17500 15972
rect 17500 15952 17552 15972
rect 17552 15952 17554 15972
rect 17498 14592 17554 14648
rect 17498 9560 17554 9616
rect 18510 23568 18566 23624
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 18418 14900 18420 14920
rect 18420 14900 18472 14920
rect 18472 14900 18474 14920
rect 18418 14864 18474 14900
rect 17682 9832 17738 9888
rect 17590 7792 17646 7848
rect 17314 7656 17370 7712
rect 17130 7112 17186 7168
rect 16946 4256 17002 4312
rect 17222 5480 17278 5536
rect 17682 7248 17738 7304
rect 17406 5752 17462 5808
rect 17590 5616 17646 5672
rect 17498 4820 17554 4856
rect 17498 4800 17500 4820
rect 17500 4800 17552 4820
rect 17552 4800 17554 4820
rect 18510 10004 18512 10024
rect 18512 10004 18564 10024
rect 18564 10004 18566 10024
rect 18510 9968 18566 10004
rect 17866 8608 17922 8664
rect 18050 8200 18106 8256
rect 17958 8064 18014 8120
rect 18050 6976 18106 7032
rect 18510 8508 18512 8528
rect 18512 8508 18564 8528
rect 18564 8508 18566 8528
rect 18510 8472 18566 8508
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 18970 12280 19026 12336
rect 19062 12144 19118 12200
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 17590 4020 17592 4040
rect 17592 4020 17644 4040
rect 17644 4020 17646 4040
rect 17590 3984 17646 4020
rect 18326 4392 18382 4448
rect 16854 3304 16910 3360
rect 15842 2216 15898 2272
rect 18602 7520 18658 7576
rect 18694 6452 18750 6488
rect 18694 6432 18696 6452
rect 18696 6432 18748 6452
rect 18748 6432 18750 6452
rect 19982 11056 20038 11112
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19246 7384 19302 7440
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 21362 13640 21418 13696
rect 20534 11600 20590 11656
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19430 6024 19486 6080
rect 20074 6332 20076 6352
rect 20076 6332 20128 6352
rect 20128 6332 20130 6352
rect 20074 6296 20130 6332
rect 19338 4936 19394 4992
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19522 5244 19524 5264
rect 19524 5244 19576 5264
rect 19576 5244 19578 5264
rect 19522 5208 19578 5244
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19522 4120 19578 4176
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20074 3848 20130 3904
rect 21086 11736 21142 11792
rect 20810 9424 20866 9480
rect 20902 8336 20958 8392
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 19430 2080 19486 2136
rect 21270 10648 21326 10704
rect 21362 6180 21418 6216
rect 21362 6160 21364 6180
rect 21364 6160 21416 6180
rect 21416 6160 21418 6180
rect 23570 19216 23626 19272
rect 24674 19216 24730 19272
rect 23294 17196 23350 17232
rect 23294 17176 23296 17196
rect 23296 17176 23348 17196
rect 23348 17176 23350 17196
rect 23846 14456 23902 14512
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 38290 38120 38346 38176
rect 38198 36760 38254 36816
rect 38198 34720 38254 34776
rect 38198 33380 38254 33416
rect 38198 33360 38200 33380
rect 38200 33360 38252 33380
rect 38252 33360 38254 33380
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 38290 31320 38346 31376
rect 38290 29960 38346 30016
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 38198 28600 38254 28656
rect 38198 26560 38254 26616
rect 38290 25236 38292 25256
rect 38292 25236 38344 25256
rect 38344 25236 38346 25256
rect 38290 25200 38346 25236
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 38290 23160 38346 23216
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 22466 10240 22522 10296
rect 22834 9016 22890 9072
rect 22098 5908 22154 5944
rect 22098 5888 22100 5908
rect 22100 5888 22152 5908
rect 22152 5888 22154 5908
rect 22098 5092 22154 5128
rect 22098 5072 22100 5092
rect 22100 5072 22152 5092
rect 22152 5072 22154 5092
rect 21454 3732 21510 3768
rect 21454 3712 21456 3732
rect 21456 3712 21508 3732
rect 21508 3712 21510 3732
rect 20810 2624 20866 2680
rect 22098 4548 22154 4584
rect 22098 4528 22100 4548
rect 22100 4528 22152 4548
rect 22152 4528 22154 4548
rect 22098 3596 22154 3632
rect 22098 3576 22100 3596
rect 22100 3576 22152 3596
rect 22152 3576 22154 3596
rect 22098 2796 22100 2816
rect 22100 2796 22152 2816
rect 22152 2796 22154 2816
rect 22098 2760 22154 2796
rect 22190 2352 22246 2408
rect 22282 1264 22338 1320
rect 23478 3476 23480 3496
rect 23480 3476 23532 3496
rect 23532 3476 23534 3496
rect 23478 3440 23534 3476
rect 23938 3032 23994 3088
rect 22742 2508 22798 2544
rect 22742 2488 22744 2508
rect 22744 2488 22796 2508
rect 22796 2488 22798 2508
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 38290 21800 38346 21856
rect 38290 19796 38292 19816
rect 38292 19796 38344 19816
rect 38344 19796 38346 19816
rect 38290 19760 38346 19796
rect 38290 18400 38346 18456
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 38198 17060 38254 17096
rect 38198 17040 38200 17060
rect 38200 17040 38252 17060
rect 38252 17040 38254 17060
rect 38290 15000 38346 15056
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 38198 13676 38200 13696
rect 38200 13676 38252 13696
rect 38252 13676 38254 13696
rect 38198 13640 38254 13676
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 38290 11600 38346 11656
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 33874 7928 33930 7984
rect 38198 10240 38254 10296
rect 38198 8880 38254 8936
rect 23570 1400 23626 1456
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38290 6840 38346 6896
rect 38198 5516 38200 5536
rect 38200 5516 38252 5536
rect 38252 5516 38254 5536
rect 38198 5480 38254 5516
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38290 3476 38292 3496
rect 38292 3476 38344 3496
rect 38344 3476 38346 3496
rect 38290 3440 38346 3476
rect 38198 2080 38254 2136
rect 37278 40 37334 96
<< metal3 >>
rect 200 39538 800 39568
rect 2773 39538 2839 39541
rect 200 39536 2839 39538
rect 200 39480 2778 39536
rect 2834 39480 2839 39536
rect 200 39478 2839 39480
rect 200 39448 800 39478
rect 2773 39475 2839 39478
rect 38285 38178 38351 38181
rect 39200 38178 39800 38208
rect 38285 38176 39800 38178
rect 38285 38120 38290 38176
rect 38346 38120 39800 38176
rect 38285 38118 39800 38120
rect 38285 38115 38351 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 3141 37498 3207 37501
rect 200 37496 3207 37498
rect 200 37440 3146 37496
rect 3202 37440 3207 37496
rect 200 37438 3207 37440
rect 200 37408 800 37438
rect 3141 37435 3207 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 38193 36818 38259 36821
rect 39200 36818 39800 36848
rect 38193 36816 39800 36818
rect 38193 36760 38198 36816
rect 38254 36760 39800 36816
rect 38193 36758 39800 36760
rect 38193 36755 38259 36758
rect 39200 36728 39800 36758
rect 7465 36546 7531 36549
rect 7598 36546 7604 36548
rect 7465 36544 7604 36546
rect 7465 36488 7470 36544
rect 7526 36488 7604 36544
rect 7465 36486 7604 36488
rect 7465 36483 7531 36486
rect 7598 36484 7604 36486
rect 7668 36484 7674 36548
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1761 36138 1827 36141
rect 200 36136 1827 36138
rect 200 36080 1766 36136
rect 1822 36080 1827 36136
rect 200 36078 1827 36080
rect 200 36048 800 36078
rect 1761 36075 1827 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 38193 34778 38259 34781
rect 39200 34778 39800 34808
rect 38193 34776 39800 34778
rect 38193 34720 38198 34776
rect 38254 34720 39800 34776
rect 38193 34718 39800 34720
rect 38193 34715 38259 34718
rect 39200 34688 39800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1761 34098 1827 34101
rect 200 34096 1827 34098
rect 200 34040 1766 34096
rect 1822 34040 1827 34096
rect 200 34038 1827 34040
rect 200 34008 800 34038
rect 1761 34035 1827 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32768
rect 1761 32738 1827 32741
rect 200 32736 1827 32738
rect 200 32680 1766 32736
rect 1822 32680 1827 32736
rect 200 32678 1827 32680
rect 200 32648 800 32678
rect 1761 32675 1827 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 38285 31378 38351 31381
rect 39200 31378 39800 31408
rect 38285 31376 39800 31378
rect 38285 31320 38290 31376
rect 38346 31320 39800 31376
rect 38285 31318 39800 31320
rect 38285 31315 38351 31318
rect 39200 31288 39800 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38285 30018 38351 30021
rect 39200 30018 39800 30048
rect 38285 30016 39800 30018
rect 38285 29960 38290 30016
rect 38346 29960 39800 30016
rect 38285 29958 39800 29960
rect 38285 29955 38351 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1761 29338 1827 29341
rect 200 29336 1827 29338
rect 200 29280 1766 29336
rect 1822 29280 1827 29336
rect 200 29278 1827 29280
rect 200 29248 800 29278
rect 1761 29275 1827 29278
rect 3918 29004 3924 29068
rect 3988 29066 3994 29068
rect 4061 29066 4127 29069
rect 3988 29064 4127 29066
rect 3988 29008 4066 29064
rect 4122 29008 4127 29064
rect 3988 29006 4127 29008
rect 3988 29004 3994 29006
rect 4061 29003 4127 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 38193 28658 38259 28661
rect 39200 28658 39800 28688
rect 38193 28656 39800 28658
rect 38193 28600 38198 28656
rect 38254 28600 39800 28656
rect 38193 28598 39800 28600
rect 38193 28595 38259 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 200 27978 800 28008
rect 1761 27978 1827 27981
rect 200 27976 1827 27978
rect 200 27920 1766 27976
rect 1822 27920 1827 27976
rect 200 27918 1827 27920
rect 200 27888 800 27918
rect 1761 27915 1827 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 38193 26618 38259 26621
rect 39200 26618 39800 26648
rect 38193 26616 39800 26618
rect 38193 26560 38198 26616
rect 38254 26560 39800 26616
rect 38193 26558 39800 26560
rect 38193 26555 38259 26558
rect 39200 26528 39800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25938 800 25968
rect 1761 25938 1827 25941
rect 200 25936 1827 25938
rect 200 25880 1766 25936
rect 1822 25880 1827 25936
rect 200 25878 1827 25880
rect 200 25848 800 25878
rect 1761 25875 1827 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 38285 25258 38351 25261
rect 39200 25258 39800 25288
rect 38285 25256 39800 25258
rect 38285 25200 38290 25256
rect 38346 25200 39800 25256
rect 38285 25198 39800 25200
rect 38285 25195 38351 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 200 24578 800 24608
rect 1761 24578 1827 24581
rect 200 24576 1827 24578
rect 200 24520 1766 24576
rect 1822 24520 1827 24576
rect 200 24518 1827 24520
rect 200 24488 800 24518
rect 1761 24515 1827 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 12014 23564 12020 23628
rect 12084 23626 12090 23628
rect 18505 23626 18571 23629
rect 12084 23624 18571 23626
rect 12084 23568 18510 23624
rect 18566 23568 18571 23624
rect 12084 23566 18571 23568
rect 12084 23564 12090 23566
rect 18505 23563 18571 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 38285 23218 38351 23221
rect 39200 23218 39800 23248
rect 38285 23216 39800 23218
rect 38285 23160 38290 23216
rect 38346 23160 39800 23216
rect 38285 23158 39800 23160
rect 38285 23155 38351 23158
rect 39200 23128 39800 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 38285 21858 38351 21861
rect 39200 21858 39800 21888
rect 38285 21856 39800 21858
rect 38285 21800 38290 21856
rect 38346 21800 39800 21856
rect 38285 21798 39800 21800
rect 38285 21795 38351 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 10501 21452 10567 21453
rect 10501 21450 10548 21452
rect 10456 21448 10548 21450
rect 10456 21392 10506 21448
rect 10456 21390 10548 21392
rect 10501 21388 10548 21390
rect 10612 21388 10618 21452
rect 10501 21387 10567 21388
rect 5758 21252 5764 21316
rect 5828 21314 5834 21316
rect 13813 21314 13879 21317
rect 5828 21312 13879 21314
rect 5828 21256 13818 21312
rect 13874 21256 13879 21312
rect 5828 21254 13879 21256
rect 5828 21252 5834 21254
rect 13813 21251 13879 21254
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1761 21178 1827 21181
rect 200 21176 1827 21178
rect 200 21120 1766 21176
rect 1822 21120 1827 21176
rect 200 21118 1827 21120
rect 200 21088 800 21118
rect 1761 21115 1827 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 2405 20362 2471 20365
rect 13997 20362 14063 20365
rect 2405 20360 14063 20362
rect 2405 20304 2410 20360
rect 2466 20304 14002 20360
rect 14058 20304 14063 20360
rect 2405 20302 14063 20304
rect 2405 20299 2471 20302
rect 13997 20299 14063 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 200 19818 800 19848
rect 1761 19818 1827 19821
rect 200 19816 1827 19818
rect 200 19760 1766 19816
rect 1822 19760 1827 19816
rect 200 19758 1827 19760
rect 200 19728 800 19758
rect 1761 19755 1827 19758
rect 38285 19818 38351 19821
rect 39200 19818 39800 19848
rect 38285 19816 39800 19818
rect 38285 19760 38290 19816
rect 38346 19760 39800 19816
rect 38285 19758 39800 19760
rect 38285 19755 38351 19758
rect 39200 19728 39800 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 9213 19410 9279 19413
rect 9438 19410 9444 19412
rect 9213 19408 9444 19410
rect 9213 19352 9218 19408
rect 9274 19352 9444 19408
rect 9213 19350 9444 19352
rect 9213 19347 9279 19350
rect 9438 19348 9444 19350
rect 9508 19348 9514 19412
rect 5942 19212 5948 19276
rect 6012 19274 6018 19276
rect 23565 19274 23631 19277
rect 24669 19274 24735 19277
rect 6012 19272 24735 19274
rect 6012 19216 23570 19272
rect 23626 19216 24674 19272
rect 24730 19216 24735 19272
rect 6012 19214 24735 19216
rect 6012 19212 6018 19214
rect 23565 19211 23631 19214
rect 24669 19211 24735 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 38285 18458 38351 18461
rect 39200 18458 39800 18488
rect 38285 18456 39800 18458
rect 38285 18400 38290 18456
rect 38346 18400 39800 18456
rect 38285 18398 39800 18400
rect 38285 18395 38351 18398
rect 39200 18368 39800 18398
rect 12249 18186 12315 18189
rect 12525 18186 12591 18189
rect 12249 18184 12591 18186
rect 12249 18128 12254 18184
rect 12310 18128 12530 18184
rect 12586 18128 12591 18184
rect 12249 18126 12591 18128
rect 12249 18123 12315 18126
rect 12525 18123 12591 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1761 17778 1827 17781
rect 200 17776 1827 17778
rect 200 17720 1766 17776
rect 1822 17720 1827 17776
rect 200 17718 1827 17720
rect 200 17688 800 17718
rect 1761 17715 1827 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 15878 17172 15884 17236
rect 15948 17234 15954 17236
rect 23289 17234 23355 17237
rect 15948 17232 23355 17234
rect 15948 17176 23294 17232
rect 23350 17176 23355 17232
rect 15948 17174 23355 17176
rect 15948 17172 15954 17174
rect 23289 17171 23355 17174
rect 3325 17098 3391 17101
rect 15326 17098 15332 17100
rect 3325 17096 15332 17098
rect 3325 17040 3330 17096
rect 3386 17040 15332 17096
rect 3325 17038 15332 17040
rect 3325 17035 3391 17038
rect 15326 17036 15332 17038
rect 15396 17036 15402 17100
rect 38193 17098 38259 17101
rect 39200 17098 39800 17128
rect 38193 17096 39800 17098
rect 38193 17040 38198 17096
rect 38254 17040 39800 17096
rect 38193 17038 39800 17040
rect 38193 17035 38259 17038
rect 39200 17008 39800 17038
rect 10225 16962 10291 16965
rect 17217 16962 17283 16965
rect 10225 16960 17283 16962
rect 10225 16904 10230 16960
rect 10286 16904 17222 16960
rect 17278 16904 17283 16960
rect 10225 16902 17283 16904
rect 10225 16899 10291 16902
rect 17217 16899 17283 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 2681 16828 2747 16829
rect 2630 16826 2636 16828
rect 2590 16766 2636 16826
rect 2700 16824 2747 16828
rect 2742 16768 2747 16824
rect 2630 16764 2636 16766
rect 2700 16764 2747 16768
rect 2681 16763 2747 16764
rect 200 16418 800 16448
rect 1761 16418 1827 16421
rect 200 16416 1827 16418
rect 200 16360 1766 16416
rect 1822 16360 1827 16416
rect 200 16358 1827 16360
rect 200 16328 800 16358
rect 1761 16355 1827 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4429 16010 4495 16013
rect 4654 16010 4660 16012
rect 4429 16008 4660 16010
rect 4429 15952 4434 16008
rect 4490 15952 4660 16008
rect 4429 15950 4660 15952
rect 4429 15947 4495 15950
rect 4654 15948 4660 15950
rect 4724 15948 4730 16012
rect 16665 16010 16731 16013
rect 17493 16010 17559 16013
rect 16665 16008 17559 16010
rect 16665 15952 16670 16008
rect 16726 15952 17498 16008
rect 17554 15952 17559 16008
rect 16665 15950 17559 15952
rect 16665 15947 16731 15950
rect 17493 15947 17559 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 2446 15404 2452 15468
rect 2516 15466 2522 15468
rect 2681 15466 2747 15469
rect 2516 15464 2747 15466
rect 2516 15408 2686 15464
rect 2742 15408 2747 15464
rect 2516 15406 2747 15408
rect 2516 15404 2522 15406
rect 2681 15403 2747 15406
rect 3233 15332 3299 15333
rect 3182 15330 3188 15332
rect 3142 15270 3188 15330
rect 3252 15328 3299 15332
rect 3294 15272 3299 15328
rect 3182 15268 3188 15270
rect 3252 15268 3299 15272
rect 3233 15267 3299 15268
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 8201 15194 8267 15197
rect 11513 15194 11579 15197
rect 8201 15192 11579 15194
rect 8201 15136 8206 15192
rect 8262 15136 11518 15192
rect 11574 15136 11579 15192
rect 8201 15134 11579 15136
rect 8201 15131 8267 15134
rect 11513 15131 11579 15134
rect 38285 15058 38351 15061
rect 39200 15058 39800 15088
rect 38285 15056 39800 15058
rect 38285 15000 38290 15056
rect 38346 15000 39800 15056
rect 38285 14998 39800 15000
rect 38285 14995 38351 14998
rect 39200 14968 39800 14998
rect 14273 14922 14339 14925
rect 18413 14922 18479 14925
rect 14273 14920 18479 14922
rect 14273 14864 14278 14920
rect 14334 14864 18418 14920
rect 18474 14864 18479 14920
rect 14273 14862 18479 14864
rect 14273 14859 14339 14862
rect 18413 14859 18479 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 14917 14650 14983 14653
rect 17493 14650 17559 14653
rect 14917 14648 17559 14650
rect 14917 14592 14922 14648
rect 14978 14592 17498 14648
rect 17554 14592 17559 14648
rect 14917 14590 17559 14592
rect 14917 14587 14983 14590
rect 17493 14587 17559 14590
rect 9254 14452 9260 14516
rect 9324 14514 9330 14516
rect 23841 14514 23907 14517
rect 9324 14512 23907 14514
rect 9324 14456 23846 14512
rect 23902 14456 23907 14512
rect 9324 14454 23907 14456
rect 9324 14452 9330 14454
rect 23841 14451 23907 14454
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 8150 13636 8156 13700
rect 8220 13698 8226 13700
rect 9489 13698 9555 13701
rect 8220 13696 9555 13698
rect 8220 13640 9494 13696
rect 9550 13640 9555 13696
rect 8220 13638 9555 13640
rect 8220 13636 8226 13638
rect 9489 13635 9555 13638
rect 11278 13636 11284 13700
rect 11348 13698 11354 13700
rect 15101 13698 15167 13701
rect 11348 13696 15167 13698
rect 11348 13640 15106 13696
rect 15162 13640 15167 13696
rect 11348 13638 15167 13640
rect 11348 13636 11354 13638
rect 15101 13635 15167 13638
rect 16062 13636 16068 13700
rect 16132 13698 16138 13700
rect 21357 13698 21423 13701
rect 16132 13696 21423 13698
rect 16132 13640 21362 13696
rect 21418 13640 21423 13696
rect 16132 13638 21423 13640
rect 16132 13636 16138 13638
rect 21357 13635 21423 13638
rect 38193 13698 38259 13701
rect 39200 13698 39800 13728
rect 38193 13696 39800 13698
rect 38193 13640 38198 13696
rect 38254 13640 39800 13696
rect 38193 13638 39800 13640
rect 38193 13635 38259 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 9029 13562 9095 13565
rect 9622 13562 9628 13564
rect 9029 13560 9628 13562
rect 9029 13504 9034 13560
rect 9090 13504 9628 13560
rect 9029 13502 9628 13504
rect 9029 13499 9095 13502
rect 9622 13500 9628 13502
rect 9692 13500 9698 13564
rect 4153 13290 4219 13293
rect 5441 13290 5507 13293
rect 4153 13288 5507 13290
rect 4153 13232 4158 13288
rect 4214 13232 5446 13288
rect 5502 13232 5507 13288
rect 4153 13230 5507 13232
rect 4153 13227 4219 13230
rect 5441 13227 5507 13230
rect 4429 13154 4495 13157
rect 7557 13154 7623 13157
rect 4429 13152 7623 13154
rect 4429 13096 4434 13152
rect 4490 13096 7562 13152
rect 7618 13096 7623 13152
rect 4429 13094 7623 13096
rect 4429 13091 4495 13094
rect 7557 13091 7623 13094
rect 19570 13088 19886 13089
rect 200 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 1761 13018 1827 13021
rect 5257 13020 5323 13021
rect 200 13016 1827 13018
rect 200 12960 1766 13016
rect 1822 12960 1827 13016
rect 200 12958 1827 12960
rect 200 12928 800 12958
rect 1761 12955 1827 12958
rect 5206 12956 5212 13020
rect 5276 13018 5323 13020
rect 5276 13016 5368 13018
rect 5318 12960 5368 13016
rect 5276 12958 5368 12960
rect 5276 12956 5323 12958
rect 5257 12955 5323 12956
rect 12065 12882 12131 12885
rect 15745 12882 15811 12885
rect 12065 12880 15811 12882
rect 12065 12824 12070 12880
rect 12126 12824 15750 12880
rect 15806 12824 15811 12880
rect 12065 12822 15811 12824
rect 12065 12819 12131 12822
rect 15745 12819 15811 12822
rect 1945 12746 2011 12749
rect 7373 12746 7439 12749
rect 1945 12744 7439 12746
rect 1945 12688 1950 12744
rect 2006 12688 7378 12744
rect 7434 12688 7439 12744
rect 1945 12686 7439 12688
rect 1945 12683 2011 12686
rect 7373 12683 7439 12686
rect 11329 12746 11395 12749
rect 14549 12746 14615 12749
rect 11329 12744 14615 12746
rect 11329 12688 11334 12744
rect 11390 12688 14554 12744
rect 14610 12688 14615 12744
rect 11329 12686 14615 12688
rect 11329 12683 11395 12686
rect 14549 12683 14615 12686
rect 5257 12610 5323 12613
rect 5390 12610 5396 12612
rect 5257 12608 5396 12610
rect 5257 12552 5262 12608
rect 5318 12552 5396 12608
rect 5257 12550 5396 12552
rect 5257 12547 5323 12550
rect 5390 12548 5396 12550
rect 5460 12548 5466 12612
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 5206 12276 5212 12340
rect 5276 12338 5282 12340
rect 5441 12338 5507 12341
rect 5276 12336 5507 12338
rect 5276 12280 5446 12336
rect 5502 12280 5507 12336
rect 5276 12278 5507 12280
rect 5276 12276 5282 12278
rect 5441 12275 5507 12278
rect 16297 12338 16363 12341
rect 18965 12338 19031 12341
rect 16297 12336 19031 12338
rect 16297 12280 16302 12336
rect 16358 12280 18970 12336
rect 19026 12280 19031 12336
rect 16297 12278 19031 12280
rect 16297 12275 16363 12278
rect 18965 12275 19031 12278
rect 2773 12202 2839 12205
rect 3233 12202 3299 12205
rect 2773 12200 3299 12202
rect 2773 12144 2778 12200
rect 2834 12144 3238 12200
rect 3294 12144 3299 12200
rect 2773 12142 3299 12144
rect 2773 12139 2839 12142
rect 3233 12139 3299 12142
rect 4061 12202 4127 12205
rect 19057 12202 19123 12205
rect 4061 12200 19123 12202
rect 4061 12144 4066 12200
rect 4122 12144 19062 12200
rect 19118 12144 19123 12200
rect 4061 12142 19123 12144
rect 4061 12139 4127 12142
rect 19057 12139 19123 12142
rect 3049 12066 3115 12069
rect 9673 12066 9739 12069
rect 3049 12064 9739 12066
rect 3049 12008 3054 12064
rect 3110 12008 9678 12064
rect 9734 12008 9739 12064
rect 3049 12006 9739 12008
rect 3049 12003 3115 12006
rect 9673 12003 9739 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 3918 11868 3924 11932
rect 3988 11930 3994 11932
rect 4245 11930 4311 11933
rect 3988 11928 4311 11930
rect 3988 11872 4250 11928
rect 4306 11872 4311 11928
rect 3988 11870 4311 11872
rect 3988 11868 3994 11870
rect 4245 11867 4311 11870
rect 6269 11930 6335 11933
rect 6637 11930 6703 11933
rect 6269 11928 6703 11930
rect 6269 11872 6274 11928
rect 6330 11872 6642 11928
rect 6698 11872 6703 11928
rect 6269 11870 6703 11872
rect 6269 11867 6335 11870
rect 6637 11867 6703 11870
rect 4061 11794 4127 11797
rect 21081 11794 21147 11797
rect 4061 11792 21147 11794
rect 4061 11736 4066 11792
rect 4122 11736 21086 11792
rect 21142 11736 21147 11792
rect 4061 11734 21147 11736
rect 4061 11731 4127 11734
rect 21081 11731 21147 11734
rect 2681 11658 2747 11661
rect 4889 11658 4955 11661
rect 2681 11656 4955 11658
rect 2681 11600 2686 11656
rect 2742 11600 4894 11656
rect 4950 11600 4955 11656
rect 2681 11598 4955 11600
rect 2681 11595 2747 11598
rect 4889 11595 4955 11598
rect 5809 11658 5875 11661
rect 20529 11658 20595 11661
rect 5809 11656 20595 11658
rect 5809 11600 5814 11656
rect 5870 11600 20534 11656
rect 20590 11600 20595 11656
rect 5809 11598 20595 11600
rect 5809 11595 5875 11598
rect 20529 11595 20595 11598
rect 38285 11658 38351 11661
rect 39200 11658 39800 11688
rect 38285 11656 39800 11658
rect 38285 11600 38290 11656
rect 38346 11600 39800 11656
rect 38285 11598 39800 11600
rect 38285 11595 38351 11598
rect 39200 11568 39800 11598
rect 6177 11522 6243 11525
rect 8109 11522 8175 11525
rect 6177 11520 8175 11522
rect 6177 11464 6182 11520
rect 6238 11464 8114 11520
rect 8170 11464 8175 11520
rect 6177 11462 8175 11464
rect 6177 11459 6243 11462
rect 8109 11459 8175 11462
rect 10777 11522 10843 11525
rect 14825 11522 14891 11525
rect 10777 11520 14891 11522
rect 10777 11464 10782 11520
rect 10838 11464 14830 11520
rect 14886 11464 14891 11520
rect 10777 11462 14891 11464
rect 10777 11459 10843 11462
rect 14825 11459 14891 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 11329 11250 11395 11253
rect 14825 11250 14891 11253
rect 11329 11248 14891 11250
rect 11329 11192 11334 11248
rect 11390 11192 14830 11248
rect 14886 11192 14891 11248
rect 11329 11190 14891 11192
rect 11329 11187 11395 11190
rect 14825 11187 14891 11190
rect 2681 11116 2747 11117
rect 2630 11114 2636 11116
rect 2590 11054 2636 11114
rect 2700 11112 2747 11116
rect 2742 11056 2747 11112
rect 2630 11052 2636 11054
rect 2700 11052 2747 11056
rect 2681 11051 2747 11052
rect 3601 11114 3667 11117
rect 9213 11114 9279 11117
rect 3601 11112 9279 11114
rect 3601 11056 3606 11112
rect 3662 11056 9218 11112
rect 9274 11056 9279 11112
rect 3601 11054 9279 11056
rect 3601 11051 3667 11054
rect 9213 11051 9279 11054
rect 11697 11114 11763 11117
rect 19977 11114 20043 11117
rect 11697 11112 20043 11114
rect 11697 11056 11702 11112
rect 11758 11056 19982 11112
rect 20038 11056 20043 11112
rect 11697 11054 20043 11056
rect 11697 11051 11763 11054
rect 19977 11051 20043 11054
rect 200 10978 800 11008
rect 3601 10978 3667 10981
rect 200 10976 3667 10978
rect 200 10920 3606 10976
rect 3662 10920 3667 10976
rect 200 10918 3667 10920
rect 200 10888 800 10918
rect 3601 10915 3667 10918
rect 9673 10978 9739 10981
rect 11881 10978 11947 10981
rect 9673 10976 11947 10978
rect 9673 10920 9678 10976
rect 9734 10920 11886 10976
rect 11942 10920 11947 10976
rect 9673 10918 11947 10920
rect 9673 10915 9739 10918
rect 11881 10915 11947 10918
rect 12341 10978 12407 10981
rect 17125 10978 17191 10981
rect 12341 10976 17191 10978
rect 12341 10920 12346 10976
rect 12402 10920 17130 10976
rect 17186 10920 17191 10976
rect 12341 10918 17191 10920
rect 12341 10915 12407 10918
rect 17125 10915 17191 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 12433 10842 12499 10845
rect 2730 10840 12499 10842
rect 2730 10784 12438 10840
rect 12494 10784 12499 10840
rect 2730 10782 12499 10784
rect 2446 10644 2452 10708
rect 2516 10706 2522 10708
rect 2730 10706 2790 10782
rect 12433 10779 12499 10782
rect 14457 10842 14523 10845
rect 16941 10842 17007 10845
rect 14457 10840 17007 10842
rect 14457 10784 14462 10840
rect 14518 10784 16946 10840
rect 17002 10784 17007 10840
rect 14457 10782 17007 10784
rect 14457 10779 14523 10782
rect 16941 10779 17007 10782
rect 2516 10646 2790 10706
rect 5441 10706 5507 10709
rect 21265 10706 21331 10709
rect 5441 10704 21331 10706
rect 5441 10648 5446 10704
rect 5502 10648 21270 10704
rect 21326 10648 21331 10704
rect 5441 10646 21331 10648
rect 2516 10644 2522 10646
rect 5441 10643 5507 10646
rect 21265 10643 21331 10646
rect 10501 10570 10567 10573
rect 13169 10570 13235 10573
rect 10501 10568 13235 10570
rect 10501 10512 10506 10568
rect 10562 10512 13174 10568
rect 13230 10512 13235 10568
rect 10501 10510 13235 10512
rect 10501 10507 10567 10510
rect 13169 10507 13235 10510
rect 13353 10570 13419 10573
rect 14365 10570 14431 10573
rect 13353 10568 14431 10570
rect 13353 10512 13358 10568
rect 13414 10512 14370 10568
rect 14426 10512 14431 10568
rect 13353 10510 14431 10512
rect 13353 10507 13419 10510
rect 14365 10507 14431 10510
rect 5993 10434 6059 10437
rect 16297 10434 16363 10437
rect 5993 10432 16363 10434
rect 5993 10376 5998 10432
rect 6054 10376 16302 10432
rect 16358 10376 16363 10432
rect 5993 10374 16363 10376
rect 5993 10371 6059 10374
rect 16297 10371 16363 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 7833 10298 7899 10301
rect 22461 10298 22527 10301
rect 7833 10296 22527 10298
rect 7833 10240 7838 10296
rect 7894 10240 22466 10296
rect 22522 10240 22527 10296
rect 7833 10238 22527 10240
rect 7833 10235 7899 10238
rect 22461 10235 22527 10238
rect 38193 10298 38259 10301
rect 39200 10298 39800 10328
rect 38193 10296 39800 10298
rect 38193 10240 38198 10296
rect 38254 10240 39800 10296
rect 38193 10238 39800 10240
rect 38193 10235 38259 10238
rect 39200 10208 39800 10238
rect 4521 10162 4587 10165
rect 4654 10162 4660 10164
rect 4521 10160 4660 10162
rect 4521 10104 4526 10160
rect 4582 10104 4660 10160
rect 4521 10102 4660 10104
rect 4521 10099 4587 10102
rect 4654 10100 4660 10102
rect 4724 10100 4730 10164
rect 9213 10162 9279 10165
rect 12341 10162 12407 10165
rect 9213 10160 12407 10162
rect 9213 10104 9218 10160
rect 9274 10104 12346 10160
rect 12402 10104 12407 10160
rect 9213 10102 12407 10104
rect 9213 10099 9279 10102
rect 12341 10099 12407 10102
rect 9949 10026 10015 10029
rect 11053 10026 11119 10029
rect 18505 10026 18571 10029
rect 9949 10024 18571 10026
rect 9949 9968 9954 10024
rect 10010 9968 11058 10024
rect 11114 9968 18510 10024
rect 18566 9968 18571 10024
rect 9949 9966 18571 9968
rect 9949 9963 10015 9966
rect 11053 9963 11119 9966
rect 18505 9963 18571 9966
rect 6453 9890 6519 9893
rect 11513 9890 11579 9893
rect 6453 9888 11579 9890
rect 6453 9832 6458 9888
rect 6514 9832 11518 9888
rect 11574 9832 11579 9888
rect 6453 9830 11579 9832
rect 6453 9827 6519 9830
rect 11513 9827 11579 9830
rect 12065 9890 12131 9893
rect 13629 9890 13695 9893
rect 17677 9890 17743 9893
rect 12065 9888 17743 9890
rect 12065 9832 12070 9888
rect 12126 9832 13634 9888
rect 13690 9832 17682 9888
rect 17738 9832 17743 9888
rect 12065 9830 17743 9832
rect 12065 9827 12131 9830
rect 13629 9827 13695 9830
rect 17677 9827 17743 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 3049 9754 3115 9757
rect 3182 9754 3188 9756
rect 3049 9752 3188 9754
rect 3049 9696 3054 9752
rect 3110 9696 3188 9752
rect 3049 9694 3188 9696
rect 3049 9691 3115 9694
rect 3182 9692 3188 9694
rect 3252 9692 3258 9756
rect 14825 9754 14891 9757
rect 16481 9754 16547 9757
rect 14825 9752 16547 9754
rect 14825 9696 14830 9752
rect 14886 9696 16486 9752
rect 16542 9696 16547 9752
rect 14825 9694 16547 9696
rect 14825 9691 14891 9694
rect 16481 9691 16547 9694
rect 200 9618 800 9648
rect 3877 9618 3943 9621
rect 7598 9618 7604 9620
rect 200 9616 3943 9618
rect 200 9560 3882 9616
rect 3938 9560 3943 9616
rect 200 9558 3943 9560
rect 200 9528 800 9558
rect 3877 9555 3943 9558
rect 4662 9558 7604 9618
rect 1853 9482 1919 9485
rect 4662 9482 4722 9558
rect 7598 9556 7604 9558
rect 7668 9556 7674 9620
rect 8201 9618 8267 9621
rect 17493 9618 17559 9621
rect 8201 9616 17559 9618
rect 8201 9560 8206 9616
rect 8262 9560 17498 9616
rect 17554 9560 17559 9616
rect 8201 9558 17559 9560
rect 8201 9555 8267 9558
rect 17493 9555 17559 9558
rect 1853 9480 4722 9482
rect 1853 9424 1858 9480
rect 1914 9424 4722 9480
rect 1853 9422 4722 9424
rect 4797 9482 4863 9485
rect 20805 9482 20871 9485
rect 4797 9480 20871 9482
rect 4797 9424 4802 9480
rect 4858 9424 20810 9480
rect 20866 9424 20871 9480
rect 4797 9422 20871 9424
rect 1853 9419 1919 9422
rect 4797 9419 4863 9422
rect 20805 9419 20871 9422
rect 9070 9284 9076 9348
rect 9140 9346 9146 9348
rect 9489 9346 9555 9349
rect 9140 9344 9555 9346
rect 9140 9288 9494 9344
rect 9550 9288 9555 9344
rect 9140 9286 9555 9288
rect 9140 9284 9146 9286
rect 9489 9283 9555 9286
rect 9673 9346 9739 9349
rect 10501 9346 10567 9349
rect 9673 9344 10567 9346
rect 9673 9288 9678 9344
rect 9734 9288 10506 9344
rect 10562 9288 10567 9344
rect 9673 9286 10567 9288
rect 9673 9283 9739 9286
rect 10501 9283 10567 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 5717 9212 5783 9213
rect 5717 9210 5764 9212
rect 5672 9208 5764 9210
rect 5672 9152 5722 9208
rect 5672 9150 5764 9152
rect 5717 9148 5764 9150
rect 5828 9148 5834 9212
rect 9213 9210 9279 9213
rect 11881 9210 11947 9213
rect 9213 9208 11947 9210
rect 9213 9152 9218 9208
rect 9274 9152 11886 9208
rect 11942 9152 11947 9208
rect 9213 9150 11947 9152
rect 5717 9147 5783 9148
rect 9213 9147 9279 9150
rect 11881 9147 11947 9150
rect 12525 9210 12591 9213
rect 17217 9210 17283 9213
rect 12525 9208 17283 9210
rect 12525 9152 12530 9208
rect 12586 9152 17222 9208
rect 17278 9152 17283 9208
rect 12525 9150 17283 9152
rect 12525 9147 12591 9150
rect 17217 9147 17283 9150
rect 3325 9074 3391 9077
rect 4521 9074 4587 9077
rect 22829 9074 22895 9077
rect 3325 9072 22895 9074
rect 3325 9016 3330 9072
rect 3386 9016 4526 9072
rect 4582 9016 22834 9072
rect 22890 9016 22895 9072
rect 3325 9014 22895 9016
rect 3325 9011 3391 9014
rect 4521 9011 4587 9014
rect 22829 9011 22895 9014
rect 9213 8938 9279 8941
rect 10542 8938 10548 8940
rect 9213 8936 10548 8938
rect 9213 8880 9218 8936
rect 9274 8880 10548 8936
rect 9213 8878 10548 8880
rect 9213 8875 9279 8878
rect 10542 8876 10548 8878
rect 10612 8938 10618 8940
rect 13445 8938 13511 8941
rect 10612 8936 13511 8938
rect 10612 8880 13450 8936
rect 13506 8880 13511 8936
rect 10612 8878 13511 8880
rect 10612 8876 10618 8878
rect 13445 8875 13511 8878
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 6269 8802 6335 8805
rect 10501 8802 10567 8805
rect 6269 8800 10567 8802
rect 6269 8744 6274 8800
rect 6330 8744 10506 8800
rect 10562 8744 10567 8800
rect 6269 8742 10567 8744
rect 6269 8739 6335 8742
rect 10501 8739 10567 8742
rect 11053 8802 11119 8805
rect 11973 8804 12039 8805
rect 11973 8802 12020 8804
rect 11053 8800 12020 8802
rect 11053 8744 11058 8800
rect 11114 8744 11978 8800
rect 11053 8742 12020 8744
rect 11053 8739 11119 8742
rect 11973 8740 12020 8742
rect 12084 8740 12090 8804
rect 12249 8802 12315 8805
rect 16297 8802 16363 8805
rect 12249 8800 16363 8802
rect 12249 8744 12254 8800
rect 12310 8744 16302 8800
rect 16358 8744 16363 8800
rect 12249 8742 16363 8744
rect 11973 8739 12039 8740
rect 12249 8739 12315 8742
rect 16297 8739 16363 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 8201 8666 8267 8669
rect 17861 8666 17927 8669
rect 8201 8664 17927 8666
rect 8201 8608 8206 8664
rect 8262 8608 17866 8664
rect 17922 8608 17927 8664
rect 8201 8606 17927 8608
rect 8201 8603 8267 8606
rect 17861 8603 17927 8606
rect 3325 8530 3391 8533
rect 18505 8530 18571 8533
rect 3325 8528 18571 8530
rect 3325 8472 3330 8528
rect 3386 8472 18510 8528
rect 18566 8472 18571 8528
rect 3325 8470 18571 8472
rect 3325 8467 3391 8470
rect 18505 8467 18571 8470
rect 8385 8394 8451 8397
rect 20897 8394 20963 8397
rect 8385 8392 20963 8394
rect 8385 8336 8390 8392
rect 8446 8336 20902 8392
rect 20958 8336 20963 8392
rect 8385 8334 20963 8336
rect 8385 8331 8451 8334
rect 20897 8331 20963 8334
rect 200 8258 800 8288
rect 3693 8258 3759 8261
rect 200 8256 3759 8258
rect 200 8200 3698 8256
rect 3754 8200 3759 8256
rect 200 8198 3759 8200
rect 200 8168 800 8198
rect 3693 8195 3759 8198
rect 9622 8196 9628 8260
rect 9692 8258 9698 8260
rect 10501 8258 10567 8261
rect 9692 8256 10567 8258
rect 9692 8200 10506 8256
rect 10562 8200 10567 8256
rect 9692 8198 10567 8200
rect 9692 8196 9698 8198
rect 10501 8195 10567 8198
rect 12249 8258 12315 8261
rect 13169 8258 13235 8261
rect 12249 8256 13235 8258
rect 12249 8200 12254 8256
rect 12310 8200 13174 8256
rect 13230 8200 13235 8256
rect 12249 8198 13235 8200
rect 12249 8195 12315 8198
rect 13169 8195 13235 8198
rect 13721 8258 13787 8261
rect 18045 8258 18111 8261
rect 13721 8256 18111 8258
rect 13721 8200 13726 8256
rect 13782 8200 18050 8256
rect 18106 8200 18111 8256
rect 13721 8198 18111 8200
rect 13721 8195 13787 8198
rect 18045 8195 18111 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 7281 8122 7347 8125
rect 8150 8122 8156 8124
rect 7281 8120 8156 8122
rect 7281 8064 7286 8120
rect 7342 8064 8156 8120
rect 7281 8062 8156 8064
rect 7281 8059 7347 8062
rect 8150 8060 8156 8062
rect 8220 8060 8226 8124
rect 8569 8122 8635 8125
rect 9121 8122 9187 8125
rect 9581 8122 9647 8125
rect 8569 8120 9647 8122
rect 8569 8064 8574 8120
rect 8630 8064 9126 8120
rect 9182 8064 9586 8120
rect 9642 8064 9647 8120
rect 8569 8062 9647 8064
rect 3877 7986 3943 7989
rect 6453 7986 6519 7989
rect 3877 7984 6519 7986
rect 3877 7928 3882 7984
rect 3938 7928 6458 7984
rect 6514 7928 6519 7984
rect 3877 7926 6519 7928
rect 3877 7923 3943 7926
rect 6453 7923 6519 7926
rect 8158 7850 8218 8060
rect 8569 8059 8635 8062
rect 9121 8059 9187 8062
rect 9581 8059 9647 8062
rect 10041 8122 10107 8125
rect 17953 8122 18019 8125
rect 10041 8120 18019 8122
rect 10041 8064 10046 8120
rect 10102 8064 17958 8120
rect 18014 8064 18019 8120
rect 10041 8062 18019 8064
rect 10041 8059 10107 8062
rect 17953 8059 18019 8062
rect 9070 7924 9076 7988
rect 9140 7986 9146 7988
rect 9581 7986 9647 7989
rect 9140 7984 9647 7986
rect 9140 7928 9586 7984
rect 9642 7928 9647 7984
rect 9140 7926 9647 7928
rect 9140 7924 9146 7926
rect 9581 7923 9647 7926
rect 10133 7986 10199 7989
rect 10317 7986 10383 7989
rect 11421 7986 11487 7989
rect 10133 7984 11487 7986
rect 10133 7928 10138 7984
rect 10194 7928 10322 7984
rect 10378 7928 11426 7984
rect 11482 7928 11487 7984
rect 10133 7926 11487 7928
rect 10133 7923 10199 7926
rect 10317 7923 10383 7926
rect 11421 7923 11487 7926
rect 12065 7986 12131 7989
rect 12525 7986 12591 7989
rect 12065 7984 12591 7986
rect 12065 7928 12070 7984
rect 12126 7928 12530 7984
rect 12586 7928 12591 7984
rect 12065 7926 12591 7928
rect 12065 7923 12131 7926
rect 12525 7923 12591 7926
rect 16297 7986 16363 7989
rect 33869 7986 33935 7989
rect 16297 7984 33935 7986
rect 16297 7928 16302 7984
rect 16358 7928 33874 7984
rect 33930 7928 33935 7984
rect 16297 7926 33935 7928
rect 16297 7923 16363 7926
rect 33869 7923 33935 7926
rect 13721 7850 13787 7853
rect 8158 7848 13787 7850
rect 8158 7792 13726 7848
rect 13782 7792 13787 7848
rect 8158 7790 13787 7792
rect 13721 7787 13787 7790
rect 14365 7850 14431 7853
rect 17585 7850 17651 7853
rect 14365 7848 17651 7850
rect 14365 7792 14370 7848
rect 14426 7792 17590 7848
rect 17646 7792 17651 7848
rect 14365 7790 17651 7792
rect 14365 7787 14431 7790
rect 17585 7787 17651 7790
rect 11421 7714 11487 7717
rect 17309 7714 17375 7717
rect 11421 7712 17375 7714
rect 11421 7656 11426 7712
rect 11482 7656 17314 7712
rect 17370 7656 17375 7712
rect 11421 7654 17375 7656
rect 11421 7651 11487 7654
rect 17309 7651 17375 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 10593 7578 10659 7581
rect 11973 7578 12039 7581
rect 18597 7578 18663 7581
rect 10593 7576 18663 7578
rect 10593 7520 10598 7576
rect 10654 7520 11978 7576
rect 12034 7520 18602 7576
rect 18658 7520 18663 7576
rect 10593 7518 18663 7520
rect 10593 7515 10659 7518
rect 11973 7515 12039 7518
rect 18597 7515 18663 7518
rect 11053 7442 11119 7445
rect 19241 7442 19307 7445
rect 11053 7440 19307 7442
rect 11053 7384 11058 7440
rect 11114 7384 19246 7440
rect 19302 7384 19307 7440
rect 11053 7382 19307 7384
rect 11053 7379 11119 7382
rect 19241 7379 19307 7382
rect 7281 7306 7347 7309
rect 17677 7306 17743 7309
rect 7281 7304 17743 7306
rect 7281 7248 7286 7304
rect 7342 7248 17682 7304
rect 17738 7248 17743 7304
rect 7281 7246 17743 7248
rect 7281 7243 7347 7246
rect 17677 7243 17743 7246
rect 4613 7170 4679 7173
rect 11278 7170 11284 7172
rect 4613 7168 11284 7170
rect 4613 7112 4618 7168
rect 4674 7112 11284 7168
rect 4613 7110 11284 7112
rect 4613 7107 4679 7110
rect 11278 7108 11284 7110
rect 11348 7170 11354 7172
rect 11421 7170 11487 7173
rect 11348 7168 11487 7170
rect 11348 7112 11426 7168
rect 11482 7112 11487 7168
rect 11348 7110 11487 7112
rect 11348 7108 11354 7110
rect 11421 7107 11487 7110
rect 13997 7170 14063 7173
rect 17125 7170 17191 7173
rect 13997 7168 17191 7170
rect 13997 7112 14002 7168
rect 14058 7112 17130 7168
rect 17186 7112 17191 7168
rect 13997 7110 17191 7112
rect 13997 7107 14063 7110
rect 17125 7107 17191 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 9489 7034 9555 7037
rect 11513 7034 11579 7037
rect 9489 7032 11579 7034
rect 9489 6976 9494 7032
rect 9550 6976 11518 7032
rect 11574 6976 11579 7032
rect 9489 6974 11579 6976
rect 9489 6971 9555 6974
rect 11513 6971 11579 6974
rect 11881 7034 11947 7037
rect 18045 7034 18111 7037
rect 11881 7032 18111 7034
rect 11881 6976 11886 7032
rect 11942 6976 18050 7032
rect 18106 6976 18111 7032
rect 11881 6974 18111 6976
rect 11881 6971 11947 6974
rect 18045 6971 18111 6974
rect 7649 6898 7715 6901
rect 15285 6900 15351 6901
rect 7649 6896 15210 6898
rect 7649 6840 7654 6896
rect 7710 6840 15210 6896
rect 7649 6838 15210 6840
rect 7649 6835 7715 6838
rect 8293 6762 8359 6765
rect 15150 6762 15210 6838
rect 15285 6896 15332 6900
rect 15396 6898 15402 6900
rect 38285 6898 38351 6901
rect 39200 6898 39800 6928
rect 15285 6840 15290 6896
rect 15285 6836 15332 6840
rect 15396 6838 15442 6898
rect 38285 6896 39800 6898
rect 38285 6840 38290 6896
rect 38346 6840 39800 6896
rect 38285 6838 39800 6840
rect 15396 6836 15402 6838
rect 15285 6835 15351 6836
rect 38285 6835 38351 6838
rect 39200 6808 39800 6838
rect 16297 6762 16363 6765
rect 8293 6760 15026 6762
rect 8293 6704 8298 6760
rect 8354 6704 15026 6760
rect 8293 6702 15026 6704
rect 15150 6760 16363 6762
rect 15150 6704 16302 6760
rect 16358 6704 16363 6760
rect 15150 6702 16363 6704
rect 8293 6699 8359 6702
rect 10225 6626 10291 6629
rect 13445 6626 13511 6629
rect 10225 6624 13511 6626
rect 10225 6568 10230 6624
rect 10286 6568 13450 6624
rect 13506 6568 13511 6624
rect 10225 6566 13511 6568
rect 14966 6626 15026 6702
rect 16297 6699 16363 6702
rect 19374 6626 19380 6628
rect 14966 6566 19380 6626
rect 10225 6563 10291 6566
rect 13445 6563 13511 6566
rect 19374 6564 19380 6566
rect 19444 6564 19450 6628
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4061 6490 4127 6493
rect 18689 6490 18755 6493
rect 4061 6488 18755 6490
rect 4061 6432 4066 6488
rect 4122 6432 18694 6488
rect 18750 6432 18755 6488
rect 4061 6430 18755 6432
rect 4061 6427 4127 6430
rect 18689 6427 18755 6430
rect 3417 6354 3483 6357
rect 20069 6354 20135 6357
rect 3417 6352 20135 6354
rect 3417 6296 3422 6352
rect 3478 6296 20074 6352
rect 20130 6296 20135 6352
rect 3417 6294 20135 6296
rect 3417 6291 3483 6294
rect 20069 6291 20135 6294
rect 200 6218 800 6248
rect 3049 6218 3115 6221
rect 200 6216 3115 6218
rect 200 6160 3054 6216
rect 3110 6160 3115 6216
rect 200 6158 3115 6160
rect 200 6128 800 6158
rect 3049 6155 3115 6158
rect 3509 6218 3575 6221
rect 21357 6218 21423 6221
rect 3509 6216 21423 6218
rect 3509 6160 3514 6216
rect 3570 6160 21362 6216
rect 21418 6160 21423 6216
rect 3509 6158 21423 6160
rect 3509 6155 3575 6158
rect 21357 6155 21423 6158
rect 10501 6082 10567 6085
rect 12709 6082 12775 6085
rect 10501 6080 12775 6082
rect 10501 6024 10506 6080
rect 10562 6024 12714 6080
rect 12770 6024 12775 6080
rect 10501 6022 12775 6024
rect 10501 6019 10567 6022
rect 12709 6019 12775 6022
rect 13169 6082 13235 6085
rect 15285 6082 15351 6085
rect 19425 6084 19491 6085
rect 13169 6080 15351 6082
rect 13169 6024 13174 6080
rect 13230 6024 15290 6080
rect 15346 6024 15351 6080
rect 13169 6022 15351 6024
rect 13169 6019 13235 6022
rect 15285 6019 15351 6022
rect 19374 6020 19380 6084
rect 19444 6082 19491 6084
rect 19444 6080 19536 6082
rect 19486 6024 19536 6080
rect 19444 6022 19536 6024
rect 19444 6020 19491 6022
rect 19425 6019 19491 6020
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 11145 5946 11211 5949
rect 22093 5946 22159 5949
rect 11145 5944 22159 5946
rect 11145 5888 11150 5944
rect 11206 5888 22098 5944
rect 22154 5888 22159 5944
rect 11145 5886 22159 5888
rect 11145 5883 11211 5886
rect 22093 5883 22159 5886
rect 1761 5810 1827 5813
rect 4153 5810 4219 5813
rect 1761 5808 4219 5810
rect 1761 5752 1766 5808
rect 1822 5752 4158 5808
rect 4214 5752 4219 5808
rect 1761 5750 4219 5752
rect 1761 5747 1827 5750
rect 4153 5747 4219 5750
rect 8201 5810 8267 5813
rect 17401 5810 17467 5813
rect 8201 5808 17467 5810
rect 8201 5752 8206 5808
rect 8262 5752 17406 5808
rect 17462 5752 17467 5808
rect 8201 5750 17467 5752
rect 8201 5747 8267 5750
rect 17401 5747 17467 5750
rect 9438 5612 9444 5676
rect 9508 5674 9514 5676
rect 10777 5674 10843 5677
rect 9508 5672 10843 5674
rect 9508 5616 10782 5672
rect 10838 5616 10843 5672
rect 9508 5614 10843 5616
rect 9508 5612 9514 5614
rect 10777 5611 10843 5614
rect 12709 5674 12775 5677
rect 17585 5674 17651 5677
rect 12709 5672 17651 5674
rect 12709 5616 12714 5672
rect 12770 5616 17590 5672
rect 17646 5616 17651 5672
rect 12709 5614 17651 5616
rect 12709 5611 12775 5614
rect 17585 5611 17651 5614
rect 11605 5538 11671 5541
rect 12893 5538 12959 5541
rect 11605 5536 12959 5538
rect 11605 5480 11610 5536
rect 11666 5480 12898 5536
rect 12954 5480 12959 5536
rect 11605 5478 12959 5480
rect 11605 5475 11671 5478
rect 12893 5475 12959 5478
rect 15009 5538 15075 5541
rect 17217 5538 17283 5541
rect 15009 5536 17283 5538
rect 15009 5480 15014 5536
rect 15070 5480 17222 5536
rect 17278 5480 17283 5536
rect 15009 5478 17283 5480
rect 15009 5475 15075 5478
rect 17217 5475 17283 5478
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 6913 5402 6979 5405
rect 10961 5402 11027 5405
rect 6913 5400 11027 5402
rect 6913 5344 6918 5400
rect 6974 5344 10966 5400
rect 11022 5344 11027 5400
rect 6913 5342 11027 5344
rect 6913 5339 6979 5342
rect 10961 5339 11027 5342
rect 12341 5402 12407 5405
rect 12801 5402 12867 5405
rect 12341 5400 12867 5402
rect 12341 5344 12346 5400
rect 12402 5344 12806 5400
rect 12862 5344 12867 5400
rect 12341 5342 12867 5344
rect 12341 5339 12407 5342
rect 12801 5339 12867 5342
rect 13629 5402 13695 5405
rect 14457 5402 14523 5405
rect 16021 5402 16087 5405
rect 13629 5400 16087 5402
rect 13629 5344 13634 5400
rect 13690 5344 14462 5400
rect 14518 5344 16026 5400
rect 16082 5344 16087 5400
rect 13629 5342 16087 5344
rect 13629 5339 13695 5342
rect 14457 5339 14523 5342
rect 16021 5339 16087 5342
rect 5349 5266 5415 5269
rect 19517 5266 19583 5269
rect 5349 5264 19583 5266
rect 5349 5208 5354 5264
rect 5410 5208 19522 5264
rect 19578 5208 19583 5264
rect 5349 5206 19583 5208
rect 5349 5203 5415 5206
rect 19517 5203 19583 5206
rect 5390 5068 5396 5132
rect 5460 5130 5466 5132
rect 22093 5130 22159 5133
rect 5460 5128 22159 5130
rect 5460 5072 22098 5128
rect 22154 5072 22159 5128
rect 5460 5070 22159 5072
rect 5460 5068 5466 5070
rect 22093 5067 22159 5070
rect 5073 4994 5139 4997
rect 19333 4994 19399 4997
rect 5073 4992 19399 4994
rect 5073 4936 5078 4992
rect 5134 4936 19338 4992
rect 19394 4936 19399 4992
rect 5073 4934 19399 4936
rect 5073 4931 5139 4934
rect 19333 4931 19399 4934
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1761 4858 1827 4861
rect 200 4856 1827 4858
rect 200 4800 1766 4856
rect 1822 4800 1827 4856
rect 200 4798 1827 4800
rect 200 4768 800 4798
rect 1761 4795 1827 4798
rect 8937 4858 9003 4861
rect 9397 4858 9463 4861
rect 8937 4856 9463 4858
rect 8937 4800 8942 4856
rect 8998 4800 9402 4856
rect 9458 4800 9463 4856
rect 8937 4798 9463 4800
rect 8937 4795 9003 4798
rect 9397 4795 9463 4798
rect 11145 4858 11211 4861
rect 17493 4858 17559 4861
rect 11145 4856 17559 4858
rect 11145 4800 11150 4856
rect 11206 4800 17498 4856
rect 17554 4800 17559 4856
rect 11145 4798 17559 4800
rect 11145 4795 11211 4798
rect 17493 4795 17559 4798
rect 8293 4722 8359 4725
rect 9397 4722 9463 4725
rect 8293 4720 9463 4722
rect 8293 4664 8298 4720
rect 8354 4664 9402 4720
rect 9458 4664 9463 4720
rect 8293 4662 9463 4664
rect 8293 4659 8359 4662
rect 9397 4659 9463 4662
rect 9673 4722 9739 4725
rect 13537 4722 13603 4725
rect 9673 4720 13603 4722
rect 9673 4664 9678 4720
rect 9734 4664 13542 4720
rect 13598 4664 13603 4720
rect 9673 4662 13603 4664
rect 9673 4659 9739 4662
rect 13537 4659 13603 4662
rect 6453 4586 6519 4589
rect 22093 4586 22159 4589
rect 6453 4584 22159 4586
rect 6453 4528 6458 4584
rect 6514 4528 22098 4584
rect 22154 4528 22159 4584
rect 6453 4526 22159 4528
rect 6453 4523 6519 4526
rect 22093 4523 22159 4526
rect 10501 4450 10567 4453
rect 12157 4450 12223 4453
rect 10501 4448 12223 4450
rect 10501 4392 10506 4448
rect 10562 4392 12162 4448
rect 12218 4392 12223 4448
rect 10501 4390 12223 4392
rect 10501 4387 10567 4390
rect 12157 4387 12223 4390
rect 13445 4450 13511 4453
rect 18321 4450 18387 4453
rect 13445 4448 18387 4450
rect 13445 4392 13450 4448
rect 13506 4392 18326 4448
rect 18382 4392 18387 4448
rect 13445 4390 18387 4392
rect 13445 4387 13511 4390
rect 18321 4387 18387 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 5625 4314 5691 4317
rect 16941 4314 17007 4317
rect 5625 4312 17007 4314
rect 5625 4256 5630 4312
rect 5686 4256 16946 4312
rect 17002 4256 17007 4312
rect 5625 4254 17007 4256
rect 5625 4251 5691 4254
rect 16941 4251 17007 4254
rect 6269 4178 6335 4181
rect 9305 4178 9371 4181
rect 6269 4176 9371 4178
rect 6269 4120 6274 4176
rect 6330 4120 9310 4176
rect 9366 4120 9371 4176
rect 6269 4118 9371 4120
rect 6269 4115 6335 4118
rect 9305 4115 9371 4118
rect 9581 4178 9647 4181
rect 19517 4178 19583 4181
rect 9581 4176 19583 4178
rect 9581 4120 9586 4176
rect 9642 4120 19522 4176
rect 19578 4120 19583 4176
rect 9581 4118 19583 4120
rect 9581 4115 9647 4118
rect 19517 4115 19583 4118
rect 5901 4044 5967 4045
rect 5901 4042 5948 4044
rect 5856 4040 5948 4042
rect 5856 3984 5906 4040
rect 5856 3982 5948 3984
rect 5901 3980 5948 3982
rect 6012 3980 6018 4044
rect 9254 3980 9260 4044
rect 9324 4042 9330 4044
rect 9765 4042 9831 4045
rect 9324 4040 9831 4042
rect 9324 3984 9770 4040
rect 9826 3984 9831 4040
rect 9324 3982 9831 3984
rect 9324 3980 9330 3982
rect 5901 3979 5967 3980
rect 9765 3979 9831 3982
rect 11053 4042 11119 4045
rect 17585 4042 17651 4045
rect 11053 4040 17651 4042
rect 11053 3984 11058 4040
rect 11114 3984 17590 4040
rect 17646 3984 17651 4040
rect 11053 3982 17651 3984
rect 11053 3979 11119 3982
rect 17585 3979 17651 3982
rect 7649 3906 7715 3909
rect 11973 3906 12039 3909
rect 20069 3906 20135 3909
rect 7649 3904 12039 3906
rect 7649 3848 7654 3904
rect 7710 3848 11978 3904
rect 12034 3848 12039 3904
rect 7649 3846 12039 3848
rect 7649 3843 7715 3846
rect 11973 3843 12039 3846
rect 15702 3904 20135 3906
rect 15702 3848 20074 3904
rect 20130 3848 20135 3904
rect 15702 3846 20135 3848
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 9765 3770 9831 3773
rect 15702 3770 15762 3846
rect 20069 3843 20135 3846
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 16021 3772 16087 3773
rect 16021 3770 16068 3772
rect 9765 3768 15762 3770
rect 9765 3712 9770 3768
rect 9826 3712 15762 3768
rect 9765 3710 15762 3712
rect 15976 3768 16068 3770
rect 15976 3712 16026 3768
rect 15976 3710 16068 3712
rect 9765 3707 9831 3710
rect 16021 3708 16068 3710
rect 16132 3708 16138 3772
rect 16205 3770 16271 3773
rect 21449 3770 21515 3773
rect 16205 3768 21515 3770
rect 16205 3712 16210 3768
rect 16266 3712 21454 3768
rect 21510 3712 21515 3768
rect 16205 3710 21515 3712
rect 16021 3707 16087 3708
rect 16205 3707 16271 3710
rect 21449 3707 21515 3710
rect 4613 3634 4679 3637
rect 22093 3634 22159 3637
rect 4613 3632 22159 3634
rect 4613 3576 4618 3632
rect 4674 3576 22098 3632
rect 22154 3576 22159 3632
rect 4613 3574 22159 3576
rect 4613 3571 4679 3574
rect 22093 3571 22159 3574
rect 23473 3498 23539 3501
rect 2730 3496 23539 3498
rect 2730 3440 23478 3496
rect 23534 3440 23539 3496
rect 2730 3438 23539 3440
rect 200 2818 800 2848
rect 2730 2818 2790 3438
rect 23473 3435 23539 3438
rect 38285 3498 38351 3501
rect 39200 3498 39800 3528
rect 38285 3496 39800 3498
rect 38285 3440 38290 3496
rect 38346 3440 39800 3496
rect 38285 3438 39800 3440
rect 38285 3435 38351 3438
rect 39200 3408 39800 3438
rect 4153 3362 4219 3365
rect 6821 3362 6887 3365
rect 12525 3362 12591 3365
rect 4153 3360 12591 3362
rect 4153 3304 4158 3360
rect 4214 3304 6826 3360
rect 6882 3304 12530 3360
rect 12586 3304 12591 3360
rect 4153 3302 12591 3304
rect 4153 3299 4219 3302
rect 6821 3299 6887 3302
rect 12525 3299 12591 3302
rect 12985 3362 13051 3365
rect 16849 3362 16915 3365
rect 12985 3360 16915 3362
rect 12985 3304 12990 3360
rect 13046 3304 16854 3360
rect 16910 3304 16915 3360
rect 12985 3302 16915 3304
rect 12985 3299 13051 3302
rect 16849 3299 16915 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 7925 3226 7991 3229
rect 7925 3224 17234 3226
rect 7925 3168 7930 3224
rect 7986 3168 17234 3224
rect 7925 3166 17234 3168
rect 7925 3163 7991 3166
rect 12157 3090 12223 3093
rect 13353 3090 13419 3093
rect 16205 3090 16271 3093
rect 12157 3088 13419 3090
rect 12157 3032 12162 3088
rect 12218 3032 13358 3088
rect 13414 3032 13419 3088
rect 12157 3030 13419 3032
rect 12157 3027 12223 3030
rect 13353 3027 13419 3030
rect 15012 3088 16271 3090
rect 15012 3032 16210 3088
rect 16266 3032 16271 3088
rect 15012 3030 16271 3032
rect 17174 3090 17234 3166
rect 23933 3090 23999 3093
rect 17174 3088 23999 3090
rect 17174 3032 23938 3088
rect 23994 3032 23999 3088
rect 17174 3030 23999 3032
rect 13077 2954 13143 2957
rect 15012 2954 15072 3030
rect 16205 3027 16271 3030
rect 23933 3027 23999 3030
rect 13077 2952 15072 2954
rect 13077 2896 13082 2952
rect 13138 2896 15072 2952
rect 13077 2894 15072 2896
rect 15193 2954 15259 2957
rect 15745 2954 15811 2957
rect 15878 2954 15884 2956
rect 15193 2952 15884 2954
rect 15193 2896 15198 2952
rect 15254 2896 15750 2952
rect 15806 2896 15884 2952
rect 15193 2894 15884 2896
rect 13077 2891 13143 2894
rect 15193 2891 15259 2894
rect 15745 2891 15811 2894
rect 15878 2892 15884 2894
rect 15948 2892 15954 2956
rect 200 2758 2790 2818
rect 7649 2818 7715 2821
rect 9254 2818 9260 2820
rect 7649 2816 9260 2818
rect 7649 2760 7654 2816
rect 7710 2760 9260 2816
rect 7649 2758 9260 2760
rect 200 2728 800 2758
rect 7649 2755 7715 2758
rect 9254 2756 9260 2758
rect 9324 2756 9330 2820
rect 10225 2818 10291 2821
rect 22093 2818 22159 2821
rect 10225 2816 22159 2818
rect 10225 2760 10230 2816
rect 10286 2760 22098 2816
rect 22154 2760 22159 2816
rect 10225 2758 22159 2760
rect 10225 2755 10291 2758
rect 22093 2755 22159 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 13537 2682 13603 2685
rect 20805 2682 20871 2685
rect 13537 2680 20871 2682
rect 13537 2624 13542 2680
rect 13598 2624 20810 2680
rect 20866 2624 20871 2680
rect 13537 2622 20871 2624
rect 13537 2619 13603 2622
rect 20805 2619 20871 2622
rect 7833 2546 7899 2549
rect 22737 2546 22803 2549
rect 7833 2544 22803 2546
rect 7833 2488 7838 2544
rect 7894 2488 22742 2544
rect 22798 2488 22803 2544
rect 7833 2486 22803 2488
rect 7833 2483 7899 2486
rect 22737 2483 22803 2486
rect 6821 2410 6887 2413
rect 22185 2410 22251 2413
rect 6821 2408 22251 2410
rect 6821 2352 6826 2408
rect 6882 2352 22190 2408
rect 22246 2352 22251 2408
rect 6821 2350 22251 2352
rect 6821 2347 6887 2350
rect 22185 2347 22251 2350
rect 1945 2274 2011 2277
rect 15837 2274 15903 2277
rect 1945 2272 15903 2274
rect 1945 2216 1950 2272
rect 2006 2216 15842 2272
rect 15898 2216 15903 2272
rect 1945 2214 15903 2216
rect 1945 2211 2011 2214
rect 15837 2211 15903 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 9489 2138 9555 2141
rect 19425 2138 19491 2141
rect 9489 2136 19491 2138
rect 9489 2080 9494 2136
rect 9550 2080 19430 2136
rect 19486 2080 19491 2136
rect 9489 2078 19491 2080
rect 9489 2075 9555 2078
rect 19425 2075 19491 2078
rect 38193 2138 38259 2141
rect 39200 2138 39800 2168
rect 38193 2136 39800 2138
rect 38193 2080 38198 2136
rect 38254 2080 39800 2136
rect 38193 2078 39800 2080
rect 38193 2075 38259 2078
rect 39200 2048 39800 2078
rect 200 1458 800 1488
rect 23565 1458 23631 1461
rect 200 1456 23631 1458
rect 200 1400 23570 1456
rect 23626 1400 23631 1456
rect 200 1398 23631 1400
rect 200 1368 800 1398
rect 23565 1395 23631 1398
rect 5165 1322 5231 1325
rect 22277 1322 22343 1325
rect 5165 1320 22343 1322
rect 5165 1264 5170 1320
rect 5226 1264 22282 1320
rect 22338 1264 22343 1320
rect 5165 1262 22343 1264
rect 5165 1259 5231 1262
rect 22277 1259 22343 1262
rect 37273 98 37339 101
rect 39200 98 39800 128
rect 37273 96 39800 98
rect 37273 40 37278 96
rect 37334 40 39800 96
rect 37273 38 39800 40
rect 37273 35 37339 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 7604 36484 7668 36548
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 3924 29004 3988 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 12020 23564 12084 23628
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 10548 21448 10612 21452
rect 10548 21392 10562 21448
rect 10562 21392 10612 21448
rect 10548 21388 10612 21392
rect 5764 21252 5828 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 9444 19348 9508 19412
rect 5948 19212 6012 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 15884 17172 15948 17236
rect 15332 17036 15396 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 2636 16824 2700 16828
rect 2636 16768 2686 16824
rect 2686 16768 2700 16824
rect 2636 16764 2700 16768
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4660 15948 4724 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 2452 15404 2516 15468
rect 3188 15328 3252 15332
rect 3188 15272 3238 15328
rect 3238 15272 3252 15328
rect 3188 15268 3252 15272
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 9260 14452 9324 14516
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 8156 13636 8220 13700
rect 11284 13636 11348 13700
rect 16068 13636 16132 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 9628 13500 9692 13564
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 5212 13016 5276 13020
rect 5212 12960 5262 13016
rect 5262 12960 5276 13016
rect 5212 12956 5276 12960
rect 5396 12548 5460 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 5212 12276 5276 12340
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 3924 11868 3988 11932
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 2636 11112 2700 11116
rect 2636 11056 2686 11112
rect 2686 11056 2700 11112
rect 2636 11052 2700 11056
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 2452 10644 2516 10708
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4660 10100 4724 10164
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 3188 9692 3252 9756
rect 7604 9556 7668 9620
rect 9076 9284 9140 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 5764 9208 5828 9212
rect 5764 9152 5778 9208
rect 5778 9152 5828 9208
rect 5764 9148 5828 9152
rect 10548 8876 10612 8940
rect 12020 8800 12084 8804
rect 12020 8744 12034 8800
rect 12034 8744 12084 8800
rect 12020 8740 12084 8744
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 9628 8196 9692 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 8156 8060 8220 8124
rect 9076 7924 9140 7988
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 11284 7108 11348 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 15332 6896 15396 6900
rect 15332 6840 15346 6896
rect 15346 6840 15396 6896
rect 15332 6836 15396 6840
rect 19380 6564 19444 6628
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 19380 6080 19444 6084
rect 19380 6024 19430 6080
rect 19430 6024 19444 6080
rect 19380 6020 19444 6024
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 9444 5612 9508 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 5396 5068 5460 5132
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 5948 4040 6012 4044
rect 5948 3984 5962 4040
rect 5962 3984 6012 4040
rect 5948 3980 6012 3984
rect 9260 3980 9324 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 16068 3768 16132 3772
rect 16068 3712 16082 3768
rect 16082 3712 16132 3768
rect 16068 3708 16132 3712
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 15884 2892 15948 2956
rect 9260 2756 9324 2820
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 7603 36548 7669 36549
rect 7603 36484 7604 36548
rect 7668 36484 7669 36548
rect 7603 36483 7669 36484
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 3923 29068 3989 29069
rect 3923 29004 3924 29068
rect 3988 29004 3989 29068
rect 3923 29003 3989 29004
rect 2635 16828 2701 16829
rect 2635 16764 2636 16828
rect 2700 16764 2701 16828
rect 2635 16763 2701 16764
rect 2451 15468 2517 15469
rect 2451 15404 2452 15468
rect 2516 15404 2517 15468
rect 2451 15403 2517 15404
rect 2454 10709 2514 15403
rect 2638 11117 2698 16763
rect 3187 15332 3253 15333
rect 3187 15268 3188 15332
rect 3252 15268 3253 15332
rect 3187 15267 3253 15268
rect 2635 11116 2701 11117
rect 2635 11052 2636 11116
rect 2700 11052 2701 11116
rect 2635 11051 2701 11052
rect 2451 10708 2517 10709
rect 2451 10644 2452 10708
rect 2516 10644 2517 10708
rect 2451 10643 2517 10644
rect 3190 9757 3250 15267
rect 3926 11933 3986 29003
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 5763 21316 5829 21317
rect 5763 21252 5764 21316
rect 5828 21252 5829 21316
rect 5763 21251 5829 21252
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4659 16012 4725 16013
rect 4659 15948 4660 16012
rect 4724 15948 4725 16012
rect 4659 15947 4725 15948
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 3923 11932 3989 11933
rect 3923 11868 3924 11932
rect 3988 11868 3989 11932
rect 3923 11867 3989 11868
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3187 9756 3253 9757
rect 3187 9692 3188 9756
rect 3252 9692 3253 9756
rect 3187 9691 3253 9692
rect 4208 9280 4528 10304
rect 4662 10165 4722 15947
rect 5211 13020 5277 13021
rect 5211 12956 5212 13020
rect 5276 12956 5277 13020
rect 5211 12955 5277 12956
rect 5214 12341 5274 12955
rect 5395 12612 5461 12613
rect 5395 12548 5396 12612
rect 5460 12548 5461 12612
rect 5395 12547 5461 12548
rect 5211 12340 5277 12341
rect 5211 12276 5212 12340
rect 5276 12276 5277 12340
rect 5211 12275 5277 12276
rect 4659 10164 4725 10165
rect 4659 10100 4660 10164
rect 4724 10100 4725 10164
rect 4659 10099 4725 10100
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 5398 5133 5458 12547
rect 5766 9213 5826 21251
rect 5947 19276 6013 19277
rect 5947 19212 5948 19276
rect 6012 19212 6013 19276
rect 5947 19211 6013 19212
rect 5763 9212 5829 9213
rect 5763 9148 5764 9212
rect 5828 9148 5829 9212
rect 5763 9147 5829 9148
rect 5395 5132 5461 5133
rect 5395 5068 5396 5132
rect 5460 5068 5461 5132
rect 5395 5067 5461 5068
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 5950 4045 6010 19211
rect 7606 9621 7666 36483
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 12019 23628 12085 23629
rect 12019 23564 12020 23628
rect 12084 23564 12085 23628
rect 12019 23563 12085 23564
rect 10547 21452 10613 21453
rect 10547 21388 10548 21452
rect 10612 21388 10613 21452
rect 10547 21387 10613 21388
rect 9443 19412 9509 19413
rect 9443 19348 9444 19412
rect 9508 19348 9509 19412
rect 9443 19347 9509 19348
rect 9259 14516 9325 14517
rect 9259 14452 9260 14516
rect 9324 14452 9325 14516
rect 9259 14451 9325 14452
rect 8155 13700 8221 13701
rect 8155 13636 8156 13700
rect 8220 13636 8221 13700
rect 8155 13635 8221 13636
rect 7603 9620 7669 9621
rect 7603 9556 7604 9620
rect 7668 9556 7669 9620
rect 7603 9555 7669 9556
rect 8158 8125 8218 13635
rect 9075 9348 9141 9349
rect 9075 9284 9076 9348
rect 9140 9284 9141 9348
rect 9075 9283 9141 9284
rect 8155 8124 8221 8125
rect 8155 8060 8156 8124
rect 8220 8060 8221 8124
rect 8155 8059 8221 8060
rect 9078 7989 9138 9283
rect 9075 7988 9141 7989
rect 9075 7924 9076 7988
rect 9140 7924 9141 7988
rect 9075 7923 9141 7924
rect 9262 4045 9322 14451
rect 9446 5677 9506 19347
rect 9627 13564 9693 13565
rect 9627 13500 9628 13564
rect 9692 13500 9693 13564
rect 9627 13499 9693 13500
rect 9630 8261 9690 13499
rect 10550 8941 10610 21387
rect 11283 13700 11349 13701
rect 11283 13636 11284 13700
rect 11348 13636 11349 13700
rect 11283 13635 11349 13636
rect 10547 8940 10613 8941
rect 10547 8876 10548 8940
rect 10612 8876 10613 8940
rect 10547 8875 10613 8876
rect 9627 8260 9693 8261
rect 9627 8196 9628 8260
rect 9692 8196 9693 8260
rect 9627 8195 9693 8196
rect 11286 7173 11346 13635
rect 12022 8805 12082 23563
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 15883 17236 15949 17237
rect 15883 17172 15884 17236
rect 15948 17172 15949 17236
rect 15883 17171 15949 17172
rect 15331 17100 15397 17101
rect 15331 17036 15332 17100
rect 15396 17036 15397 17100
rect 15331 17035 15397 17036
rect 12019 8804 12085 8805
rect 12019 8740 12020 8804
rect 12084 8740 12085 8804
rect 12019 8739 12085 8740
rect 11283 7172 11349 7173
rect 11283 7108 11284 7172
rect 11348 7108 11349 7172
rect 11283 7107 11349 7108
rect 15334 6901 15394 17035
rect 15331 6900 15397 6901
rect 15331 6836 15332 6900
rect 15396 6836 15397 6900
rect 15331 6835 15397 6836
rect 9443 5676 9509 5677
rect 9443 5612 9444 5676
rect 9508 5612 9509 5676
rect 9443 5611 9509 5612
rect 5947 4044 6013 4045
rect 5947 3980 5948 4044
rect 6012 3980 6013 4044
rect 5947 3979 6013 3980
rect 9259 4044 9325 4045
rect 9259 3980 9260 4044
rect 9324 3980 9325 4044
rect 9259 3979 9325 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 9262 2821 9322 3979
rect 15886 2957 15946 17171
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 16067 13700 16133 13701
rect 16067 13636 16068 13700
rect 16132 13636 16133 13700
rect 16067 13635 16133 13636
rect 16070 3773 16130 13635
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19379 6628 19445 6629
rect 19379 6564 19380 6628
rect 19444 6564 19445 6628
rect 19379 6563 19445 6564
rect 19382 6085 19442 6563
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19379 6084 19445 6085
rect 19379 6020 19380 6084
rect 19444 6020 19445 6084
rect 19379 6019 19445 6020
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 16067 3772 16133 3773
rect 16067 3708 16068 3772
rect 16132 3708 16133 3772
rect 16067 3707 16133 3708
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 15883 2956 15949 2957
rect 15883 2892 15884 2956
rect 15948 2892 15949 2956
rect 15883 2891 15949 2892
rect 9259 2820 9325 2821
rect 9259 2756 9260 2820
rect 9324 2756 9325 2820
rect 9259 2755 9325 2756
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23552 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 23736 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform 1 0 22080 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1667941163
transform 1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1667941163
transform 1 0 13064 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1667941163
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1667941163
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_181 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1667941163
transform 1 0 20240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_212
timestamp 1667941163
transform 1 0 20608 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1667941163
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_258 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 1667941163
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_294
timestamp 1667941163
transform 1 0 28152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1667941163
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_322
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1667941163
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_342
timestamp 1667941163
transform 1 0 32568 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 1667941163
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1667941163
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 1667941163
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_399
timestamp 1667941163
transform 1 0 37812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_26
timestamp 1667941163
transform 1 0 3496 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_32
timestamp 1667941163
transform 1 0 4048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_65
timestamp 1667941163
transform 1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1667941163
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_97
timestamp 1667941163
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1667941163
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1667941163
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1667941163
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1667941163
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1667941163
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1667941163
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1667941163
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1667941163
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_242
timestamp 1667941163
transform 1 0 23368 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_246
timestamp 1667941163
transform 1 0 23736 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_251
timestamp 1667941163
transform 1 0 24196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_263
timestamp 1667941163
transform 1 0 25300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp 1667941163
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1667941163
transform 1 0 2208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1667941163
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_47
timestamp 1667941163
transform 1 0 5428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1667941163
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_114
timestamp 1667941163
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1667941163
transform 1 0 16192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_171
timestamp 1667941163
transform 1 0 16836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178
timestamp 1667941163
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1667941163
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1667941163
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_216
timestamp 1667941163
transform 1 0 20976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_223
timestamp 1667941163
transform 1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_227
timestamp 1667941163
transform 1 0 21988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_230
timestamp 1667941163
transform 1 0 22264 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_238
timestamp 1667941163
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_244
timestamp 1667941163
transform 1 0 23552 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1667941163
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_280
timestamp 1667941163
transform 1 0 26864 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_292
timestamp 1667941163
transform 1 0 27968 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1667941163
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1667941163
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_14
timestamp 1667941163
transform 1 0 2392 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_26
timestamp 1667941163
transform 1 0 3496 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_32
timestamp 1667941163
transform 1 0 4048 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1667941163
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_68
timestamp 1667941163
transform 1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_95
timestamp 1667941163
transform 1 0 9844 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1667941163
transform 1 0 10212 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1667941163
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1667941163
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1667941163
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1667941163
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_177
timestamp 1667941163
transform 1 0 17388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1667941163
transform 1 0 18032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_191
timestamp 1667941163
transform 1 0 18676 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_198
timestamp 1667941163
transform 1 0 19320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1667941163
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1667941163
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1667941163
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_286
timestamp 1667941163
transform 1 0 27416 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_298
timestamp 1667941163
transform 1 0 28520 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_310
timestamp 1667941163
transform 1 0 29624 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_322
timestamp 1667941163
transform 1 0 30728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1667941163
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1667941163
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_14
timestamp 1667941163
transform 1 0 2392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_18
timestamp 1667941163
transform 1 0 2760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1667941163
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1667941163
transform 1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 1667941163
transform 1 0 6992 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1667941163
transform 1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_75
timestamp 1667941163
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_91
timestamp 1667941163
transform 1 0 9476 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_95
timestamp 1667941163
transform 1 0 9844 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1667941163
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_126
timestamp 1667941163
transform 1 0 12696 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_152
timestamp 1667941163
transform 1 0 15088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_159
timestamp 1667941163
transform 1 0 15732 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_166
timestamp 1667941163
transform 1 0 16376 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1667941163
transform 1 0 17020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_180
timestamp 1667941163
transform 1 0 17664 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1667941163
transform 1 0 18400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1667941163
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_202
timestamp 1667941163
transform 1 0 19688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_216
timestamp 1667941163
transform 1 0 20976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1667941163
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1667941163
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_237
timestamp 1667941163
transform 1 0 22908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1667941163
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_13
timestamp 1667941163
transform 1 0 2300 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1667941163
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_42
timestamp 1667941163
transform 1 0 4968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1667941163
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1667941163
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1667941163
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_136
timestamp 1667941163
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_156
timestamp 1667941163
transform 1 0 15456 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1667941163
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_174
timestamp 1667941163
transform 1 0 17112 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1667941163
transform 1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1667941163
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_202
timestamp 1667941163
transform 1 0 19688 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_209
timestamp 1667941163
transform 1 0 20332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1667941163
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_230
timestamp 1667941163
transform 1 0 22264 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_325
timestamp 1667941163
transform 1 0 31004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_342
timestamp 1667941163
transform 1 0 32568 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_354
timestamp 1667941163
transform 1 0 33672 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_366
timestamp 1667941163
transform 1 0 34776 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_378
timestamp 1667941163
transform 1 0 35880 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1667941163
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_398
timestamp 1667941163
transform 1 0 37720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_37
timestamp 1667941163
transform 1 0 4508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1667941163
transform 1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_73
timestamp 1667941163
transform 1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1667941163
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_91
timestamp 1667941163
transform 1 0 9476 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_98
timestamp 1667941163
transform 1 0 10120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_125
timestamp 1667941163
transform 1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1667941163
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1667941163
transform 1 0 16744 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_184
timestamp 1667941163
transform 1 0 18032 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1667941163
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_202
timestamp 1667941163
transform 1 0 19688 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_216
timestamp 1667941163
transform 1 0 20976 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1667941163
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_230
timestamp 1667941163
transform 1 0 22264 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_242
timestamp 1667941163
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1667941163
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_258
timestamp 1667941163
transform 1 0 24840 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_270
timestamp 1667941163
transform 1 0 25944 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_282
timestamp 1667941163
transform 1 0 27048 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_294
timestamp 1667941163
transform 1 0 28152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1667941163
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_371
timestamp 1667941163
transform 1 0 35236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_383
timestamp 1667941163
transform 1 0 36340 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_395
timestamp 1667941163
transform 1 0 37444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33
timestamp 1667941163
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_40
timestamp 1667941163
transform 1 0 4784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_47
timestamp 1667941163
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1667941163
transform 1 0 6808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp 1667941163
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_99
timestamp 1667941163
transform 1 0 10212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1667941163
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_135
timestamp 1667941163
transform 1 0 13524 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_159
timestamp 1667941163
transform 1 0 15732 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_180
timestamp 1667941163
transform 1 0 17664 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_187
timestamp 1667941163
transform 1 0 18308 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_194
timestamp 1667941163
transform 1 0 18952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1667941163
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1667941163
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1667941163
transform 1 0 20884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_229
timestamp 1667941163
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_233
timestamp 1667941163
transform 1 0 22540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_245
timestamp 1667941163
transform 1 0 23644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_257
timestamp 1667941163
transform 1 0 24748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1667941163
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1667941163
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_312
timestamp 1667941163
transform 1 0 29808 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_324
timestamp 1667941163
transform 1 0 30912 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_54
timestamp 1667941163
transform 1 0 6072 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_96
timestamp 1667941163
transform 1 0 9936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_129
timestamp 1667941163
transform 1 0 12972 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_151
timestamp 1667941163
transform 1 0 14996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_159
timestamp 1667941163
transform 1 0 15732 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_168
timestamp 1667941163
transform 1 0 16560 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_175
timestamp 1667941163
transform 1 0 17204 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_182
timestamp 1667941163
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_202
timestamp 1667941163
transform 1 0 19688 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_206
timestamp 1667941163
transform 1 0 20056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1667941163
transform 1 0 20424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_222
timestamp 1667941163
transform 1 0 21528 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_230
timestamp 1667941163
transform 1 0 22264 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_235
timestamp 1667941163
transform 1 0 22724 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp 1667941163
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_337
timestamp 1667941163
transform 1 0 32108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_349
timestamp 1667941163
transform 1 0 33212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1667941163
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_25
timestamp 1667941163
transform 1 0 3404 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1667941163
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1667941163
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_70
timestamp 1667941163
transform 1 0 7544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_97
timestamp 1667941163
transform 1 0 10028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1667941163
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1667941163
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_148
timestamp 1667941163
transform 1 0 14720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_156
timestamp 1667941163
transform 1 0 15456 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1667941163
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp 1667941163
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_188
timestamp 1667941163
transform 1 0 18400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_195
timestamp 1667941163
transform 1 0 19044 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_202
timestamp 1667941163
transform 1 0 19688 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_210
timestamp 1667941163
transform 1 0 20424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_214
timestamp 1667941163
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_236
timestamp 1667941163
transform 1 0 22816 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_311
timestamp 1667941163
transform 1 0 29716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_323
timestamp 1667941163
transform 1 0 30820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_358
timestamp 1667941163
transform 1 0 34040 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_370
timestamp 1667941163
transform 1 0 35144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_382
timestamp 1667941163
transform 1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1667941163
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_401
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_47
timestamp 1667941163
transform 1 0 5428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_69
timestamp 1667941163
transform 1 0 7452 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1667941163
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1667941163
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_118
timestamp 1667941163
transform 1 0 11960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1667941163
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_129
timestamp 1667941163
transform 1 0 12972 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1667941163
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_151
timestamp 1667941163
transform 1 0 14996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1667941163
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1667941163
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_173
timestamp 1667941163
transform 1 0 17020 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1667941163
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1667941163
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_213
timestamp 1667941163
transform 1 0 20700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_225
timestamp 1667941163
transform 1 0 21804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_229
timestamp 1667941163
transform 1 0 22172 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_236
timestamp 1667941163
transform 1 0 22816 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1667941163
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_292
timestamp 1667941163
transform 1 0 27968 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1667941163
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_32
timestamp 1667941163
transform 1 0 4048 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1667941163
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_47
timestamp 1667941163
transform 1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_63
timestamp 1667941163
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_84
timestamp 1667941163
transform 1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1667941163
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1667941163
transform 1 0 13524 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_146
timestamp 1667941163
transform 1 0 14536 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1667941163
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1667941163
transform 1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_191
timestamp 1667941163
transform 1 0 18676 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_203
timestamp 1667941163
transform 1 0 19780 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1667941163
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1667941163
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_298
timestamp 1667941163
transform 1 0 28520 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_310
timestamp 1667941163
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_322
timestamp 1667941163
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1667941163
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_52
timestamp 1667941163
transform 1 0 5888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1667941163
transform 1 0 6624 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1667941163
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1667941163
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_117
timestamp 1667941163
transform 1 0 11868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_126
timestamp 1667941163
transform 1 0 12696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1667941163
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_151
timestamp 1667941163
transform 1 0 14996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_158
timestamp 1667941163
transform 1 0 15640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_170
timestamp 1667941163
transform 1 0 16744 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_176
timestamp 1667941163
transform 1 0 17296 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_180
timestamp 1667941163
transform 1 0 17664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1667941163
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_220
timestamp 1667941163
transform 1 0 21344 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1667941163
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_261
timestamp 1667941163
transform 1 0 25116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_273
timestamp 1667941163
transform 1 0 26220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_285
timestamp 1667941163
transform 1 0 27324 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_297
timestamp 1667941163
transform 1 0 28428 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_305
timestamp 1667941163
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1667941163
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1667941163
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_85
timestamp 1667941163
transform 1 0 8924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1667941163
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1667941163
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1667941163
transform 1 0 12420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_130
timestamp 1667941163
transform 1 0 13064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_144
timestamp 1667941163
transform 1 0 14352 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1667941163
transform 1 0 15180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_180
timestamp 1667941163
transform 1 0 17664 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_186
timestamp 1667941163
transform 1 0 18216 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_190
timestamp 1667941163
transform 1 0 18584 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_202
timestamp 1667941163
transform 1 0 19688 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp 1667941163
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_243
timestamp 1667941163
transform 1 0 23460 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_255
timestamp 1667941163
transform 1 0 24564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_267
timestamp 1667941163
transform 1 0 25668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_39
timestamp 1667941163
transform 1 0 4692 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp 1667941163
transform 1 0 5520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_72
timestamp 1667941163
transform 1 0 7728 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_78
timestamp 1667941163
transform 1 0 8280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_94
timestamp 1667941163
transform 1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_118
timestamp 1667941163
transform 1 0 11960 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1667941163
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1667941163
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_151
timestamp 1667941163
transform 1 0 14996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_157
timestamp 1667941163
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_161
timestamp 1667941163
transform 1 0 15916 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_168
timestamp 1667941163
transform 1 0 16560 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_181
timestamp 1667941163
transform 1 0 17756 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1667941163
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1667941163
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_210
timestamp 1667941163
transform 1 0 20424 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_222
timestamp 1667941163
transform 1 0 21528 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_234
timestamp 1667941163
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_238
timestamp 1667941163
transform 1 0 23000 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1667941163
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_353
timestamp 1667941163
transform 1 0 33580 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1667941163
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_8
timestamp 1667941163
transform 1 0 1840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_40
timestamp 1667941163
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1667941163
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_89
timestamp 1667941163
transform 1 0 9292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_135
timestamp 1667941163
transform 1 0 13524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_141
timestamp 1667941163
transform 1 0 14076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1667941163
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1667941163
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1667941163
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_179
timestamp 1667941163
transform 1 0 17572 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1667941163
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_194
timestamp 1667941163
transform 1 0 18952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_198
timestamp 1667941163
transform 1 0 19320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_202
timestamp 1667941163
transform 1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_206
timestamp 1667941163
transform 1 0 20056 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_210
timestamp 1667941163
transform 1 0 20424 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_233
timestamp 1667941163
transform 1 0 22540 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_241
timestamp 1667941163
transform 1 0 23276 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_245
timestamp 1667941163
transform 1 0 23644 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_252
timestamp 1667941163
transform 1 0 24288 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_264
timestamp 1667941163
transform 1 0 25392 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1667941163
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_286
timestamp 1667941163
transform 1 0 27416 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_298
timestamp 1667941163
transform 1 0 28520 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_310
timestamp 1667941163
transform 1 0 29624 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_322
timestamp 1667941163
transform 1 0 30728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1667941163
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_370
timestamp 1667941163
transform 1 0 35144 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1667941163
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_54
timestamp 1667941163
transform 1 0 6072 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_94
timestamp 1667941163
transform 1 0 9752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1667941163
transform 1 0 11960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp 1667941163
transform 1 0 12696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_152
timestamp 1667941163
transform 1 0 15088 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1667941163
transform 1 0 16100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1667941163
transform 1 0 17204 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_179
timestamp 1667941163
transform 1 0 17572 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1667941163
transform 1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_187
timestamp 1667941163
transform 1 0 18308 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1667941163
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1667941163
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_206
timestamp 1667941163
transform 1 0 20056 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1667941163
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_222
timestamp 1667941163
transform 1 0 21528 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_237
timestamp 1667941163
transform 1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1667941163
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_258
timestamp 1667941163
transform 1 0 24840 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_270
timestamp 1667941163
transform 1 0 25944 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_282
timestamp 1667941163
transform 1 0 27048 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_294
timestamp 1667941163
transform 1 0 28152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1667941163
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_314
timestamp 1667941163
transform 1 0 29992 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_326
timestamp 1667941163
transform 1 0 31096 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_338
timestamp 1667941163
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_350
timestamp 1667941163
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1667941163
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1667941163
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_34
timestamp 1667941163
transform 1 0 4232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_46
timestamp 1667941163
transform 1 0 5336 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_50
timestamp 1667941163
transform 1 0 5704 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_67
timestamp 1667941163
transform 1 0 7268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_74
timestamp 1667941163
transform 1 0 7912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1667941163
transform 1 0 10120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1667941163
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1667941163
transform 1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_146
timestamp 1667941163
transform 1 0 14536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1667941163
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1667941163
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1667941163
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_182
timestamp 1667941163
transform 1 0 17848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1667941163
transform 1 0 18492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1667941163
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_213
timestamp 1667941163
transform 1 0 20700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1667941163
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_230
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_252
timestamp 1667941163
transform 1 0 24288 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_259
timestamp 1667941163
transform 1 0 24932 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_266
timestamp 1667941163
transform 1 0 25576 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1667941163
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_357
timestamp 1667941163
transform 1 0 33948 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_363
timestamp 1667941163
transform 1 0 34500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_375
timestamp 1667941163
transform 1 0 35604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_387
timestamp 1667941163
transform 1 0 36708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_401
timestamp 1667941163
transform 1 0 37996 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1667941163
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_43
timestamp 1667941163
transform 1 0 5060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_67
timestamp 1667941163
transform 1 0 7268 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_96
timestamp 1667941163
transform 1 0 9936 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_104
timestamp 1667941163
transform 1 0 10672 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1667941163
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1667941163
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1667941163
transform 1 0 14720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1667941163
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_173
timestamp 1667941163
transform 1 0 17020 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_179
timestamp 1667941163
transform 1 0 17572 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_183
timestamp 1667941163
transform 1 0 17940 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1667941163
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_204
timestamp 1667941163
transform 1 0 19872 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1667941163
transform 1 0 21160 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_225
timestamp 1667941163
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_232
timestamp 1667941163
transform 1 0 22448 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_240
timestamp 1667941163
transform 1 0 23184 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1667941163
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_263
timestamp 1667941163
transform 1 0 25300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_275
timestamp 1667941163
transform 1 0 26404 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_287
timestamp 1667941163
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_299
timestamp 1667941163
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_376
timestamp 1667941163
transform 1 0 35696 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_388
timestamp 1667941163
transform 1 0 36800 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_400
timestamp 1667941163
transform 1 0 37904 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1667941163
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_26
timestamp 1667941163
transform 1 0 3496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1667941163
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_67
timestamp 1667941163
transform 1 0 7268 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1667941163
transform 1 0 8280 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_90
timestamp 1667941163
transform 1 0 9384 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 1667941163
transform 1 0 10120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_103
timestamp 1667941163
transform 1 0 10580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1667941163
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_119
timestamp 1667941163
transform 1 0 12052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1667941163
transform 1 0 13248 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_136
timestamp 1667941163
transform 1 0 13616 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1667941163
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_152
timestamp 1667941163
transform 1 0 15088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_156
timestamp 1667941163
transform 1 0 15456 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1667941163
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1667941163
transform 1 0 17572 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_183
timestamp 1667941163
transform 1 0 17940 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1667941163
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_191
timestamp 1667941163
transform 1 0 18676 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1667941163
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1667941163
transform 1 0 20148 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_214
timestamp 1667941163
transform 1 0 20792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_218
timestamp 1667941163
transform 1 0 21160 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_230
timestamp 1667941163
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_247
timestamp 1667941163
transform 1 0 23828 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_254
timestamp 1667941163
transform 1 0 24472 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_266
timestamp 1667941163
transform 1 0 25576 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1667941163
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1667941163
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1667941163
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_38
timestamp 1667941163
transform 1 0 4600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_62
timestamp 1667941163
transform 1 0 6808 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_71
timestamp 1667941163
transform 1 0 7636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1667941163
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_92
timestamp 1667941163
transform 1 0 9568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1667941163
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1667941163
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_113
timestamp 1667941163
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_125
timestamp 1667941163
transform 1 0 12604 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_147
timestamp 1667941163
transform 1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_154
timestamp 1667941163
transform 1 0 15272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_166
timestamp 1667941163
transform 1 0 16376 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_172
timestamp 1667941163
transform 1 0 16928 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1667941163
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_185
timestamp 1667941163
transform 1 0 18124 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1667941163
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1667941163
transform 1 0 20884 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_223
timestamp 1667941163
transform 1 0 21620 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1667941163
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_240
timestamp 1667941163
transform 1 0 23184 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1667941163
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_349
timestamp 1667941163
transform 1 0 33212 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_353
timestamp 1667941163
transform 1 0 33580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1667941163
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1667941163
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_29
timestamp 1667941163
transform 1 0 3772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_38
timestamp 1667941163
transform 1 0 4600 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_45
timestamp 1667941163
transform 1 0 5244 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1667941163
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_65
timestamp 1667941163
transform 1 0 7084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1667941163
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_79
timestamp 1667941163
transform 1 0 8372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_85
timestamp 1667941163
transform 1 0 8924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_89
timestamp 1667941163
transform 1 0 9292 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1667941163
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1667941163
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 1667941163
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_134
timestamp 1667941163
transform 1 0 13432 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_148
timestamp 1667941163
transform 1 0 14720 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1667941163
transform 1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_194
timestamp 1667941163
transform 1 0 18952 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_202
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_206
timestamp 1667941163
transform 1 0 20056 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_235
timestamp 1667941163
transform 1 0 22724 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1667941163
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_254
timestamp 1667941163
transform 1 0 24472 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_266
timestamp 1667941163
transform 1 0 25576 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1667941163
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_18
timestamp 1667941163
transform 1 0 2760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_22
timestamp 1667941163
transform 1 0 3128 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_39
timestamp 1667941163
transform 1 0 4692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_43
timestamp 1667941163
transform 1 0 5060 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_59
timestamp 1667941163
transform 1 0 6532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_63
timestamp 1667941163
transform 1 0 6900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_70
timestamp 1667941163
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_96
timestamp 1667941163
transform 1 0 9936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1667941163
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_110
timestamp 1667941163
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1667941163
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1667941163
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1667941163
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1667941163
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_160
timestamp 1667941163
transform 1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_173
timestamp 1667941163
transform 1 0 17020 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_182
timestamp 1667941163
transform 1 0 17848 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_216
timestamp 1667941163
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_220
timestamp 1667941163
transform 1 0 21344 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_229
timestamp 1667941163
transform 1 0 22172 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_236
timestamp 1667941163
transform 1 0 22816 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1667941163
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_295
timestamp 1667941163
transform 1 0 28244 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1667941163
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1667941163
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1667941163
transform 1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1667941163
transform 1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_25
timestamp 1667941163
transform 1 0 3404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_32
timestamp 1667941163
transform 1 0 4048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_46
timestamp 1667941163
transform 1 0 5336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1667941163
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1667941163
transform 1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1667941163
transform 1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_83
timestamp 1667941163
transform 1 0 8740 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_87
timestamp 1667941163
transform 1 0 9108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_96
timestamp 1667941163
transform 1 0 9936 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1667941163
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1667941163
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_128
timestamp 1667941163
transform 1 0 12880 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1667941163
transform 1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_148
timestamp 1667941163
transform 1 0 14720 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1667941163
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1667941163
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_183
timestamp 1667941163
transform 1 0 17940 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_187
timestamp 1667941163
transform 1 0 18308 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1667941163
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_208
timestamp 1667941163
transform 1 0 20240 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_216
timestamp 1667941163
transform 1 0 20976 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1667941163
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1667941163
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_242
timestamp 1667941163
transform 1 0 23368 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_254
timestamp 1667941163
transform 1 0 24472 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_266
timestamp 1667941163
transform 1 0 25576 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_8
timestamp 1667941163
transform 1 0 1840 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_17
timestamp 1667941163
transform 1 0 2668 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1667941163
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1667941163
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_47
timestamp 1667941163
transform 1 0 5428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_58
timestamp 1667941163
transform 1 0 6440 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1667941163
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_91
timestamp 1667941163
transform 1 0 9476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_98
timestamp 1667941163
transform 1 0 10120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_110
timestamp 1667941163
transform 1 0 11224 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_126
timestamp 1667941163
transform 1 0 12696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1667941163
transform 1 0 14720 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_160
timestamp 1667941163
transform 1 0 15824 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_166
timestamp 1667941163
transform 1 0 16376 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_175
timestamp 1667941163
transform 1 0 17204 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_183
timestamp 1667941163
transform 1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1667941163
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_212
timestamp 1667941163
transform 1 0 20608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_216
timestamp 1667941163
transform 1 0 20976 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_225
timestamp 1667941163
transform 1 0 21804 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_232
timestamp 1667941163
transform 1 0 22448 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_239
timestamp 1667941163
transform 1 0 23092 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1667941163
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_372
timestamp 1667941163
transform 1 0 35328 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_384
timestamp 1667941163
transform 1 0 36432 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_396
timestamp 1667941163
transform 1 0 37536 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_10
timestamp 1667941163
transform 1 0 2024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_14
timestamp 1667941163
transform 1 0 2392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_18
timestamp 1667941163
transform 1 0 2760 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_25
timestamp 1667941163
transform 1 0 3404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1667941163
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1667941163
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_63
timestamp 1667941163
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_67
timestamp 1667941163
transform 1 0 7268 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_74
timestamp 1667941163
transform 1 0 7912 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_87
timestamp 1667941163
transform 1 0 9108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1667941163
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_100
timestamp 1667941163
transform 1 0 10304 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1667941163
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1667941163
transform 1 0 12420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_128
timestamp 1667941163
transform 1 0 12880 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1667941163
transform 1 0 13248 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_142
timestamp 1667941163
transform 1 0 14168 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_148
timestamp 1667941163
transform 1 0 14720 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1667941163
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1667941163
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_179
timestamp 1667941163
transform 1 0 17572 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_187
timestamp 1667941163
transform 1 0 18308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_202
timestamp 1667941163
transform 1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_214
timestamp 1667941163
transform 1 0 20792 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1667941163
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1667941163
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1667941163
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_250
timestamp 1667941163
transform 1 0 24104 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_262
timestamp 1667941163
transform 1 0 25208 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1667941163
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_357
timestamp 1667941163
transform 1 0 33948 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_362
timestamp 1667941163
transform 1 0 34408 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_374
timestamp 1667941163
transform 1 0 35512 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_386
timestamp 1667941163
transform 1 0 36616 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_9
timestamp 1667941163
transform 1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_16
timestamp 1667941163
transform 1 0 2576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1667941163
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_34
timestamp 1667941163
transform 1 0 4232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1667941163
transform 1 0 4600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_42
timestamp 1667941163
transform 1 0 4968 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_48
timestamp 1667941163
transform 1 0 5520 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_52
timestamp 1667941163
transform 1 0 5888 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_64
timestamp 1667941163
transform 1 0 6992 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_72
timestamp 1667941163
transform 1 0 7728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1667941163
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_95
timestamp 1667941163
transform 1 0 9844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_99
timestamp 1667941163
transform 1 0 10212 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_103
timestamp 1667941163
transform 1 0 10580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_110
timestamp 1667941163
transform 1 0 11224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1667941163
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1667941163
transform 1 0 12512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_131
timestamp 1667941163
transform 1 0 13156 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1667941163
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_151
timestamp 1667941163
transform 1 0 14996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_164
timestamp 1667941163
transform 1 0 16192 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1667941163
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_208
timestamp 1667941163
transform 1 0 20240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1667941163
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_232
timestamp 1667941163
transform 1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_239
timestamp 1667941163
transform 1 0 23092 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1667941163
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1667941163
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_11
timestamp 1667941163
transform 1 0 2116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_19
timestamp 1667941163
transform 1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_26
timestamp 1667941163
transform 1 0 3496 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_34
timestamp 1667941163
transform 1 0 4232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_46
timestamp 1667941163
transform 1 0 5336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_50
timestamp 1667941163
transform 1 0 5704 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_64
timestamp 1667941163
transform 1 0 6992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1667941163
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1667941163
transform 1 0 8464 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1667941163
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_96
timestamp 1667941163
transform 1 0 9936 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_103
timestamp 1667941163
transform 1 0 10580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1667941163
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_131
timestamp 1667941163
transform 1 0 13156 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_138
timestamp 1667941163
transform 1 0 13800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_150
timestamp 1667941163
transform 1 0 14904 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1667941163
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_179
timestamp 1667941163
transform 1 0 17572 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_185
timestamp 1667941163
transform 1 0 18124 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_194
timestamp 1667941163
transform 1 0 18952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_206
timestamp 1667941163
transform 1 0 20056 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_214
timestamp 1667941163
transform 1 0 20792 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1667941163
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_235
timestamp 1667941163
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_242
timestamp 1667941163
transform 1 0 23368 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_256
timestamp 1667941163
transform 1 0 24656 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_268
timestamp 1667941163
transform 1 0 25760 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_10
timestamp 1667941163
transform 1 0 2024 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_17
timestamp 1667941163
transform 1 0 2668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1667941163
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_45
timestamp 1667941163
transform 1 0 5244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_57
timestamp 1667941163
transform 1 0 6348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1667941163
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1667941163
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1667941163
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_94
timestamp 1667941163
transform 1 0 9752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_107
timestamp 1667941163
transform 1 0 10948 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_115
timestamp 1667941163
transform 1 0 11684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_119
timestamp 1667941163
transform 1 0 12052 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_126
timestamp 1667941163
transform 1 0 12696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_150
timestamp 1667941163
transform 1 0 14904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1667941163
transform 1 0 16100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_175
timestamp 1667941163
transform 1 0 17204 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1667941163
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1667941163
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_211
timestamp 1667941163
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1667941163
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_225
timestamp 1667941163
transform 1 0 21804 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1667941163
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1667941163
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_329
timestamp 1667941163
transform 1 0 31372 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_351
timestamp 1667941163
transform 1 0 33396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1667941163
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1667941163
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_63
timestamp 1667941163
transform 1 0 6900 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_73
timestamp 1667941163
transform 1 0 7820 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1667941163
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_89
timestamp 1667941163
transform 1 0 9292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1667941163
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_103
timestamp 1667941163
transform 1 0 10580 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_119
timestamp 1667941163
transform 1 0 12052 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 1667941163
transform 1 0 12696 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_138
timestamp 1667941163
transform 1 0 13800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_145
timestamp 1667941163
transform 1 0 14444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1667941163
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1667941163
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_180
timestamp 1667941163
transform 1 0 17664 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_189
timestamp 1667941163
transform 1 0 18492 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_201
timestamp 1667941163
transform 1 0 19596 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1667941163
transform 1 0 20332 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1667941163
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_231
timestamp 1667941163
transform 1 0 22356 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_240
timestamp 1667941163
transform 1 0 23184 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1667941163
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_254
timestamp 1667941163
transform 1 0 24472 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_266
timestamp 1667941163
transform 1 0 25576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_69
timestamp 1667941163
transform 1 0 7452 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_99
timestamp 1667941163
transform 1 0 10212 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_108
timestamp 1667941163
transform 1 0 11040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1667941163
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_124
timestamp 1667941163
transform 1 0 12512 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1667941163
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_155
timestamp 1667941163
transform 1 0 15364 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_159
timestamp 1667941163
transform 1 0 15732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_166
timestamp 1667941163
transform 1 0 16376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1667941163
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_180
timestamp 1667941163
transform 1 0 17664 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_212
timestamp 1667941163
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_224
timestamp 1667941163
transform 1 0 21712 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1667941163
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_350
timestamp 1667941163
transform 1 0 33304 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1667941163
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_405
timestamp 1667941163
transform 1 0 38364 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_74
timestamp 1667941163
transform 1 0 7912 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_80
timestamp 1667941163
transform 1 0 8464 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_84
timestamp 1667941163
transform 1 0 8832 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_91
timestamp 1667941163
transform 1 0 9476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1667941163
transform 1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_127
timestamp 1667941163
transform 1 0 12788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_144
timestamp 1667941163
transform 1 0 14352 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_151
timestamp 1667941163
transform 1 0 14996 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1667941163
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1667941163
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_188
timestamp 1667941163
transform 1 0 18400 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_200
timestamp 1667941163
transform 1 0 19504 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_213
timestamp 1667941163
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1667941163
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_231
timestamp 1667941163
transform 1 0 22356 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_235
timestamp 1667941163
transform 1 0 22724 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_250
timestamp 1667941163
transform 1 0 24104 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_257
timestamp 1667941163
transform 1 0 24748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1667941163
transform 1 0 25852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1667941163
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_8
timestamp 1667941163
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1667941163
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 1667941163
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_75
timestamp 1667941163
transform 1 0 8004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_91
timestamp 1667941163
transform 1 0 9476 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_103
timestamp 1667941163
transform 1 0 10580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1667941163
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_117
timestamp 1667941163
transform 1 0 11868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_124
timestamp 1667941163
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_131
timestamp 1667941163
transform 1 0 13156 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1667941163
transform 1 0 14720 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_155
timestamp 1667941163
transform 1 0 15364 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_167
timestamp 1667941163
transform 1 0 16468 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_182
timestamp 1667941163
transform 1 0 17848 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_190
timestamp 1667941163
transform 1 0 18584 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_208
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_215
timestamp 1667941163
transform 1 0 20884 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1667941163
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_243
timestamp 1667941163
transform 1 0 23460 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1667941163
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_258
timestamp 1667941163
transform 1 0 24840 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1667941163
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1667941163
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_75
timestamp 1667941163
transform 1 0 8004 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1667941163
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_91
timestamp 1667941163
transform 1 0 9476 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_97
timestamp 1667941163
transform 1 0 10028 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1667941163
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1667941163
transform 1 0 11960 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_130
timestamp 1667941163
transform 1 0 13064 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_136
timestamp 1667941163
transform 1 0 13616 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_140
timestamp 1667941163
transform 1 0 13984 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_147
timestamp 1667941163
transform 1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1667941163
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_185
timestamp 1667941163
transform 1 0 18124 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_191
timestamp 1667941163
transform 1 0 18676 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_195
timestamp 1667941163
transform 1 0 19044 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_199
timestamp 1667941163
transform 1 0 19412 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_208
timestamp 1667941163
transform 1 0 20240 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1667941163
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_231
timestamp 1667941163
transform 1 0 22356 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1667941163
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_247
timestamp 1667941163
transform 1 0 23828 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_254
timestamp 1667941163
transform 1 0 24472 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_266
timestamp 1667941163
transform 1 0 25576 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_71
timestamp 1667941163
transform 1 0 7636 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_75
timestamp 1667941163
transform 1 0 8004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1667941163
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_100
timestamp 1667941163
transform 1 0 10304 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_108
timestamp 1667941163
transform 1 0 11040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_118
timestamp 1667941163
transform 1 0 11960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_126
timestamp 1667941163
transform 1 0 12696 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_131
timestamp 1667941163
transform 1 0 13156 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1667941163
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_167
timestamp 1667941163
transform 1 0 16468 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_174
timestamp 1667941163
transform 1 0 17112 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_186
timestamp 1667941163
transform 1 0 18216 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_190
timestamp 1667941163
transform 1 0 18584 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_207
timestamp 1667941163
transform 1 0 20148 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_214
timestamp 1667941163
transform 1 0 20792 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_222
timestamp 1667941163
transform 1 0 21528 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1667941163
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_241
timestamp 1667941163
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1667941163
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1667941163
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_41
timestamp 1667941163
transform 1 0 4876 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1667941163
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_75
timestamp 1667941163
transform 1 0 8004 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_79
timestamp 1667941163
transform 1 0 8372 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_86
timestamp 1667941163
transform 1 0 9016 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_92
timestamp 1667941163
transform 1 0 9568 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_96
timestamp 1667941163
transform 1 0 9936 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_103
timestamp 1667941163
transform 1 0 10580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_123
timestamp 1667941163
transform 1 0 12420 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_139
timestamp 1667941163
transform 1 0 13892 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_146
timestamp 1667941163
transform 1 0 14536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_153
timestamp 1667941163
transform 1 0 15180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1667941163
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1667941163
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_177
timestamp 1667941163
transform 1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_184
timestamp 1667941163
transform 1 0 18032 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1667941163
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_208
timestamp 1667941163
transform 1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_215
timestamp 1667941163
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_236
timestamp 1667941163
transform 1 0 22816 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_248
timestamp 1667941163
transform 1 0 23920 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_260
timestamp 1667941163
transform 1 0 25024 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_272
timestamp 1667941163
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1667941163
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_367
timestamp 1667941163
transform 1 0 34868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_379
timestamp 1667941163
transform 1 0 35972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_38
timestamp 1667941163
transform 1 0 4600 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_50
timestamp 1667941163
transform 1 0 5704 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_62
timestamp 1667941163
transform 1 0 6808 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_74
timestamp 1667941163
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_100
timestamp 1667941163
transform 1 0 10304 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_106
timestamp 1667941163
transform 1 0 10856 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1667941163
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_117
timestamp 1667941163
transform 1 0 11868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_124
timestamp 1667941163
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1667941163
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_152
timestamp 1667941163
transform 1 0 15088 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_160
timestamp 1667941163
transform 1 0 15824 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_171
timestamp 1667941163
transform 1 0 16836 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_182
timestamp 1667941163
transform 1 0 17848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_202
timestamp 1667941163
transform 1 0 19688 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_210
timestamp 1667941163
transform 1 0 20424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_214
timestamp 1667941163
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_298
timestamp 1667941163
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1667941163
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1667941163
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1667941163
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_44
timestamp 1667941163
transform 1 0 5152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_50
timestamp 1667941163
transform 1 0 5704 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_133
timestamp 1667941163
transform 1 0 13340 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_138
timestamp 1667941163
transform 1 0 13800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_145
timestamp 1667941163
transform 1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_152
timestamp 1667941163
transform 1 0 15088 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1667941163
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_180
timestamp 1667941163
transform 1 0 17664 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_188
timestamp 1667941163
transform 1 0 18400 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_192
timestamp 1667941163
transform 1 0 18768 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_199
timestamp 1667941163
transform 1 0 19412 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_206
timestamp 1667941163
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1667941163
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_117
timestamp 1667941163
transform 1 0 11868 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_125
timestamp 1667941163
transform 1 0 12604 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_129
timestamp 1667941163
transform 1 0 12972 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1667941163
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1667941163
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_154
timestamp 1667941163
transform 1 0 15272 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_161
timestamp 1667941163
transform 1 0 15916 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1667941163
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_185
timestamp 1667941163
transform 1 0 18124 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_207
timestamp 1667941163
transform 1 0 20148 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_75
timestamp 1667941163
transform 1 0 8004 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_87
timestamp 1667941163
transform 1 0 9108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_99
timestamp 1667941163
transform 1 0 10212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_132
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_144
timestamp 1667941163
transform 1 0 14352 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_152
timestamp 1667941163
transform 1 0 15088 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_157
timestamp 1667941163
transform 1 0 15548 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_182
timestamp 1667941163
transform 1 0 17848 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_186
timestamp 1667941163
transform 1 0 18216 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_190
timestamp 1667941163
transform 1 0 18584 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_197
timestamp 1667941163
transform 1 0 19228 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_210
timestamp 1667941163
transform 1 0 20424 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_365
timestamp 1667941163
transform 1 0 34684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_369
timestamp 1667941163
transform 1 0 35052 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_381
timestamp 1667941163
transform 1 0 36156 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1667941163
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_401
timestamp 1667941163
transform 1 0 37996 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1667941163
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_179
timestamp 1667941163
transform 1 0 17572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_183
timestamp 1667941163
transform 1 0 17940 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_187
timestamp 1667941163
transform 1 0 18308 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_203
timestamp 1667941163
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_213
timestamp 1667941163
transform 1 0 20700 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_225
timestamp 1667941163
transform 1 0 21804 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_237
timestamp 1667941163
transform 1 0 22908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1667941163
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_21
timestamp 1667941163
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_33
timestamp 1667941163
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1667941163
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_173
timestamp 1667941163
transform 1 0 17020 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_177
timestamp 1667941163
transform 1 0 17388 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_189
timestamp 1667941163
transform 1 0 18492 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_203
timestamp 1667941163
transform 1 0 19780 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_210
timestamp 1667941163
transform 1 0 20424 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1667941163
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_365
timestamp 1667941163
transform 1 0 34684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_369
timestamp 1667941163
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_381
timestamp 1667941163
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1667941163
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1667941163
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_297
timestamp 1667941163
transform 1 0 28428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp 1667941163
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_31
timestamp 1667941163
transform 1 0 3956 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1667941163
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1667941163
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_8
timestamp 1667941163
transform 1 0 1840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1667941163
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_314
timestamp 1667941163
transform 1 0 29992 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_326
timestamp 1667941163
transform 1 0 31096 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_338
timestamp 1667941163
transform 1 0 32200 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_350
timestamp 1667941163
transform 1 0 33304 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1667941163
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_72
timestamp 1667941163
transform 1 0 7728 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1667941163
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1667941163
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1667941163
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1667941163
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1667941163
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_342
timestamp 1667941163
transform 1 0 32568 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_354
timestamp 1667941163
transform 1 0 33672 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_366
timestamp 1667941163
transform 1 0 34776 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_378
timestamp 1667941163
transform 1 0 35880 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_390
timestamp 1667941163
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_61
timestamp 1667941163
transform 1 0 6716 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_66
timestamp 1667941163
transform 1 0 7176 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_78
timestamp 1667941163
transform 1 0 8280 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_314
timestamp 1667941163
transform 1 0 29992 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_326
timestamp 1667941163
transform 1 0 31096 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_338
timestamp 1667941163
transform 1 0 32200 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_350
timestamp 1667941163
transform 1 0 33304 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1667941163
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_186
timestamp 1667941163
transform 1 0 18216 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_198
timestamp 1667941163
transform 1 0 19320 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_210
timestamp 1667941163
transform 1 0 20424 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1667941163
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_301
timestamp 1667941163
transform 1 0 28796 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_307
timestamp 1667941163
transform 1 0 29348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_319
timestamp 1667941163
transform 1 0 30452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1667941163
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_9
timestamp 1667941163
transform 1 0 1932 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1667941163
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_34
timestamp 1667941163
transform 1 0 4232 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_46
timestamp 1667941163
transform 1 0 5336 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_52
timestamp 1667941163
transform 1 0 5888 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_56
timestamp 1667941163
transform 1 0 6256 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_68
timestamp 1667941163
transform 1 0 7360 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1667941163
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_173
timestamp 1667941163
transform 1 0 17020 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_202
timestamp 1667941163
transform 1 0 19688 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_214
timestamp 1667941163
transform 1 0 20792 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_229
timestamp 1667941163
transform 1 0 22172 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_241
timestamp 1667941163
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1667941163
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_370
timestamp 1667941163
transform 1 0 35144 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_382
timestamp 1667941163
transform 1 0 36248 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_394
timestamp 1667941163
transform 1 0 37352 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1667941163
transform 1 0 38456 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_160
timestamp 1667941163
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_401
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_8
timestamp 1667941163
transform 1 0 1840 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1667941163
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_36
timestamp 1667941163
transform 1 0 4416 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_48
timestamp 1667941163
transform 1 0 5520 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_60
timestamp 1667941163
transform 1 0 6624 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_72
timestamp 1667941163
transform 1 0 7728 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_173
timestamp 1667941163
transform 1 0 17020 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_178
timestamp 1667941163
transform 1 0 17480 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_190
timestamp 1667941163
transform 1 0 18584 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_370
timestamp 1667941163
transform 1 0 35144 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_382
timestamp 1667941163
transform 1 0 36248 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_394
timestamp 1667941163
transform 1 0 37352 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1667941163
transform 1 0 38456 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_321
timestamp 1667941163
transform 1 0 30636 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_325
timestamp 1667941163
transform 1 0 31004 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_333
timestamp 1667941163
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1667941163
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_90
timestamp 1667941163
transform 1 0 9384 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_264
timestamp 1667941163
transform 1 0 25392 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_273
timestamp 1667941163
transform 1 0 26220 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_285
timestamp 1667941163
transform 1 0 27324 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_297
timestamp 1667941163
transform 1 0 28428 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp 1667941163
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_314
timestamp 1667941163
transform 1 0 29992 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_326
timestamp 1667941163
transform 1 0 31096 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_338
timestamp 1667941163
transform 1 0 32200 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_350
timestamp 1667941163
transform 1 0 33304 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 1667941163
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_62
timestamp 1667941163
transform 1 0 6808 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_74
timestamp 1667941163
transform 1 0 7912 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_86
timestamp 1667941163
transform 1 0 9016 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_98
timestamp 1667941163
transform 1 0 10120 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1667941163
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_243
timestamp 1667941163
transform 1 0 23460 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_255
timestamp 1667941163
transform 1 0 24564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_267
timestamp 1667941163
transform 1 0 25668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_368
timestamp 1667941163
transform 1 0 34960 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_380
timestamp 1667941163
transform 1 0 36064 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_8
timestamp 1667941163
transform 1 0 1840 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1667941163
transform 1 0 2944 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1667941163
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_68
timestamp 1667941163
transform 1 0 7360 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_80
timestamp 1667941163
transform 1 0 8464 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_227
timestamp 1667941163
transform 1 0 21988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_239
timestamp 1667941163
transform 1 0 23092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_272
timestamp 1667941163
transform 1 0 26128 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_284
timestamp 1667941163
transform 1 0 27232 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_296
timestamp 1667941163
transform 1 0 28336 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_314
timestamp 1667941163
transform 1 0 29992 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_326
timestamp 1667941163
transform 1 0 31096 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_338
timestamp 1667941163
transform 1 0 32200 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_350
timestamp 1667941163
transform 1 0 33304 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1667941163
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_370
timestamp 1667941163
transform 1 0 35144 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_382
timestamp 1667941163
transform 1 0 36248 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_394
timestamp 1667941163
transform 1 0 37352 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1667941163
transform 1 0 38456 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1667941163
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1667941163
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1667941163
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1667941163
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_73
timestamp 1667941163
transform 1 0 7820 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_77
timestamp 1667941163
transform 1 0 8188 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_89
timestamp 1667941163
transform 1 0 9292 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_101
timestamp 1667941163
transform 1 0 10396 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_109
timestamp 1667941163
transform 1 0 11132 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_117
timestamp 1667941163
transform 1 0 11868 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_121
timestamp 1667941163
transform 1 0 12236 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_133
timestamp 1667941163
transform 1 0 13340 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_145
timestamp 1667941163
transform 1 0 14444 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_157
timestamp 1667941163
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_165
timestamp 1667941163
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_190
timestamp 1667941163
transform 1 0 18584 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_202
timestamp 1667941163
transform 1 0 19688 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_207
timestamp 1667941163
transform 1 0 20148 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1667941163
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_286
timestamp 1667941163
transform 1 0 27416 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_298
timestamp 1667941163
transform 1 0 28520 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_310
timestamp 1667941163
transform 1 0 29624 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_322
timestamp 1667941163
transform 1 0 30728 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1667941163
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_352
timestamp 1667941163
transform 1 0 33488 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_364
timestamp 1667941163
transform 1 0 34592 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_376
timestamp 1667941163
transform 1 0 35696 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1667941163
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_49
timestamp 1667941163
transform 1 0 5612 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_117
timestamp 1667941163
transform 1 0 11868 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_122
timestamp 1667941163
transform 1 0 12328 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_134
timestamp 1667941163
transform 1 0 13432 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_149
timestamp 1667941163
transform 1 0 14812 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_155
timestamp 1667941163
transform 1 0 15364 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_170
timestamp 1667941163
transform 1 0 16744 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_176
timestamp 1667941163
transform 1 0 17296 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_180
timestamp 1667941163
transform 1 0 17664 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1667941163
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_220
timestamp 1667941163
transform 1 0 21344 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_232
timestamp 1667941163
transform 1 0 22448 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_243
timestamp 1667941163
transform 1 0 23460 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_317
timestamp 1667941163
transform 1 0 30268 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_322
timestamp 1667941163
transform 1 0 30728 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_334
timestamp 1667941163
transform 1 0 31832 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_346
timestamp 1667941163
transform 1 0 32936 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_358
timestamp 1667941163
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_11
timestamp 1667941163
transform 1 0 2116 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_17
timestamp 1667941163
transform 1 0 2668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_29
timestamp 1667941163
transform 1 0 3772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_41
timestamp 1667941163
transform 1 0 4876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1667941163
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_20
timestamp 1667941163
transform 1 0 2944 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_401
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_16
timestamp 1667941163
transform 1 0 2576 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_28
timestamp 1667941163
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_40
timestamp 1667941163
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1667941163
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_16
timestamp 1667941163
transform 1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_43
timestamp 1667941163
transform 1 0 5060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_49
timestamp 1667941163
transform 1 0 5612 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1667941163
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_65
timestamp 1667941163
transform 1 0 7084 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1667941163
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_104
timestamp 1667941163
transform 1 0 10672 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_118
timestamp 1667941163
transform 1 0 11960 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1667941163
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_149
timestamp 1667941163
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_203
timestamp 1667941163
transform 1 0 19780 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_211
timestamp 1667941163
transform 1 0 20516 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_216
timestamp 1667941163
transform 1 0 20976 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_233
timestamp 1667941163
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1667941163
transform 1 0 26220 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1667941163
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_286
timestamp 1667941163
transform 1 0 27416 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_298
timestamp 1667941163
transform 1 0 28520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1667941163
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_342
timestamp 1667941163
transform 1 0 32568 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_356
timestamp 1667941163
transform 1 0 33856 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_382
timestamp 1667941163
transform 1 0 36248 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_386
timestamp 1667941163
transform 1 0 36616 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0410_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17572 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0411_
timestamp 1667941163
transform 1 0 15180 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12420 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0413_
timestamp 1667941163
transform 1 0 14904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0414_
timestamp 1667941163
transform 1 0 16744 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1667941163
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0416_
timestamp 1667941163
transform 1 0 5704 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 4508 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_
timestamp 1667941163
transform 1 0 5060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 5336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 4968 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 22448 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 23276 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 23092 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 24196 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 23552 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform 1 0 21804 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 17296 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 21160 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 20516 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform 1 0 16100 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 16652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 12880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 10948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 10304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 10948 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 7728 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 18952 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform 1 0 18032 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 16652 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform 1 0 18676 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 22632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 24656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 18308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1667941163
transform 1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1667941163
transform 1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform 1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 22448 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform 1 0 14996 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 11592 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 11592 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform 1 0 11684 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 15088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 9476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 9016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 10304 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform 1 0 10948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform 1 0 8004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0480_
timestamp 1667941163
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1667941163
transform 1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 16100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0486_
timestamp 1667941163
transform 1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1667941163
transform 1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0488_
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1667941163
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1667941163
transform 1 0 7268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0493_
timestamp 1667941163
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1667941163
transform 1 0 16100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0495_
timestamp 1667941163
transform 1 0 15824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1667941163
transform 1 0 6624 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0499_
timestamp 1667941163
transform 1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0500_
timestamp 1667941163
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0501_
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 16100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1667941163
transform 1 0 16744 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0505_
timestamp 1667941163
transform 1 0 17480 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1667941163
transform 1 0 20148 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 20792 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 23184 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0510_
timestamp 1667941163
transform 1 0 23552 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0511_
timestamp 1667941163
transform 1 0 24196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0512_
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1667941163
transform 1 0 3220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 3128 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1667941163
transform 1 0 3772 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 20516 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0522_
timestamp 1667941163
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0523_
timestamp 1667941163
transform 1 0 19872 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0524_
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform 1 0 20608 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1667941163
transform 1 0 24380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 10580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1667941163
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0532_
timestamp 1667941163
transform 1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0533_
timestamp 1667941163
transform 1 0 14260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 18032 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1667941163
transform 1 0 15640 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 13432 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0540_
timestamp 1667941163
transform 1 0 14904 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0541_
timestamp 1667941163
transform 1 0 12052 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0542_
timestamp 1667941163
transform 1 0 14260 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 13248 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform 1 0 12880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1667941163
transform 1 0 15456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 16928 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 14076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0550_
timestamp 1667941163
transform 1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1667941163
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1667941163
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 15824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 9200 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0558_
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1667941163
transform 1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1667941163
transform 1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 10948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 10764 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0564_
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform 1 0 23184 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0568_
timestamp 1667941163
transform 1 0 20976 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0569_
timestamp 1667941163
transform 1 0 17572 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1667941163
transform 1 0 15640 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 21528 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 14168 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1667941163
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0577_
timestamp 1667941163
transform 1 0 15640 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1667941163
transform 1 0 15272 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 14996 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform 1 0 17572 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1667941163
transform 1 0 18492 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 13524 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 11960 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1667941163
transform 1 0 12972 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0586_
timestamp 1667941163
transform 1 0 12696 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0587_
timestamp 1667941163
transform 1 0 14352 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 14352 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0590_
timestamp 1667941163
transform 1 0 14720 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 15456 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1667941163
transform 1 0 15456 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0595_
timestamp 1667941163
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0596_
timestamp 1667941163
transform 1 0 20516 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1667941163
transform 1 0 19596 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 18216 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1667941163
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 23552 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1667941163
transform 1 0 23736 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0604_
timestamp 1667941163
transform 1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0605_
timestamp 1667941163
transform 1 0 24472 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1667941163
transform 1 0 25208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1667941163
transform 1 0 22264 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0609_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 11776 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 10948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0613_
timestamp 1667941163
transform 1 0 11592 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1667941163
transform 1 0 12880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1667941163
transform 1 0 14168 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 11776 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1667941163
transform 1 0 12420 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1667941163
transform 1 0 12420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 21160 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1667941163
transform 1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0622_
timestamp 1667941163
transform 1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0623_
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1667941163
transform 1 0 14720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1667941163
transform 1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1667941163
transform 1 0 23092 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 11592 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 10948 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1667941163
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 1667941163
transform 1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0632_
timestamp 1667941163
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1667941163
transform 1 0 14352 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1667941163
transform 1 0 18400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1667941163
transform 1 0 17664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1667941163
transform 1 0 6808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0640_
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0641_
timestamp 1667941163
transform 1 0 4324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1667941163
transform 1 0 6532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1667941163
transform 1 0 6992 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1667941163
transform 1 0 7820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 12144 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1667941163
transform 1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0649_
timestamp 1667941163
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 1667941163
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1667941163
transform 1 0 10764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1667941163
transform 1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1667941163
transform 1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 8464 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1667941163
transform 1 0 8372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0659_
timestamp 1667941163
transform 1 0 7176 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1667941163
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1667941163
transform 1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1667941163
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 16928 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 14904 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0667_
timestamp 1667941163
transform 1 0 12144 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0668_
timestamp 1667941163
transform 1 0 14996 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1667941163
transform 1 0 17572 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 20700 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1667941163
transform 1 0 20608 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1667941163
transform 1 0 19780 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 12880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 16836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0675_
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0676_
timestamp 1667941163
transform 1 0 17112 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0677_
timestamp 1667941163
transform 1 0 14444 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1667941163
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1667941163
transform 1 0 18768 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1667941163
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1667941163
transform 1 0 11224 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0685_
timestamp 1667941163
transform 1 0 14260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1667941163
transform 1 0 10304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1667941163
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0690_
timestamp 1667941163
transform 1 0 14628 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 23184 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 22632 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 21712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0694_
timestamp 1667941163
transform 1 0 21252 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0695_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0696_
timestamp 1667941163
transform 1 0 24196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1667941163
transform 1 0 23368 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 28336 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 25944 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 15364 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 6900 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 29716 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 33028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 18308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 9108 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 6532 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 6164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 5060 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 17940 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 3956 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 31832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 33120 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 33304 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 29716 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 7636 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 7360 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 29716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 34132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 29716 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 35420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 8004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 19412 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 7452 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 17112 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 11960 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0737_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 30728 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 2392 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 30452 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 20148 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 31464 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0748_
timestamp 1667941163
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 13432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 28244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 5612 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 28704 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 33856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 29716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 34592 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 22632 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 21712 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 37444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 8372 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 16744 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 9752 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 7636 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 7268 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 32292 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 28244 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 7728 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 29532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 31096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 21896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 19872 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 8096 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 12052 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 23184 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 15548 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 14720 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 17204 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 34132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 4324 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 29072 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0793_
timestamp 1667941163
transform 1 0 15088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0794_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0795_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2944 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 19412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0806_
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 2576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 18676 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 19320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 2392 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 23092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0817_
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0828_
timestamp 1667941163
transform 1 0 3956 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 18400 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 17756 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 18768 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 18400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0839_
timestamp 1667941163
transform 1 0 1840 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 2300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 3956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0850_
timestamp 1667941163
transform 1 0 1840 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 7544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 5152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 5336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 4508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 2944 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 3128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0861_
timestamp 1667941163
transform 1 0 1656 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1667941163
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1667941163
transform 1 0 4416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1667941163
transform 1 0 20700 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1667941163
transform 1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1667941163
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1667941163
transform 1 0 18768 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1667941163
transform 1 0 19412 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1667941163
transform 1 0 20056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1667941163
transform 1 0 17204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1667941163
transform 1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1667941163
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1667941163
transform 1 0 9936 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1667941163
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _0878_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0879_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0880_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6808 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0881_
timestamp 1667941163
transform 1 0 3956 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0882_
timestamp 1667941163
transform 1 0 4140 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0883_
timestamp 1667941163
transform 1 0 5060 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0884_
timestamp 1667941163
transform 1 0 2392 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0885_
timestamp 1667941163
transform 1 0 4508 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0886_
timestamp 1667941163
transform 1 0 11960 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0887_
timestamp 1667941163
transform 1 0 10580 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0888_
timestamp 1667941163
transform 1 0 13892 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0889_
timestamp 1667941163
transform 1 0 11684 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0890_
timestamp 1667941163
transform 1 0 11684 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0891_
timestamp 1667941163
transform 1 0 10304 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0892_
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0893_
timestamp 1667941163
transform 1 0 7912 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0894_
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0895_
timestamp 1667941163
transform 1 0 2024 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0896_
timestamp 1667941163
transform 1 0 11684 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0897_
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0898_
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0899_
timestamp 1667941163
transform 1 0 7728 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0901_
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0902_
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0903_
timestamp 1667941163
transform 1 0 9476 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0904_
timestamp 1667941163
transform 1 0 4140 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0905_
timestamp 1667941163
transform 1 0 7912 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 11684 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0907_
timestamp 1667941163
transform 1 0 6624 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0908_
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0909_
timestamp 1667941163
transform 1 0 8096 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0910_
timestamp 1667941163
transform 1 0 6808 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0911_
timestamp 1667941163
transform 1 0 10488 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 14260 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0913_
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 9200 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0915_
timestamp 1667941163
transform 1 0 9108 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0916_
timestamp 1667941163
transform 1 0 1932 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0917_
timestamp 1667941163
transform 1 0 3956 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1667941163
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1667941163
transform 1 0 1656 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0921_
timestamp 1667941163
transform 1 0 2300 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 6716 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0923_
timestamp 1667941163
transform 1 0 3864 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 9384 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 10120 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 1656 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0927_
timestamp 1667941163
transform 1 0 11684 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 8280 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0929_
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 5888 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 6808 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 1564 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0934_
timestamp 1667941163
transform 1 0 4968 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0936_
timestamp 1667941163
transform 1 0 4048 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 5428 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0938_
timestamp 1667941163
transform 1 0 2852 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 1656 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0940_
timestamp 1667941163
transform 1 0 6624 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0941_
timestamp 1667941163
transform 1 0 4140 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0942_
timestamp 1667941163
transform 1 0 6992 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1667941163
transform 1 0 1656 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1667941163
transform 1 0 10120 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0946_
timestamp 1667941163
transform 1 0 5520 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0947_
timestamp 1667941163
transform 1 0 3956 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0948_
timestamp 1667941163
transform 1 0 14260 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0949_
timestamp 1667941163
transform 1 0 13984 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0950_
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform 1 0 1656 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0952_
timestamp 1667941163
transform 1 0 9292 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 13984 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1667941163
transform 1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 34868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 4048 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1667941163
transform 1 0 27140 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1667941163
transform 1 0 16468 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 15088 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 5244 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1667941163
transform 1 0 23184 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1667941163
transform 1 0 34960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1667941163
transform 1 0 32292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 34776 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 1748 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 21068 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 36248 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 34684 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 34776 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 27140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 4968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 34224 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 7912 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 38088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 4140 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform 1 0 5704 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 18308 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 4416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 1748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 5428 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 35052 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1030_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1031_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1031__100 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23276 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1032_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1033_
timestamp 1667941163
transform 1 0 22356 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1034_
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1035_
timestamp 1667941163
transform 1 0 23092 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1036_
timestamp 1667941163
transform 1 0 17572 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1037__101
timestamp 1667941163
transform 1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1037_
timestamp 1667941163
transform 1 0 13064 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1038_
timestamp 1667941163
transform 1 0 13984 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1039_
timestamp 1667941163
transform 1 0 15640 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1040_
timestamp 1667941163
transform 1 0 10488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1041_
timestamp 1667941163
transform 1 0 18216 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1042_
timestamp 1667941163
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1043__102
timestamp 1667941163
transform 1 0 20608 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1043_
timestamp 1667941163
transform 1 0 18400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1044_
timestamp 1667941163
transform 1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1045_
timestamp 1667941163
transform 1 0 14628 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1046_
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1047_
timestamp 1667941163
transform 1 0 17480 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1048_
timestamp 1667941163
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1049__103
timestamp 1667941163
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1049_
timestamp 1667941163
transform 1 0 19504 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1050_
timestamp 1667941163
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1051_
timestamp 1667941163
transform 1 0 17020 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1052_
timestamp 1667941163
transform 1 0 20056 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1053_
timestamp 1667941163
transform 1 0 15088 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1054_
timestamp 1667941163
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1055__104
timestamp 1667941163
transform 1 0 8096 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1055_
timestamp 1667941163
transform 1 0 9844 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1056_
timestamp 1667941163
transform 1 0 9200 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1057_
timestamp 1667941163
transform 1 0 7820 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1058_
timestamp 1667941163
transform 1 0 10120 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1059_
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1060_
timestamp 1667941163
transform 1 0 12420 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1061_
timestamp 1667941163
transform 1 0 11408 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1061__105
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1062_
timestamp 1667941163
transform 1 0 12052 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1063_
timestamp 1667941163
transform 1 0 12512 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1064_
timestamp 1667941163
transform 1 0 9476 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1065_
timestamp 1667941163
transform 1 0 11868 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1066_
timestamp 1667941163
transform 1 0 6532 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1067_
timestamp 1667941163
transform 1 0 7360 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1067__106
timestamp 1667941163
transform 1 0 6716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1068_
timestamp 1667941163
transform 1 0 8648 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1069_
timestamp 1667941163
transform 1 0 7636 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1070_
timestamp 1667941163
transform 1 0 6256 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1071_
timestamp 1667941163
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1072_
timestamp 1667941163
transform 1 0 16192 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1073_
timestamp 1667941163
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1073__107
timestamp 1667941163
transform 1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1074_
timestamp 1667941163
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1075_
timestamp 1667941163
transform 1 0 13892 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 18216 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1077_
timestamp 1667941163
transform 1 0 12144 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1078_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1079__108
timestamp 1667941163
transform 1 0 22172 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1079_
timestamp 1667941163
transform 1 0 21068 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1080_
timestamp 1667941163
transform 1 0 21712 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1081_
timestamp 1667941163
transform 1 0 18492 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1082_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1083_
timestamp 1667941163
transform 1 0 20608 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1084_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1085_
timestamp 1667941163
transform 1 0 16468 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1085__109
timestamp 1667941163
transform 1 0 13524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1086_
timestamp 1667941163
transform 1 0 14168 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1087_
timestamp 1667941163
transform 1 0 15456 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1088_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1089_
timestamp 1667941163
transform 1 0 12052 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1090_
timestamp 1667941163
transform 1 0 23276 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1091__110
timestamp 1667941163
transform 1 0 24196 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1091_
timestamp 1667941163
transform 1 0 22448 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1092_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1093_
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1094_
timestamp 1667941163
transform 1 0 21528 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1095_
timestamp 1667941163
transform 1 0 22080 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform 1 0 19504 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1097_
timestamp 1667941163
transform 1 0 19320 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1097__111
timestamp 1667941163
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1098_
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1099_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1100_
timestamp 1667941163
transform 1 0 18768 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1101_
timestamp 1667941163
transform 1 0 15548 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1102_
timestamp 1667941163
transform 1 0 16008 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1103__112
timestamp 1667941163
transform 1 0 14260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1103_
timestamp 1667941163
transform 1 0 15732 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1104_
timestamp 1667941163
transform 1 0 12880 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1105_
timestamp 1667941163
transform 1 0 14260 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1106_
timestamp 1667941163
transform 1 0 15732 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1107_
timestamp 1667941163
transform 1 0 11868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1108_
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1109__113
timestamp 1667941163
transform 1 0 19136 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1109_
timestamp 1667941163
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1110_
timestamp 1667941163
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1111_
timestamp 1667941163
transform 1 0 15456 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1112_
timestamp 1667941163
transform 1 0 19504 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1113_
timestamp 1667941163
transform 1 0 13156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1114_
timestamp 1667941163
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1115__114
timestamp 1667941163
transform 1 0 19412 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1116_
timestamp 1667941163
transform 1 0 20608 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1117_
timestamp 1667941163
transform 1 0 15548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1118_
timestamp 1667941163
transform 1 0 20424 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1119_
timestamp 1667941163
transform 1 0 21712 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1120_
timestamp 1667941163
transform 1 0 13156 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1121__115
timestamp 1667941163
transform 1 0 12880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1121_
timestamp 1667941163
transform 1 0 14260 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1122_
timestamp 1667941163
transform 1 0 20516 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1123_
timestamp 1667941163
transform 1 0 12604 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1124_
timestamp 1667941163
transform 1 0 13064 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1125_
timestamp 1667941163
transform 1 0 20976 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1126_
timestamp 1667941163
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1127_
timestamp 1667941163
transform 1 0 16836 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1127__116
timestamp 1667941163
transform 1 0 14444 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1128_
timestamp 1667941163
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1129_
timestamp 1667941163
transform 1 0 14260 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1130_
timestamp 1667941163
transform 1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1131_
timestamp 1667941163
transform 1 0 15824 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 17112 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1133_
timestamp 1667941163
transform 1 0 16468 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1133__117
timestamp 1667941163
transform 1 0 15548 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1134_
timestamp 1667941163
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1136_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1137_
timestamp 1667941163
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1139_
timestamp 1667941163
transform 1 0 16468 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1139__118
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1140_
timestamp 1667941163
transform 1 0 14352 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform 1 0 15548 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1142_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1143_
timestamp 1667941163
transform 1 0 12696 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 19872 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1145_
timestamp 1667941163
transform 1 0 18216 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1145__119
timestamp 1667941163
transform 1 0 15456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1146_
timestamp 1667941163
transform 1 0 18400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 19780 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1148_
timestamp 1667941163
transform 1 0 18124 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1149_
timestamp 1667941163
transform 1 0 18768 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1150__120
timestamp 1667941163
transform 1 0 3772 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1150_
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1151_
timestamp 1667941163
transform 1 0 3864 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1152_
timestamp 1667941163
transform 1 0 6532 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1153_
timestamp 1667941163
transform 1 0 4600 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1154__121
timestamp 1667941163
transform 1 0 25300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1154_
timestamp 1667941163
transform 1 0 23460 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1155_
timestamp 1667941163
transform 1 0 23092 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 23000 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1157_
timestamp 1667941163
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1158__122
timestamp 1667941163
transform 1 0 21252 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1158_
timestamp 1667941163
transform 1 0 20148 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1159_
timestamp 1667941163
transform 1 0 19504 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1160_
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1161_
timestamp 1667941163
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1162__123
timestamp 1667941163
transform 1 0 7176 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 6992 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1163_
timestamp 1667941163
transform 1 0 9200 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1164_
timestamp 1667941163
transform 1 0 8280 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1165_
timestamp 1667941163
transform 1 0 10488 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 16836 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1166__124
timestamp 1667941163
transform 1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1167_
timestamp 1667941163
transform 1 0 13064 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 14260 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1169_
timestamp 1667941163
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1170_
timestamp 1667941163
transform 1 0 10120 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1170__125
timestamp 1667941163
transform 1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1171_
timestamp 1667941163
transform 1 0 14260 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1172_
timestamp 1667941163
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1173_
timestamp 1667941163
transform 1 0 11408 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1174__126
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1174_
timestamp 1667941163
transform 1 0 17204 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 14260 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1176_
timestamp 1667941163
transform 1 0 12972 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1177_
timestamp 1667941163
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1178_
timestamp 1667941163
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1178__127
timestamp 1667941163
transform 1 0 8096 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1179_
timestamp 1667941163
transform 1 0 13432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1180_
timestamp 1667941163
transform 1 0 9200 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1181_
timestamp 1667941163
transform 1 0 11960 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1182__128
timestamp 1667941163
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 10396 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 13156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 13984 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform 1 0 12328 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1186__129
timestamp 1667941163
transform 1 0 18124 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1187_
timestamp 1667941163
transform 1 0 12328 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1188_
timestamp 1667941163
transform 1 0 17020 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1189_
timestamp 1667941163
transform 1 0 15364 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1190__130
timestamp 1667941163
transform 1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1190_
timestamp 1667941163
transform 1 0 23184 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 20516 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1192_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform 1 0 20792 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1194__131
timestamp 1667941163
transform 1 0 20148 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1194_
timestamp 1667941163
transform 1 0 19872 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1195_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 19596 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1197_
timestamp 1667941163
transform 1 0 19044 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1198__132
timestamp 1667941163
transform 1 0 8740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1198_
timestamp 1667941163
transform 1 0 8740 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1199_
timestamp 1667941163
transform 1 0 11224 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1200_
timestamp 1667941163
transform 1 0 9568 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 11684 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1202__133
timestamp 1667941163
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 15272 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform 1 0 16008 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1204_
timestamp 1667941163
transform 1 0 15364 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1205_
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1206__134
timestamp 1667941163
transform 1 0 17112 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1206_
timestamp 1667941163
transform 1 0 17020 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1207_
timestamp 1667941163
transform 1 0 20424 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1208_
timestamp 1667941163
transform 1 0 17296 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 20700 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1210__135
timestamp 1667941163
transform 1 0 22540 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1210_
timestamp 1667941163
transform 1 0 22448 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1211_
timestamp 1667941163
transform 1 0 22172 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1212_
timestamp 1667941163
transform 1 0 22632 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 22448 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 4508 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1214__136
timestamp 1667941163
transform 1 0 4692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 4324 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1216_
timestamp 1667941163
transform 1 0 5152 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1217_
timestamp 1667941163
transform 1 0 3956 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1218_
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1218__137
timestamp 1667941163
transform 1 0 21160 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1219_
timestamp 1667941163
transform 1 0 16192 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1220_
timestamp 1667941163
transform 1 0 19412 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1221_
timestamp 1667941163
transform 1 0 13892 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 1564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 38088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 38088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 23920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 38088 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 22448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 38088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 1564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 36708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 38088 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 20700 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 12972 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 38088 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 38088 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1667941163
transform 1 0 2576 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 36708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 36708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 1564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 38088 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 30452 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 2300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 38088 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 14904 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 9108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 5244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 37996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 1564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 37996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 18584 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 19872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
<< labels >>
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 ccff_head
port 0 nsew signal input
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 2 nsew signal input
flabel metal3 s 39200 11568 39800 11688 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 3 nsew signal input
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 4 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 5 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_right_in[13]
port 6 nsew signal input
flabel metal2 s 15474 200 15530 800 0 FreeSans 224 90 0 0 chanx_right_in[14]
port 7 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chanx_right_in[15]
port 8 nsew signal input
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 9 nsew signal input
flabel metal3 s 39200 31288 39800 31408 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 10 nsew signal input
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_right_in[18]
port 11 nsew signal input
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_right_in[1]
port 12 nsew signal input
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 13 nsew signal input
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 14 nsew signal input
flabel metal3 s 39200 19728 39800 19848 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 15 nsew signal input
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chanx_right_in[5]
port 16 nsew signal input
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 17 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 18 nsew signal input
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 19 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 20 nsew signal input
flabel metal3 s 39200 34688 39800 34808 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 21 nsew signal tristate
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 22 nsew signal tristate
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 23 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 24 nsew signal tristate
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_right_out[13]
port 25 nsew signal tristate
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 26 nsew signal tristate
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 27 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 28 nsew signal tristate
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 29 nsew signal tristate
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 30 nsew signal tristate
flabel metal3 s 39200 36728 39800 36848 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 31 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 32 nsew signal tristate
flabel metal2 s 23846 39200 23902 39800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 33 nsew signal tristate
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 34 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 35 nsew signal tristate
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 36 nsew signal tristate
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 37 nsew signal tristate
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 38 nsew signal tristate
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 39 nsew signal tristate
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal2 s 20626 39200 20682 39800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal3 s 200 2728 800 2848 0 FreeSans 480 0 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal2 s 34794 39200 34850 39800 0 FreeSans 224 90 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal2 s 2594 200 2650 800 0 FreeSans 224 90 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal3 s 200 16328 800 16448 0 FreeSans 480 0 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal3 s 200 8168 800 8288 0 FreeSans 480 0 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal3 s 200 12928 800 13048 0 FreeSans 480 0 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 pReset
port 78 nsew signal input
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 prog_clk
port 79 nsew signal input
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 80 nsew signal input
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 81 nsew signal input
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 82 nsew signal input
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 83 nsew signal input
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 84 nsew signal input
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 85 nsew signal input
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 86 nsew signal input
flabel metal2 s 7746 200 7802 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 87 nsew signal input
flabel metal2 s 12254 200 12310 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 88 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 89 nsew signal input
flabel metal3 s 39200 23128 39800 23248 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 90 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 91 nsew signal input
flabel metal2 s 31574 39200 31630 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 92 nsew signal input
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 93 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 94 nsew signal input
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 95 nsew signal input
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 96 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 97 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 98 nsew signal input
flabel metal3 s 39200 18368 39800 18488 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 99 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 16928 2006 16928 2006 0 _0000_
rlabel metal1 6263 2346 6263 2346 0 _0001_
rlabel metal2 10258 2941 10258 2941 0 _0002_
rlabel metal1 17526 4182 17526 4182 0 _0003_
rlabel metal1 19550 3910 19550 3910 0 _0004_
rlabel metal1 13853 2346 13853 2346 0 _0005_
rlabel via2 17526 4811 17526 4811 0 _0006_
rlabel metal1 18446 3570 18446 3570 0 _0007_
rlabel metal1 12013 5678 12013 5678 0 _0008_
rlabel metal1 16843 5610 16843 5610 0 _0009_
rlabel metal1 18124 5338 18124 5338 0 _0010_
rlabel metal1 19964 4794 19964 4794 0 _0011_
rlabel metal1 18216 4046 18216 4046 0 _0012_
rlabel via2 18538 8517 18538 8517 0 _0013_
rlabel metal2 19182 2482 19182 2482 0 _0014_
rlabel metal2 2898 15198 2898 15198 0 _0015_
rlabel metal1 2070 16966 2070 16966 0 _0016_
rlabel metal1 3273 12886 3273 12886 0 _0017_
rlabel metal1 21022 5338 21022 5338 0 _0018_
rlabel metal1 21022 3910 21022 3910 0 _0019_
rlabel metal3 5359 12580 5359 12580 0 _0020_
rlabel metal1 9154 5746 9154 5746 0 _0021_
rlabel metal1 19780 6766 19780 6766 0 _0022_
rlabel metal2 7314 6494 7314 6494 0 _0023_
rlabel metal3 2599 15436 2599 15436 0 _0024_
rlabel metal1 6762 6086 6762 6086 0 _0025_
rlabel metal1 7130 5882 7130 5882 0 _0026_
rlabel metal1 6808 7514 6808 7514 0 _0027_
rlabel metal1 5474 6290 5474 6290 0 _0028_
rlabel metal1 6256 5338 6256 5338 0 _0029_
rlabel metal1 4416 5338 4416 5338 0 _0030_
rlabel metal1 5658 13192 5658 13192 0 _0031_
rlabel metal1 7038 6154 7038 6154 0 _0032_
rlabel metal3 3818 11628 3818 11628 0 _0033_
rlabel metal1 3404 15878 3404 15878 0 _0034_
rlabel metal1 21390 5882 21390 5882 0 _0035_
rlabel metal1 21528 4794 21528 4794 0 _0036_
rlabel metal1 20332 4658 20332 4658 0 _0037_
rlabel metal2 5612 14212 5612 14212 0 _0038_
rlabel metal1 20884 5882 20884 5882 0 _0039_
rlabel metal1 20976 4794 20976 4794 0 _0040_
rlabel metal2 13662 12920 13662 12920 0 _0041_
rlabel metal2 18906 7888 18906 7888 0 _0042_
rlabel metal3 14996 6664 14996 6664 0 _0043_
rlabel metal1 20424 4998 20424 4998 0 _0044_
rlabel metal1 16567 3434 16567 3434 0 _0045_
rlabel metal2 17986 3230 17986 3230 0 _0046_
rlabel metal2 18906 2040 18906 2040 0 _0047_
rlabel metal1 3733 2346 3733 2346 0 _0048_
rlabel metal2 10074 3400 10074 3400 0 _0049_
rlabel metal1 10810 4488 10810 4488 0 _0050_
rlabel via2 21390 6171 21390 6171 0 _0051_
rlabel via2 20102 6341 20102 6341 0 _0052_
rlabel metal1 14996 1122 14996 1122 0 _0053_
rlabel via2 19550 5253 19550 5253 0 _0054_
rlabel metal3 13754 1292 13754 1292 0 _0055_
rlabel metal2 20286 1751 20286 1751 0 _0056_
rlabel metal2 20102 1853 20102 1853 0 _0057_
rlabel metal1 6263 4522 6263 4522 0 _0058_
rlabel metal3 17204 2652 17204 2652 0 _0059_
rlabel metal1 12427 4522 12427 4522 0 _0060_
rlabel via3 15341 6868 15341 6868 0 _0061_
rlabel metal1 13570 4216 13570 4216 0 _0062_
rlabel via3 2691 16796 2691 16796 0 _0063_
rlabel metal2 11178 6307 11178 6307 0 _0064_
rlabel metal1 18768 6426 18768 6426 0 _0065_
rlabel metal1 19366 6426 19366 6426 0 _0066_
rlabel metal1 13110 1530 13110 1530 0 _0067_
rlabel metal1 2530 6392 2530 6392 0 _0068_
rlabel metal2 18354 3791 18354 3791 0 _0069_
rlabel via2 22770 2499 22770 2499 0 _0070_
rlabel metal2 19366 2210 19366 2210 0 _0071_
rlabel metal2 19550 3927 19550 3927 0 _0072_
rlabel metal1 15785 2414 15785 2414 0 _0073_
rlabel metal2 13294 1802 13294 1802 0 _0074_
rlabel via2 21482 3723 21482 3723 0 _0075_
rlabel metal1 13570 9146 13570 9146 0 _0076_
rlabel metal2 16790 16966 16790 16966 0 _0077_
rlabel metal1 5244 15130 5244 15130 0 _0078_
rlabel metal1 5290 16218 5290 16218 0 _0079_
rlabel metal1 23782 17306 23782 17306 0 _0080_
rlabel metal1 23000 20570 23000 20570 0 _0081_
rlabel metal1 20976 21862 20976 21862 0 _0082_
rlabel metal2 16146 24004 16146 24004 0 _0083_
rlabel metal1 16238 7344 16238 7344 0 _0084_
rlabel metal1 12696 16762 12696 16762 0 _0085_
rlabel metal1 10764 21658 10764 21658 0 _0086_
rlabel metal1 8602 20944 8602 20944 0 _0087_
rlabel metal1 18906 23018 18906 23018 0 _0088_
rlabel metal1 23460 11322 23460 11322 0 _0089_
rlabel metal2 18354 24004 18354 24004 0 _0090_
rlabel metal2 20654 8058 20654 8058 0 _0091_
rlabel metal2 22678 7242 22678 7242 0 _0092_
rlabel metal2 11638 21148 11638 21148 0 _0093_
rlabel metal1 16928 19346 16928 19346 0 _0094_
rlabel metal1 9522 11118 9522 11118 0 _0095_
rlabel metal1 16790 3604 16790 3604 0 _0096_
rlabel metal1 11040 16558 11040 16558 0 _0097_
rlabel metal2 8234 13498 8234 13498 0 _0098_
rlabel metal1 11316 6154 11316 6154 0 _0099_
rlabel metal1 16284 6426 16284 6426 0 _0100_
rlabel metal2 9430 9588 9430 9588 0 _0101_
rlabel metal1 9752 16218 9752 16218 0 _0102_
rlabel metal2 17710 6783 17710 6783 0 _0103_
rlabel metal2 16146 4998 16146 4998 0 _0104_
rlabel metal1 6624 14246 6624 14246 0 _0105_
rlabel metal1 7314 17612 7314 17612 0 _0106_
rlabel metal1 16974 18938 16974 18938 0 _0107_
rlabel metal1 20608 10234 20608 10234 0 _0108_
rlabel metal1 24012 13498 24012 13498 0 _0109_
rlabel metal1 24426 10778 24426 10778 0 _0110_
rlabel metal2 3450 14586 3450 14586 0 _0111_
rlabel metal1 4002 15028 4002 15028 0 _0112_
rlabel metal1 20102 12852 20102 12852 0 _0113_
rlabel metal1 20838 19856 20838 19856 0 _0114_
rlabel metal2 24610 16286 24610 16286 0 _0115_
rlabel metal1 12006 12852 12006 12852 0 _0116_
rlabel metal2 14306 8602 14306 8602 0 _0117_
rlabel viali 15870 10031 15870 10031 0 _0118_
rlabel metal1 14950 11832 14950 11832 0 _0119_
rlabel viali 16330 13905 16330 13905 0 _0120_
rlabel metal1 15272 13906 15272 13906 0 _0121_
rlabel metal1 13018 9520 13018 9520 0 _0122_
rlabel metal2 9890 6596 9890 6596 0 _0123_
rlabel metal1 15502 11322 15502 11322 0 _0124_
rlabel metal1 21344 17646 21344 17646 0 _0125_
rlabel metal1 11178 19890 11178 19890 0 _0126_
rlabel metal1 11270 18598 11270 18598 0 _0127_
rlabel metal1 23184 16218 23184 16218 0 _0128_
rlabel metal1 17572 6970 17572 6970 0 _0129_
rlabel metal1 21436 11866 21436 11866 0 _0130_
rlabel metal1 15410 21658 15410 21658 0 _0131_
rlabel metal2 15226 23290 15226 23290 0 _0132_
rlabel metal1 18170 21862 18170 21862 0 _0133_
rlabel metal2 12926 23290 12926 23290 0 _0134_
rlabel metal1 14720 22610 14720 22610 0 _0135_
rlabel metal1 14352 19482 14352 19482 0 _0136_
rlabel metal1 18400 17646 18400 17646 0 _0137_
rlabel metal1 20286 12614 20286 12614 0 _0138_
rlabel metal1 18262 16524 18262 16524 0 _0139_
rlabel metal1 23644 16966 23644 16966 0 _0140_
rlabel metal1 24978 19482 24978 19482 0 _0141_
rlabel metal1 23552 18938 23552 18938 0 _0142_
rlabel metal2 11822 16490 11822 16490 0 _0143_
rlabel metal1 12926 17272 12926 17272 0 _0144_
rlabel metal2 12374 17884 12374 17884 0 _0145_
rlabel metal1 23276 15674 23276 15674 0 _0146_
rlabel metal1 14950 16524 14950 16524 0 _0147_
rlabel metal1 23414 14994 23414 14994 0 _0148_
rlabel metal1 10534 14348 10534 14348 0 _0149_
rlabel metal1 14582 13260 14582 13260 0 _0150_
rlabel metal2 18446 11764 18446 11764 0 _0151_
rlabel metal1 6440 14042 6440 14042 0 _0152_
rlabel metal1 5106 13498 5106 13498 0 _0153_
rlabel metal2 8050 15436 8050 15436 0 _0154_
rlabel metal2 10534 12988 10534 12988 0 _0155_
rlabel metal1 10672 12206 10672 12206 0 _0156_
rlabel metal1 9384 17850 9384 17850 0 _0157_
rlabel metal2 8602 17782 8602 17782 0 _0158_
rlabel metal1 7314 15130 7314 15130 0 _0159_
rlabel metal1 8602 19788 8602 19788 0 _0160_
rlabel metal1 12328 14586 12328 14586 0 _0161_
rlabel metal1 16422 13158 16422 13158 0 _0162_
rlabel metal1 20332 13498 20332 13498 0 _0163_
rlabel metal1 17388 18938 17388 18938 0 _0164_
rlabel metal2 14490 20468 14490 20468 0 _0165_
rlabel metal1 18860 20570 18860 20570 0 _0166_
rlabel metal2 14490 12580 14490 12580 0 _0167_
rlabel metal1 10994 18258 10994 18258 0 _0168_
rlabel metal2 14858 17850 14858 17850 0 _0169_
rlabel viali 22218 12817 22218 12817 0 _0170_
rlabel metal1 23920 12614 23920 12614 0 _0171_
rlabel metal1 17066 3502 17066 3502 0 _0172_
rlabel metal3 15732 3808 15732 3808 0 _0173_
rlabel metal1 22908 2414 22908 2414 0 _0174_
rlabel metal1 17802 4080 17802 4080 0 _0175_
rlabel metal1 17204 4590 17204 4590 0 _0176_
rlabel metal1 2162 17170 2162 17170 0 _0177_
rlabel metal1 3174 16116 3174 16116 0 _0178_
rlabel metal1 18814 7344 18814 7344 0 _0179_
rlabel metal2 24702 12002 24702 12002 0 _0180_
rlabel metal1 23644 10778 23644 10778 0 _0181_
rlabel metal2 22218 13396 22218 13396 0 _0182_
rlabel metal1 22678 11866 22678 11866 0 _0183_
rlabel metal1 21758 13498 21758 13498 0 _0184_
rlabel metal2 23322 9860 23322 9860 0 _0185_
rlabel metal1 17480 17646 17480 17646 0 _0186_
rlabel via2 12558 18139 12558 18139 0 _0187_
rlabel metal2 14168 13838 14168 13838 0 _0188_
rlabel metal1 15410 11186 15410 11186 0 _0189_
rlabel metal1 10718 19346 10718 19346 0 _0190_
rlabel metal1 18308 12954 18308 12954 0 _0191_
rlabel metal1 15502 20434 15502 20434 0 _0192_
rlabel metal2 18722 21284 18722 21284 0 _0193_
rlabel metal1 17388 20434 17388 20434 0 _0194_
rlabel metal1 13938 20978 13938 20978 0 _0195_
rlabel metal1 19642 21012 19642 21012 0 _0196_
rlabel metal1 17342 20978 17342 20978 0 _0197_
rlabel metal1 18216 14450 18216 14450 0 _0198_
rlabel metal1 19918 14042 19918 14042 0 _0199_
rlabel metal2 12650 15708 12650 15708 0 _0200_
rlabel metal1 17158 11866 17158 11866 0 _0201_
rlabel metal2 20838 15300 20838 15300 0 _0202_
rlabel metal2 15042 15062 15042 15062 0 _0203_
rlabel metal2 7222 16048 7222 16048 0 _0204_
rlabel metal1 9246 19890 9246 19890 0 _0205_
rlabel metal1 9200 17170 9200 17170 0 _0206_
rlabel metal1 8510 15130 8510 15130 0 _0207_
rlabel metal2 10350 21148 10350 21148 0 _0208_
rlabel metal1 8832 16626 8832 16626 0 _0209_
rlabel metal1 12604 12886 12604 12886 0 _0210_
rlabel metal2 9062 18530 9062 18530 0 _0211_
rlabel metal1 10534 12614 10534 12614 0 _0212_
rlabel metal1 12558 12104 12558 12104 0 _0213_
rlabel metal1 9108 18802 9108 18802 0 _0214_
rlabel metal1 11592 13362 11592 13362 0 _0215_
rlabel metal1 6670 14790 6670 14790 0 _0216_
rlabel metal1 7728 15130 7728 15130 0 _0217_
rlabel metal1 8602 12818 8602 12818 0 _0218_
rlabel metal1 6992 13838 6992 13838 0 _0219_
rlabel metal2 6486 16796 6486 16796 0 _0220_
rlabel metal1 9384 7786 9384 7786 0 _0221_
rlabel metal1 14490 13498 14490 13498 0 _0222_
rlabel metal1 18400 13294 18400 13294 0 _0223_
rlabel metal1 10534 14586 10534 14586 0 _0224_
rlabel metal2 11730 14824 11730 14824 0 _0225_
rlabel metal2 18630 10404 18630 10404 0 _0226_
rlabel metal2 11086 14722 11086 14722 0 _0227_
rlabel metal1 17204 15402 17204 15402 0 _0228_
rlabel metal1 23046 15130 23046 15130 0 _0229_
rlabel metal1 21942 16626 21942 16626 0 _0230_
rlabel metal1 16836 16150 16836 16150 0 _0231_
rlabel metal2 22678 14756 22678 14756 0 _0232_
rlabel metal2 21298 15878 21298 15878 0 _0233_
rlabel metal1 17066 18360 17066 18360 0 _0234_
rlabel metal1 16698 17578 16698 17578 0 _0235_
rlabel metal1 14398 17068 14398 17068 0 _0236_
rlabel metal1 14858 18326 14858 18326 0 _0237_
rlabel metal1 17066 17068 17066 17068 0 _0238_
rlabel metal2 11086 18292 11086 18292 0 _0239_
rlabel metal1 24380 19414 24380 19414 0 _0240_
rlabel metal2 24610 20196 24610 20196 0 _0241_
rlabel metal2 22862 16932 22862 16932 0 _0242_
rlabel metal1 23414 18394 23414 18394 0 _0243_
rlabel metal1 23023 19958 23023 19958 0 _0244_
rlabel metal1 23138 16014 23138 16014 0 _0245_
rlabel metal1 19596 14246 19596 14246 0 _0246_
rlabel metal1 18768 16422 18768 16422 0 _0247_
rlabel metal1 18906 17850 18906 17850 0 _0248_
rlabel metal2 20102 12546 20102 12546 0 _0249_
rlabel metal1 18676 18394 18676 18394 0 _0250_
rlabel metal1 15686 10778 15686 10778 0 _0251_
rlabel metal1 15548 22406 15548 22406 0 _0252_
rlabel metal1 14858 19890 14858 19890 0 _0253_
rlabel metal1 12926 22066 12926 22066 0 _0254_
rlabel metal1 14076 22406 14076 22406 0 _0255_
rlabel metal1 15226 20570 15226 20570 0 _0256_
rlabel metal2 12098 22780 12098 22780 0 _0257_
rlabel metal1 17066 22712 17066 22712 0 _0258_
rlabel metal1 18492 22066 18492 22066 0 _0259_
rlabel metal1 15732 21522 15732 21522 0 _0260_
rlabel metal1 14996 22678 14996 22678 0 _0261_
rlabel metal1 19596 21522 19596 21522 0 _0262_
rlabel metal1 13432 21522 13432 21522 0 _0263_
rlabel metal1 16422 8058 16422 8058 0 _0264_
rlabel metal2 21206 11934 21206 11934 0 _0265_
rlabel metal1 20930 17306 20930 17306 0 _0266_
rlabel metal2 18262 8058 18262 8058 0 _0267_
rlabel metal1 20654 12172 20654 12172 0 _0268_
rlabel metal1 21574 8874 21574 8874 0 _0269_
rlabel metal1 13202 19414 13202 19414 0 _0270_
rlabel metal2 13478 19278 13478 19278 0 _0271_
rlabel metal1 20838 17850 20838 17850 0 _0272_
rlabel metal1 12650 18632 12650 18632 0 _0273_
rlabel metal1 12696 16218 12696 16218 0 _0274_
rlabel metal2 21206 18972 21206 18972 0 _0275_
rlabel metal2 13202 7344 13202 7344 0 _0276_
rlabel metal2 17066 12818 17066 12818 0 _0277_
rlabel metal2 13294 9180 13294 9180 0 _0278_
rlabel metal2 9338 6800 9338 6800 0 _0279_
rlabel metal1 16192 10778 16192 10778 0 _0280_
rlabel metal1 16560 6834 16560 6834 0 _0281_
rlabel metal1 16284 13770 16284 13770 0 _0282_
rlabel metal1 15502 13804 15502 13804 0 _0283_
rlabel via2 15778 12835 15778 12835 0 _0284_
rlabel metal1 17066 14008 17066 14008 0 _0285_
rlabel metal1 13984 15130 13984 15130 0 _0286_
rlabel metal1 13432 10234 13432 10234 0 _0287_
rlabel metal2 18078 9384 18078 9384 0 _0288_
rlabel metal1 16192 10234 16192 10234 0 _0289_
rlabel metal1 14582 12852 14582 12852 0 _0290_
rlabel metal2 15042 9044 15042 9044 0 _0291_
rlabel metal1 17066 10540 17066 10540 0 _0292_
rlabel metal2 12926 13668 12926 13668 0 _0293_
rlabel metal2 20102 19550 20102 19550 0 _0294_
rlabel metal1 18446 17068 18446 17068 0 _0295_
rlabel metal1 20102 12954 20102 12954 0 _0296_
rlabel metal1 20332 18666 20332 18666 0 _0297_
rlabel metal2 16238 15334 16238 15334 0 _0298_
rlabel metal1 19182 12750 19182 12750 0 _0299_
rlabel metal1 4140 10098 4140 10098 0 _0300_
rlabel metal2 4094 14076 4094 14076 0 _0301_
rlabel metal2 1702 12517 1702 12517 0 _0302_
rlabel metal2 4830 11220 4830 11220 0 _0303_
rlabel metal2 24610 11560 24610 11560 0 _0304_
rlabel metal1 23782 13838 23782 13838 0 _0305_
rlabel metal1 22678 12886 22678 12886 0 _0306_
rlabel metal2 22494 14076 22494 14076 0 _0307_
rlabel metal2 20838 10948 20838 10948 0 _0308_
rlabel metal2 17526 19890 17526 19890 0 _0309_
rlabel metal1 20240 10778 20240 10778 0 _0310_
rlabel metal1 17342 18802 17342 18802 0 _0311_
rlabel metal1 7176 17850 7176 17850 0 _0312_
rlabel metal1 6394 9894 6394 9894 0 _0313_
rlabel metal1 8142 16150 8142 16150 0 _0314_
rlabel metal1 10212 14042 10212 14042 0 _0315_
rlabel metal1 16468 5338 16468 5338 0 _0316_
rlabel metal1 13340 4658 13340 4658 0 _0317_
rlabel metal1 14628 4522 14628 4522 0 _0318_
rlabel metal1 11270 7310 11270 7310 0 _0319_
rlabel metal1 10350 17544 10350 17544 0 _0320_
rlabel metal1 14490 9996 14490 9996 0 _0321_
rlabel metal2 9338 15912 9338 15912 0 _0322_
rlabel metal1 12604 8058 12604 8058 0 _0323_
rlabel metal2 17434 8296 17434 8296 0 _0324_
rlabel metal1 15686 6766 15686 6766 0 _0325_
rlabel metal1 13800 5610 13800 5610 0 _0326_
rlabel metal1 15502 4726 15502 4726 0 _0327_
rlabel metal1 8096 13498 8096 13498 0 _0328_
rlabel metal1 13524 16082 13524 16082 0 _0329_
rlabel metal1 9292 14042 9292 14042 0 _0330_
rlabel metal1 11086 15538 11086 15538 0 _0331_
rlabel metal1 10672 3094 10672 3094 0 _0332_
rlabel metal2 13386 11492 13386 11492 0 _0333_
rlabel metal2 11086 4556 11086 4556 0 _0334_
rlabel metal1 10258 10132 10258 10132 0 _0335_
rlabel metal2 16882 19584 16882 19584 0 _0336_
rlabel metal1 12558 20332 12558 20332 0 _0337_
rlabel metal2 17250 20026 17250 20026 0 _0338_
rlabel metal2 12834 19482 12834 19482 0 _0339_
rlabel metal1 22954 6970 22954 6970 0 _0340_
rlabel metal1 20608 8058 20608 8058 0 _0341_
rlabel metal2 22218 7582 22218 7582 0 _0342_
rlabel metal2 21022 7004 21022 7004 0 _0343_
rlabel metal1 20102 24072 20102 24072 0 _0344_
rlabel metal1 19642 23188 19642 23188 0 _0345_
rlabel metal1 19458 23766 19458 23766 0 _0346_
rlabel metal2 18170 24548 18170 24548 0 _0347_
rlabel metal2 8970 20604 8970 20604 0 _0348_
rlabel metal2 10994 21420 10994 21420 0 _0349_
rlabel metal2 9798 21148 9798 21148 0 _0350_
rlabel metal1 11500 21454 11500 21454 0 _0351_
rlabel metal1 14490 17000 14490 17000 0 _0352_
rlabel metal1 16146 7514 16146 7514 0 _0353_
rlabel metal1 15088 15674 15088 15674 0 _0354_
rlabel metal2 16974 7684 16974 7684 0 _0355_
rlabel metal2 17250 23902 17250 23902 0 _0356_
rlabel metal1 20608 22202 20608 22202 0 _0357_
rlabel metal2 17526 23528 17526 23528 0 _0358_
rlabel metal1 20424 22746 20424 22746 0 _0359_
rlabel metal1 22379 20842 22379 20842 0 _0360_
rlabel metal1 23322 17714 23322 17714 0 _0361_
rlabel metal1 22724 19482 22724 19482 0 _0362_
rlabel metal1 23046 17850 23046 17850 0 _0363_
rlabel metal2 4738 17374 4738 17374 0 _0364_
rlabel metal1 5014 15334 5014 15334 0 _0365_
rlabel metal2 5382 14552 5382 14552 0 _0366_
rlabel metal1 4416 14450 4416 14450 0 _0367_
rlabel metal1 16514 16966 16514 16966 0 _0368_
rlabel metal1 15824 12138 15824 12138 0 _0369_
rlabel metal1 18906 14586 18906 14586 0 _0370_
rlabel metal1 15272 5338 15272 5338 0 _0371_
rlabel metal1 7176 37298 7176 37298 0 ccff_head
rlabel metal1 4048 37094 4048 37094 0 ccff_tail
rlabel metal3 1234 27948 1234 27948 0 chanx_right_in[0]
rlabel metal2 38318 11679 38318 11679 0 chanx_right_in[10]
rlabel via2 38318 25245 38318 25245 0 chanx_right_in[11]
rlabel metal1 22724 37230 22724 37230 0 chanx_right_in[12]
rlabel metal2 10258 3604 10258 3604 0 chanx_right_in[13]
rlabel metal2 15502 1078 15502 1078 0 chanx_right_in[14]
rlabel metal2 32246 1588 32246 1588 0 chanx_right_in[15]
rlabel metal3 12136 1428 12136 1428 0 chanx_right_in[16]
rlabel metal2 38318 31569 38318 31569 0 chanx_right_in[17]
rlabel metal2 4554 891 4554 891 0 chanx_right_in[18]
rlabel metal2 34178 1588 34178 1588 0 chanx_right_in[1]
rlabel metal3 1234 32708 1234 32708 0 chanx_right_in[2]
rlabel metal1 33672 37230 33672 37230 0 chanx_right_in[3]
rlabel via2 38318 19805 38318 19805 0 chanx_right_in[4]
rlabel metal1 11776 37230 11776 37230 0 chanx_right_in[5]
rlabel metal3 1924 37468 1924 37468 0 chanx_right_in[6]
rlabel metal3 1234 25908 1234 25908 0 chanx_right_in[7]
rlabel metal2 38686 1554 38686 1554 0 chanx_right_in[8]
rlabel metal3 1234 17748 1234 17748 0 chanx_right_in[9]
rlabel metal2 38226 34833 38226 34833 0 chanx_right_out[0]
rlabel via2 38226 5525 38226 5525 0 chanx_right_out[10]
rlabel metal1 25944 37094 25944 37094 0 chanx_right_out[11]
rlabel metal3 1234 21148 1234 21148 0 chanx_right_out[12]
rlabel metal1 14996 37094 14996 37094 0 chanx_right_out[13]
rlabel metal1 16836 37094 16836 37094 0 chanx_right_out[14]
rlabel metal1 29486 37094 29486 37094 0 chanx_right_out[15]
rlabel metal3 1234 29308 1234 29308 0 chanx_right_out[16]
rlabel metal1 38272 36890 38272 36890 0 chanx_right_out[17]
rlabel via2 38226 33371 38226 33371 0 chanx_right_out[18]
rlabel metal2 38226 36941 38226 36941 0 chanx_right_out[1]
rlabel metal2 38226 8857 38226 8857 0 chanx_right_out[2]
rlabel metal1 24334 37094 24334 37094 0 chanx_right_out[3]
rlabel metal1 18216 37094 18216 37094 0 chanx_right_out[4]
rlabel metal3 1234 4828 1234 4828 0 chanx_right_out[5]
rlabel metal1 1794 37128 1794 37128 0 chanx_right_out[6]
rlabel metal1 9200 4454 9200 4454 0 chanx_right_out[7]
rlabel metal2 38226 28815 38226 28815 0 chanx_right_out[8]
rlabel metal2 37398 1520 37398 1520 0 chanx_right_out[9]
rlabel metal2 38318 15249 38318 15249 0 chany_top_in[0]
rlabel metal1 20838 37230 20838 37230 0 chany_top_in[10]
rlabel metal1 13064 37230 13064 37230 0 chany_top_in[11]
rlabel metal1 37122 3026 37122 3026 0 chany_top_in[12]
rlabel metal2 38318 30107 38318 30107 0 chany_top_in[13]
rlabel metal1 38180 36142 38180 36142 0 chany_top_in[14]
rlabel via3 3243 15300 3243 15300 0 chany_top_in[15]
rlabel metal2 13570 1163 13570 1163 0 chany_top_in[16]
rlabel metal3 38786 6868 38786 6868 0 chany_top_in[17]
rlabel metal3 1234 22508 1234 22508 0 chany_top_in[18]
rlabel metal3 1717 2788 1717 2788 0 chany_top_in[1]
rlabel metal3 1234 30668 1234 30668 0 chany_top_in[2]
rlabel metal1 10488 37230 10488 37230 0 chany_top_in[3]
rlabel metal2 29026 1588 29026 1588 0 chany_top_in[4]
rlabel metal1 34960 37230 34960 37230 0 chany_top_in[5]
rlabel metal2 24518 1588 24518 1588 0 chany_top_in[6]
rlabel metal2 2622 2132 2622 2132 0 chany_top_in[7]
rlabel metal3 1234 19788 1234 19788 0 chany_top_in[8]
rlabel metal2 35466 1588 35466 1588 0 chany_top_in[9]
rlabel via2 38226 17051 38226 17051 0 chany_top_out[0]
rlabel metal2 38226 10353 38226 10353 0 chany_top_out[10]
rlabel metal2 27738 1520 27738 1520 0 chany_top_out[11]
rlabel metal3 1234 34068 1234 34068 0 chany_top_out[12]
rlabel metal2 38226 2465 38226 2465 0 chany_top_out[13]
rlabel metal1 5336 37094 5336 37094 0 chany_top_out[14]
rlabel via2 38226 13685 38226 13685 0 chany_top_out[15]
rlabel via2 1794 16405 1794 16405 0 chany_top_out[16]
rlabel metal2 30958 1520 30958 1520 0 chany_top_out[17]
rlabel metal2 38226 26673 38226 26673 0 chany_top_out[18]
rlabel metal2 18722 1520 18722 1520 0 chany_top_out[1]
rlabel metal3 1234 24548 1234 24548 0 chany_top_out[2]
rlabel metal2 20010 1520 20010 1520 0 chany_top_out[3]
rlabel metal2 46 1044 46 1044 0 chany_top_out[4]
rlabel metal2 23230 1520 23230 1520 0 chany_top_out[5]
rlabel via2 3726 8245 3726 8245 0 chany_top_out[6]
rlabel metal1 19504 37094 19504 37094 0 chany_top_out[7]
rlabel metal3 1234 12988 1234 12988 0 chany_top_out[8]
rlabel metal1 1242 36890 1242 36890 0 chany_top_out[9]
rlabel metal1 15042 20468 15042 20468 0 mem_right_track_0.DFFR_0_.D
rlabel metal2 8050 3876 8050 3876 0 mem_right_track_0.DFFR_0_.Q
rlabel metal1 13524 5134 13524 5134 0 mem_right_track_0.DFFR_1_.Q
rlabel metal1 14214 22542 14214 22542 0 mem_right_track_10.DFFR_0_.D
rlabel metal1 22494 16082 22494 16082 0 mem_right_track_10.DFFR_0_.Q
rlabel metal2 13478 7072 13478 7072 0 mem_right_track_10.DFFR_1_.Q
rlabel metal2 21758 18496 21758 18496 0 mem_right_track_12.DFFR_0_.Q
rlabel metal2 10902 2244 10902 2244 0 mem_right_track_12.DFFR_1_.Q
rlabel metal1 8418 8840 8418 8840 0 mem_right_track_14.DFFR_0_.Q
rlabel metal2 9614 8177 9614 8177 0 mem_right_track_14.DFFR_1_.Q
rlabel metal1 13110 14348 13110 14348 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 13754 14382 13754 14382 0 mem_right_track_16.DFFR_1_.Q
rlabel metal2 9706 7021 9706 7021 0 mem_right_track_18.DFFR_0_.Q
rlabel metal1 1978 12104 1978 12104 0 mem_right_track_18.DFFR_1_.Q
rlabel metal1 23920 17170 23920 17170 0 mem_right_track_2.DFFR_0_.Q
rlabel metal2 23598 18751 23598 18751 0 mem_right_track_2.DFFR_1_.Q
rlabel metal2 20102 8738 20102 8738 0 mem_right_track_20.DFFR_0_.Q
rlabel metal2 20838 8653 20838 8653 0 mem_right_track_20.DFFR_1_.Q
rlabel metal1 16882 23120 16882 23120 0 mem_right_track_22.DFFR_0_.Q
rlabel metal2 18538 23647 18538 23647 0 mem_right_track_22.DFFR_1_.Q
rlabel metal2 13478 8653 13478 8653 0 mem_right_track_24.DFFR_0_.Q
rlabel metal1 9890 21522 9890 21522 0 mem_right_track_24.DFFR_1_.Q
rlabel metal1 16836 7378 16836 7378 0 mem_right_track_26.DFFR_0_.Q
rlabel metal1 13846 15470 13846 15470 0 mem_right_track_26.DFFR_1_.Q
rlabel metal2 19826 22372 19826 22372 0 mem_right_track_28.DFFR_0_.Q
rlabel metal1 16330 23664 16330 23664 0 mem_right_track_28.DFFR_1_.Q
rlabel via2 23322 17187 23322 17187 0 mem_right_track_30.DFFR_0_.Q
rlabel metal1 22494 19380 22494 19380 0 mem_right_track_30.DFFR_1_.Q
rlabel metal1 4232 2618 4232 2618 0 mem_right_track_32.DFFR_0_.Q
rlabel metal1 5750 14960 5750 14960 0 mem_right_track_32.DFFR_1_.Q
rlabel metal2 9614 2006 9614 2006 0 mem_right_track_34.DFFR_0_.Q
rlabel metal2 17618 14484 17618 14484 0 mem_right_track_34.DFFR_1_.Q
rlabel metal1 16238 14994 16238 14994 0 mem_right_track_36.DFFR_0_.Q
rlabel metal2 14582 1870 14582 1870 0 mem_right_track_4.DFFR_0_.Q
rlabel metal1 17296 2278 17296 2278 0 mem_right_track_4.DFFR_1_.Q
rlabel metal1 12006 23052 12006 23052 0 mem_right_track_6.DFFR_0_.Q
rlabel metal2 14490 16252 14490 16252 0 mem_right_track_6.DFFR_1_.Q
rlabel metal2 13570 19788 13570 19788 0 mem_right_track_8.DFFR_0_.Q
rlabel metal1 22218 12716 22218 12716 0 mem_top_track_0.DFFR_0_.Q
rlabel via2 3358 9061 3358 9061 0 mem_top_track_0.DFFR_1_.Q
rlabel metal1 8510 14926 8510 14926 0 mem_top_track_10.DFFR_0_.D
rlabel metal1 8418 18802 8418 18802 0 mem_top_track_10.DFFR_0_.Q
rlabel metal2 12742 6239 12742 6239 0 mem_top_track_10.DFFR_1_.Q
rlabel metal1 7268 13906 7268 13906 0 mem_top_track_12.DFFR_0_.Q
rlabel metal2 13478 6375 13478 6375 0 mem_top_track_12.DFFR_1_.Q
rlabel metal2 9982 7616 9982 7616 0 mem_top_track_14.DFFR_0_.Q
rlabel metal2 12006 13226 12006 13226 0 mem_top_track_14.DFFR_1_.Q
rlabel metal1 2024 13974 2024 13974 0 mem_top_track_16.DFFR_0_.Q
rlabel metal1 1610 10676 1610 10676 0 mem_top_track_16.DFFR_1_.Q
rlabel metal2 22586 14093 22586 14093 0 mem_top_track_18.DFFR_0_.Q
rlabel metal1 13708 16558 13708 16558 0 mem_top_track_18.DFFR_1_.Q
rlabel metal1 8188 19346 8188 19346 0 mem_top_track_2.DFFR_0_.Q
rlabel metal2 14858 11169 14858 11169 0 mem_top_track_2.DFFR_1_.Q
rlabel metal1 23230 14450 23230 14450 0 mem_top_track_20.DFFR_0_.Q
rlabel metal2 12466 13260 12466 13260 0 mem_top_track_20.DFFR_1_.Q
rlabel metal1 7314 12886 7314 12886 0 mem_top_track_22.DFFR_0_.Q
rlabel metal2 20378 10336 20378 10336 0 mem_top_track_22.DFFR_1_.Q
rlabel metal1 6854 14348 6854 14348 0 mem_top_track_24.DFFR_0_.Q
rlabel metal1 7774 16082 7774 16082 0 mem_top_track_24.DFFR_1_.Q
rlabel metal1 18216 7786 18216 7786 0 mem_top_track_26.DFFR_0_.Q
rlabel metal2 1886 7752 1886 7752 0 mem_top_track_26.DFFR_1_.Q
rlabel metal1 9292 8942 9292 8942 0 mem_top_track_28.DFFR_0_.Q
rlabel metal1 9522 15470 9522 15470 0 mem_top_track_28.DFFR_1_.Q
rlabel metal3 9016 9860 9016 9860 0 mem_top_track_30.DFFR_0_.Q
rlabel metal2 16330 6511 16330 6511 0 mem_top_track_30.DFFR_1_.Q
rlabel metal3 6026 13124 6026 13124 0 mem_top_track_32.DFFR_0_.Q
rlabel metal1 8832 13906 8832 13906 0 mem_top_track_32.DFFR_1_.Q
rlabel metal2 9522 13124 9522 13124 0 mem_top_track_34.DFFR_0_.Q
rlabel metal1 6624 13362 6624 13362 0 mem_top_track_34.DFFR_1_.Q
rlabel metal1 11592 19822 11592 19822 0 mem_top_track_36.DFFR_0_.Q
rlabel metal1 17388 18734 17388 18734 0 mem_top_track_4.DFFR_0_.Q
rlabel metal1 12926 20876 12926 20876 0 mem_top_track_4.DFFR_1_.Q
rlabel metal2 20746 14722 20746 14722 0 mem_top_track_6.DFFR_0_.Q
rlabel metal1 10948 4522 10948 4522 0 mem_top_track_6.DFFR_1_.Q
rlabel metal1 8832 17170 8832 17170 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 11454 19346 11454 19346 0 mux_right_track_0.INVTX1_0_.out
rlabel metal2 12558 8109 12558 8109 0 mux_right_track_0.INVTX1_1_.out
rlabel metal2 22034 17034 22034 17034 0 mux_right_track_0.INVTX1_2_.out
rlabel metal1 15456 18190 15456 18190 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16974 18020 16974 18020 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 29716 26350 29716 26350 0 mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 29946 26554 29946 26554 0 mux_right_track_0.out
rlabel metal1 23414 9010 23414 9010 0 mux_right_track_10.INVTX1_0_.out
rlabel metal1 19780 21454 19780 21454 0 mux_right_track_10.INVTX1_1_.out
rlabel metal1 22218 17782 22218 17782 0 mux_right_track_10.INVTX1_2_.out
rlabel metal1 21620 20366 21620 20366 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 19550 11356 19550 11356 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 1886 11730 1886 11730 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 2024 16082 2024 16082 0 mux_right_track_10.out
rlabel metal2 30590 26894 30590 26894 0 mux_right_track_12.INVTX1_0_.out
rlabel metal1 13110 9044 13110 9044 0 mux_right_track_12.INVTX1_2_.out
rlabel metal1 20332 18598 20332 18598 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13800 17850 13800 17850 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 2438 27999 2438 27999 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 2530 36278 2530 36278 0 mux_right_track_12.out
rlabel metal1 19803 6834 19803 6834 0 mux_right_track_14.INVTX1_0_.out
rlabel metal2 31602 17374 31602 17374 0 mux_right_track_14.INVTX1_2_.out
rlabel metal1 14674 7854 14674 7854 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16836 12614 16836 12614 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15778 7718 15778 7718 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 17342 5202 17342 5202 0 mux_right_track_14.out
rlabel metal1 12880 11118 12880 11118 0 mux_right_track_16.INVTX1_0_.out
rlabel metal1 13524 9350 13524 9350 0 mux_right_track_16.INVTX1_2_.out
rlabel metal1 16376 12954 16376 12954 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17204 15674 17204 15674 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 28842 17476 28842 17476 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30498 21114 30498 21114 0 mux_right_track_16.out
rlabel metal2 12466 14892 12466 14892 0 mux_right_track_18.INVTX1_0_.out
rlabel metal1 15180 12954 15180 12954 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17250 10744 17250 10744 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 28290 8942 28290 8942 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 32119 5202 32119 5202 0 mux_right_track_18.out
rlabel metal1 22126 15980 22126 15980 0 mux_right_track_2.INVTX1_0_.out
rlabel metal2 29854 27302 29854 27302 0 mux_right_track_2.INVTX1_2_.out
rlabel metal1 22862 17306 22862 17306 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22862 20128 22862 20128 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 23690 19040 23690 19040 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 29900 28730 29900 28730 0 mux_right_track_2.out
rlabel metal1 20838 6732 20838 6732 0 mux_right_track_20.INVTX1_0_.out
rlabel metal2 22126 7820 22126 7820 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 26772 7310 26772 7310 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 29670 5882 29670 5882 0 mux_right_track_20.out
rlabel metal1 19550 34510 19550 34510 0 mux_right_track_22.INVTX1_0_.out
rlabel metal1 19596 23630 19596 23630 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 20654 26928 20654 26928 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 22724 35054 22724 35054 0 mux_right_track_22.out
rlabel metal1 11960 34918 11960 34918 0 mux_right_track_24.INVTX1_0_.out
rlabel metal1 21068 32198 21068 32198 0 mux_right_track_24.INVTX1_1_.out
rlabel metal1 10626 21046 10626 21046 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9108 20298 9108 20298 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 5520 20434 5520 20434 0 mux_right_track_24.out
rlabel metal2 33902 7735 33902 7735 0 mux_right_track_26.INVTX1_0_.out
rlabel metal1 15686 20910 15686 20910 0 mux_right_track_26.INVTX1_1_.out
rlabel metal1 16468 16626 16468 16626 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16054 17204 16054 17204 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15502 35054 15502 35054 0 mux_right_track_26.out
rlabel metal2 20746 25228 20746 25228 0 mux_right_track_28.INVTX1_0_.out
rlabel metal1 20562 23222 20562 23222 0 mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17434 27166 17434 27166 0 mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17020 30906 17020 30906 0 mux_right_track_28.out
rlabel metal1 23506 18224 23506 18224 0 mux_right_track_30.INVTX1_0_.out
rlabel metal1 22816 18054 22816 18054 0 mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 23230 20434 23230 20434 0 mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 27370 34374 27370 34374 0 mux_right_track_30.out
rlabel metal2 2714 14926 2714 14926 0 mux_right_track_32.INVTX1_0_.out
rlabel metal1 4968 14314 4968 14314 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 4876 17102 4876 17102 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 4462 25874 4462 25874 0 mux_right_track_32.out
rlabel metal1 14582 7310 14582 7310 0 mux_right_track_34.INVTX1_0_.out
rlabel metal1 19044 16626 19044 16626 0 mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 29118 23358 29118 23358 0 mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 29670 29274 29670 29274 0 mux_right_track_34.out
rlabel metal1 19136 10166 19136 10166 0 mux_right_track_36.INVTX1_0_.out
rlabel metal1 19642 14858 19642 14858 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19504 17238 19504 17238 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 28750 22236 28750 22236 0 mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 31786 25466 31786 25466 0 mux_right_track_36.out
rlabel metal2 11362 12801 11362 12801 0 mux_right_track_4.INVTX1_0_.out
rlabel metal1 19964 13362 19964 13362 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19734 17306 19734 17306 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 20102 13940 20102 13940 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 36478 11356 36478 11356 0 mux_right_track_4.out
rlabel metal1 10258 22610 10258 22610 0 mux_right_track_6.INVTX1_0_.out
rlabel metal1 13846 22066 13846 22066 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16146 21522 16146 21522 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15824 22066 15824 22066 0 mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 20654 35054 20654 35054 0 mux_right_track_6.out
rlabel metal1 12144 34510 12144 34510 0 mux_right_track_8.INVTX1_0_.out
rlabel metal1 14904 21386 14904 21386 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19412 21658 19412 21658 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 17618 26146 17618 26146 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 17434 29818 17434 29818 0 mux_right_track_8.out
rlabel metal1 20654 16660 20654 16660 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 20332 13838 20332 13838 0 mux_top_track_0.INVTX1_1_.out
rlabel metal2 29578 8738 29578 8738 0 mux_top_track_0.INVTX1_2_.out
rlabel metal2 22402 14008 22402 14008 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23414 12308 23414 12308 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23322 13362 23322 13362 0 mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30222 14586 30222 14586 0 mux_top_track_0.out
rlabel metal1 9292 31790 9292 31790 0 mux_top_track_10.INVTX1_0_.out
rlabel via1 13110 6749 13110 6749 0 mux_top_track_10.INVTX1_1_.out
rlabel metal1 7590 18666 7590 18666 0 mux_top_track_10.INVTX1_2_.out
rlabel metal1 12604 13158 12604 13158 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel via1 12558 18581 12558 18581 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 13248 12750 13248 12750 0 mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 18814 6970 18814 6970 0 mux_top_track_10.out
rlabel metal1 8740 12750 8740 12750 0 mux_top_track_12.INVTX1_1_.out
rlabel metal2 6302 19006 6302 19006 0 mux_top_track_12.INVTX1_2_.out
rlabel metal1 9476 12614 9476 12614 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 7360 16966 7360 16966 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 6624 15470 6624 15470 0 mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 4646 15028 4646 15028 0 mux_top_track_12.out
rlabel metal3 4025 29036 4025 29036 0 mux_top_track_14.INVTX1_1_.out
rlabel metal2 21482 6426 21482 6426 0 mux_top_track_14.INVTX1_2_.out
rlabel metal1 12006 14994 12006 14994 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 18630 13906 18630 13906 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17342 14450 17342 14450 0 mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 18308 29274 18308 29274 0 mux_top_track_14.out
rlabel metal2 1978 14314 1978 14314 0 mux_top_track_16.INVTX1_1_.out
rlabel metal1 4830 13702 4830 13702 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 6900 12614 6900 12614 0 mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 3450 15470 3450 15470 0 mux_top_track_16.out
rlabel metal1 22494 16626 22494 16626 0 mux_top_track_18.INVTX1_1_.out
rlabel metal1 23230 14960 23230 14960 0 mux_top_track_18.INVTX1_2_.out
rlabel metal1 21114 16422 21114 16422 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20516 15606 20516 15606 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 7130 33184 7130 33184 0 mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 7222 34612 7222 34612 0 mux_top_track_18.out
rlabel metal1 22264 31926 22264 31926 0 mux_top_track_2.INVTX1_1_.out
rlabel metal1 8786 20026 8786 20026 0 mux_top_track_2.INVTX1_2_.out
rlabel metal1 18584 14042 18584 14042 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13938 18054 13938 18054 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15732 13498 15732 13498 0 mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 16882 3026 16882 3026 0 mux_top_track_2.out
rlabel metal1 24334 13872 24334 13872 0 mux_top_track_20.INVTX1_1_.out
rlabel metal1 23184 12750 23184 12750 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24242 11594 24242 11594 0 mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 30866 10846 30866 10846 0 mux_top_track_20.out
rlabel metal1 20700 20570 20700 20570 0 mux_top_track_22.INVTX1_1_.out
rlabel metal1 19596 18870 19596 18870 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20976 10982 20976 10982 0 mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 24794 8092 24794 8092 0 mux_top_track_22.out
rlabel metal2 25254 26044 25254 26044 0 mux_top_track_24.INVTX1_0_.out
rlabel metal1 9384 12274 9384 12274 0 mux_top_track_24.INVTX1_1_.out
rlabel metal1 10902 15674 10902 15674 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 6854 29614 6854 29614 0 mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 6118 30260 6118 30260 0 mux_top_track_24.out
rlabel metal1 8694 31790 8694 31790 0 mux_top_track_26.INVTX1_0_.out
rlabel metal1 13110 4556 13110 4556 0 mux_top_track_26.INVTX1_1_.out
rlabel metal1 13478 4590 13478 4590 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 36685 5202 36685 5202 0 mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 37950 5202 37950 5202 0 mux_top_track_26.out
rlabel metal2 18354 8840 18354 8840 0 mux_top_track_28.INVTX1_1_.out
rlabel metal2 14674 11220 14674 11220 0 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 10350 31790 10350 31790 0 mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 9890 33286 9890 33286 0 mux_top_track_28.out
rlabel metal2 14214 9911 14214 9911 0 mux_top_track_30.INVTX1_1_.out
rlabel metal1 14352 6630 14352 6630 0 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 24886 9622 24886 9622 0 mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 28842 10778 28842 10778 0 mux_top_track_30.out
rlabel metal2 32430 21726 32430 21726 0 mux_top_track_32.INVTX1_1_.out
rlabel metal1 12926 15674 12926 15674 0 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 8602 14620 8602 14620 0 mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 5198 13940 5198 13940 0 mux_top_track_32.out
rlabel metal1 12190 11798 12190 11798 0 mux_top_track_34.INVTX1_1_.out
rlabel metal1 13570 9894 13570 9894 0 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 19826 3842 19826 3842 0 mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 26726 3910 26726 3910 0 mux_top_track_34.out
rlabel metal1 8740 23494 8740 23494 0 mux_top_track_36.INVTX1_1_.out
rlabel metal1 15502 19482 15502 19482 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 24886 20842 24886 20842 0 mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 30084 22066 30084 22066 0 mux_top_track_36.out
rlabel metal2 29854 33728 29854 33728 0 mux_top_track_4.INVTX1_2_.out
rlabel metal1 16422 20842 16422 20842 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17940 21386 17940 21386 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15640 20230 15640 20230 0 mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6946 22610 6946 22610 0 mux_top_track_4.out
rlabel metal2 23138 15708 23138 15708 0 mux_top_track_6.INVTX1_2_.out
rlabel metal1 14766 15334 14766 15334 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20332 15130 20332 15130 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17756 13498 17756 13498 0 mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 17526 4114 17526 4114 0 mux_top_track_6.out
rlabel metal1 10534 33286 10534 33286 0 mux_top_track_8.INVTX1_2_.out
rlabel metal1 9752 16422 9752 16422 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9246 19686 9246 19686 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 2530 14348 2530 14348 0 mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 2162 17646 2162 17646 0 mux_top_track_8.out
rlabel metal3 7567 36516 7567 36516 0 net1
rlabel metal2 37030 29988 37030 29988 0 net10
rlabel metal1 23736 11186 23736 11186 0 net100
rlabel metal2 11270 18700 11270 18700 0 net101
rlabel metal1 18446 21556 18446 21556 0 net102
rlabel metal1 19044 14926 19044 14926 0 net103
rlabel metal2 9890 20094 9890 20094 0 net104
rlabel metal2 9706 18530 9706 18530 0 net105
rlabel metal1 7084 17102 7084 17102 0 net106
rlabel metal1 18308 12274 18308 12274 0 net107
rlabel metal1 21666 15538 21666 15538 0 net108
rlabel metal1 15042 17306 15042 17306 0 net109
rlabel metal2 20562 9707 20562 9707 0 net11
rlabel metal1 22494 20468 22494 20468 0 net110
rlabel metal1 19044 16558 19044 16558 0 net111
rlabel metal1 15640 19822 15640 19822 0 net112
rlabel metal1 18722 22542 18722 22542 0 net113
rlabel metal2 19458 11254 19458 11254 0 net114
rlabel metal2 14306 19278 14306 19278 0 net115
rlabel metal1 16790 12750 16790 12750 0 net116
rlabel metal1 16054 14450 16054 14450 0 net117
rlabel metal1 16422 10098 16422 10098 0 net118
rlabel metal1 18262 17204 18262 17204 0 net119
rlabel metal1 34822 2618 34822 2618 0 net12
rlabel metal1 3910 16014 3910 16014 0 net120
rlabel metal1 24472 11662 24472 11662 0 net121
rlabel metal1 20746 11186 20746 11186 0 net122
rlabel metal2 7130 18462 7130 18462 0 net123
rlabel metal2 16514 5984 16514 5984 0 net124
rlabel metal1 10304 17306 10304 17306 0 net125
rlabel metal2 17342 8670 17342 8670 0 net126
rlabel metal1 8050 14042 8050 14042 0 net127
rlabel metal1 10442 3094 10442 3094 0 net128
rlabel metal2 18170 19618 18170 19618 0 net129
rlabel metal2 5566 30634 5566 30634 0 net13
rlabel metal2 23322 7582 23322 7582 0 net130
rlabel metal2 20010 24480 20010 24480 0 net131
rlabel metal2 8786 20944 8786 20944 0 net132
rlabel metal2 15410 18734 15410 18734 0 net133
rlabel metal2 17158 24242 17158 24242 0 net134
rlabel metal2 22586 21216 22586 21216 0 net135
rlabel metal1 4692 16626 4692 16626 0 net136
rlabel metal2 21206 16966 21206 16966 0 net137
rlabel metal1 31694 36890 31694 36890 0 net14
rlabel metal2 37030 19210 37030 19210 0 net15
rlabel metal1 11270 37094 11270 37094 0 net16
rlabel metal1 4784 37162 4784 37162 0 net17
rlabel metal1 3358 26486 3358 26486 0 net18
rlabel metal2 35650 2448 35650 2448 0 net19
rlabel metal1 2760 27846 2760 27846 0 net2
rlabel metal1 1748 14994 1748 14994 0 net20
rlabel metal2 38134 15878 38134 15878 0 net21
rlabel metal1 20332 34578 20332 34578 0 net22
rlabel metal1 12558 35054 12558 35054 0 net23
rlabel metal1 36248 3162 36248 3162 0 net24
rlabel metal2 34178 28730 34178 28730 0 net25
rlabel metal1 36340 36006 36340 36006 0 net26
rlabel metal1 2530 15470 2530 15470 0 net27
rlabel metal1 15594 7378 15594 7378 0 net28
rlabel metal1 37536 7514 37536 7514 0 net29
rlabel metal2 34638 12580 34638 12580 0 net3
rlabel metal1 3588 22406 3588 22406 0 net30
rlabel metal1 19458 12784 19458 12784 0 net31
rlabel metal2 3818 29002 3818 29002 0 net32
rlabel metal1 11224 37162 11224 37162 0 net33
rlabel metal1 29118 2618 29118 2618 0 net34
rlabel metal1 33396 37162 33396 37162 0 net35
rlabel metal1 21114 6834 21114 6834 0 net36
rlabel metal2 12604 10676 12604 10676 0 net37
rlabel metal2 5566 18156 5566 18156 0 net38
rlabel metal1 35006 2550 35006 2550 0 net39
rlabel metal2 34638 23324 34638 23324 0 net4
rlabel metal2 20838 2074 20838 2074 0 net40
rlabel metal1 36340 37094 36340 37094 0 net41
rlabel metal1 25208 32402 25208 32402 0 net42
rlabel metal1 16330 2550 16330 2550 0 net43
rlabel metal2 36754 33932 36754 33932 0 net44
rlabel metal2 31418 8262 31418 8262 0 net45
rlabel metal1 5520 8466 5520 8466 0 net46
rlabel metal2 38134 19788 38134 19788 0 net47
rlabel metal2 12834 7497 12834 7497 0 net48
rlabel metal2 19458 2193 19458 2193 0 net49
rlabel metal1 22218 37094 22218 37094 0 net5
rlabel metal2 7130 14450 7130 14450 0 net50
rlabel metal2 34546 22508 34546 22508 0 net51
rlabel metal1 21160 2618 21160 2618 0 net52
rlabel metal1 29302 31892 29302 31892 0 net53
rlabel metal1 25162 31824 25162 31824 0 net54
rlabel metal1 4186 36890 4186 36890 0 net55
rlabel metal2 9154 34442 9154 34442 0 net56
rlabel metal1 25714 2618 25714 2618 0 net57
rlabel metal1 4922 8058 4922 8058 0 net58
rlabel metal1 2162 36006 2162 36006 0 net59
rlabel metal1 8096 4794 8096 4794 0 net6
rlabel metal2 34546 18122 34546 18122 0 net60
rlabel metal1 18354 19822 18354 19822 0 net61
rlabel metal1 35190 30906 35190 30906 0 net62
rlabel metal1 36961 5678 36961 5678 0 net63
rlabel metal1 25300 37230 25300 37230 0 net64
rlabel metal1 5106 20570 5106 20570 0 net65
rlabel metal1 15042 35258 15042 35258 0 net66
rlabel metal2 16882 36244 16882 36244 0 net67
rlabel metal1 28796 37230 28796 37230 0 net68
rlabel metal1 4094 28968 4094 28968 0 net69
rlabel metal1 17158 2618 17158 2618 0 net7
rlabel metal1 38042 36720 38042 36720 0 net70
rlabel metal1 35144 29818 35144 29818 0 net71
rlabel metal1 38042 37196 38042 37196 0 net72
rlabel metal2 38042 9690 38042 9690 0 net73
rlabel metal1 23782 37230 23782 37230 0 net74
rlabel metal1 17802 35258 17802 35258 0 net75
rlabel metal1 1656 15878 1656 15878 0 net76
rlabel metal1 2116 36890 2116 36890 0 net77
rlabel metal2 15962 4896 15962 4896 0 net78
rlabel metal2 38042 26894 38042 26894 0 net79
rlabel metal1 31280 2618 31280 2618 0 net8
rlabel metal1 37490 2448 37490 2448 0 net80
rlabel metal1 36984 17170 36984 17170 0 net81
rlabel metal1 38042 10608 38042 10608 0 net82
rlabel metal1 27830 2448 27830 2448 0 net83
rlabel metal1 4140 30906 4140 30906 0 net84
rlabel metal2 38042 4012 38042 4012 0 net85
rlabel metal1 6026 37230 6026 37230 0 net86
rlabel metal2 34270 12886 34270 12886 0 net87
rlabel metal2 1702 15300 1702 15300 0 net88
rlabel metal1 31050 2448 31050 2448 0 net89
rlabel metal3 17204 3128 17204 3128 0 net9
rlabel metal2 34822 25398 34822 25398 0 net90
rlabel metal1 17756 2890 17756 2890 0 net91
rlabel metal2 5474 23766 5474 23766 0 net92
rlabel metal1 19688 2482 19688 2482 0 net93
rlabel metal1 1840 17510 1840 17510 0 net94
rlabel metal1 23322 2380 23322 2380 0 net95
rlabel metal2 4692 13158 4692 13158 0 net96
rlabel metal1 18906 34714 18906 34714 0 net97
rlabel metal1 1610 14416 1610 14416 0 net98
rlabel metal1 2852 36686 2852 36686 0 net99
rlabel metal2 20470 2108 20470 2108 0 pReset
rlabel metal2 1610 13600 1610 13600 0 prog_clk
rlabel metal1 36846 37230 36846 37230 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 27232 37230 27232 37230 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 16790 1588 16790 1588 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 36938 36788 36938 36788 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel via2 38318 3485 38318 3485 0 right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 3910 9095 3910 9095 0 right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 38318 21913 38318 21913 0 right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal1 7544 4590 7544 4590 0 right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 18814 2074 18814 2074 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal3 1234 14348 1234 14348 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 38318 23443 38318 23443 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 21298 1588 21298 1588 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 32154 37230 32154 37230 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 30544 37230 30544 37230 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 2254 37230 2254 37230 0 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 8878 37230 8878 37230 0 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 26450 1588 26450 1588 0 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 3634 9435 3634 9435 0 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal3 1234 36108 1234 36108 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 38318 18581 38318 18581 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
