magic
tech sky130A
magscale 1 2
timestamp 1672416659
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 1844 39362 37584
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 3238 39200 3294 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 14186 39200 14242 39800
rect 16118 39200 16174 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 23202 39200 23258 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 34150 39200 34206 39800
rect 36082 39200 36138 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 5170 200 5226 800
rect 7102 200 7158 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 12254 200 12310 800
rect 14186 200 14242 800
rect 16118 200 16174 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 23202 200 23258 800
rect 25134 200 25190 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 36082 200 36138 800
rect 38014 200 38070 800
rect 39302 200 39358 800
<< obsm2 >>
rect 130 39144 1250 39200
rect 1418 39144 3182 39200
rect 3350 39144 5114 39200
rect 5282 39144 7046 39200
rect 7214 39144 8978 39200
rect 9146 39144 10266 39200
rect 10434 39144 12198 39200
rect 12366 39144 14130 39200
rect 14298 39144 16062 39200
rect 16230 39144 17994 39200
rect 18162 39144 19926 39200
rect 20094 39144 21214 39200
rect 21382 39144 23146 39200
rect 23314 39144 25078 39200
rect 25246 39144 27010 39200
rect 27178 39144 28942 39200
rect 29110 39144 30230 39200
rect 30398 39144 32162 39200
rect 32330 39144 34094 39200
rect 34262 39144 36026 39200
rect 36194 39144 37958 39200
rect 38126 39144 39246 39200
rect 20 856 39356 39144
rect 130 734 1250 856
rect 1418 734 3182 856
rect 3350 734 5114 856
rect 5282 734 7046 856
rect 7214 734 8978 856
rect 9146 734 10266 856
rect 10434 734 12198 856
rect 12366 734 14130 856
rect 14298 734 16062 856
rect 16230 734 17994 856
rect 18162 734 19282 856
rect 19450 734 21214 856
rect 21382 734 23146 856
rect 23314 734 25078 856
rect 25246 734 27010 856
rect 27178 734 28942 856
rect 29110 734 30230 856
rect 30398 734 32162 856
rect 32330 734 34094 856
rect 34262 734 36026 856
rect 36194 734 37958 856
rect 38126 734 39246 856
<< metal3 >>
rect 200 38088 800 38208
rect 39200 38088 39800 38208
rect 200 36048 800 36168
rect 39200 36048 39800 36168
rect 200 34008 800 34128
rect 39200 34008 39800 34128
rect 200 31968 800 32088
rect 39200 31968 39800 32088
rect 200 30608 800 30728
rect 39200 29928 39800 30048
rect 200 28568 800 28688
rect 39200 28568 39800 28688
rect 200 26528 800 26648
rect 39200 26528 39800 26648
rect 200 24488 800 24608
rect 39200 24488 39800 24608
rect 200 22448 800 22568
rect 39200 22448 39800 22568
rect 200 20408 800 20528
rect 39200 20408 39800 20528
rect 200 19048 800 19168
rect 39200 19048 39800 19168
rect 200 17008 800 17128
rect 39200 17008 39800 17128
rect 200 14968 800 15088
rect 39200 14968 39800 15088
rect 200 12928 800 13048
rect 39200 12928 39800 13048
rect 200 10888 800 11008
rect 39200 10888 39800 11008
rect 200 9528 800 9648
rect 39200 8848 39800 8968
rect 200 7488 800 7608
rect 39200 7488 39800 7608
rect 200 5448 800 5568
rect 39200 5448 39800 5568
rect 200 3408 800 3528
rect 39200 3408 39800 3528
rect 200 1368 800 1488
rect 39200 1368 39800 1488
<< obsm3 >>
rect 880 38008 39120 38181
rect 800 36248 39200 38008
rect 880 35968 39120 36248
rect 800 34208 39200 35968
rect 880 33928 39120 34208
rect 800 32168 39200 33928
rect 880 31888 39120 32168
rect 800 30808 39200 31888
rect 880 30528 39200 30808
rect 800 30128 39200 30528
rect 800 29848 39120 30128
rect 800 28768 39200 29848
rect 880 28488 39120 28768
rect 800 26728 39200 28488
rect 880 26448 39120 26728
rect 800 24688 39200 26448
rect 880 24408 39120 24688
rect 800 22648 39200 24408
rect 880 22368 39120 22648
rect 800 20608 39200 22368
rect 880 20328 39120 20608
rect 800 19248 39200 20328
rect 880 18968 39120 19248
rect 800 17208 39200 18968
rect 880 16928 39120 17208
rect 800 15168 39200 16928
rect 880 14888 39120 15168
rect 800 13128 39200 14888
rect 880 12848 39120 13128
rect 800 11088 39200 12848
rect 880 10808 39120 11088
rect 800 9728 39200 10808
rect 880 9448 39200 9728
rect 800 9048 39200 9448
rect 800 8768 39120 9048
rect 800 7688 39200 8768
rect 880 7408 39120 7688
rect 800 5648 39200 7408
rect 880 5368 39120 5648
rect 800 3608 39200 5368
rect 880 3328 39120 3608
rect 800 1568 39200 3328
rect 880 1395 39120 1568
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 26371 7515 26437 23629
<< labels >>
rlabel metal3 s 39200 17008 39800 17128 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 39200 34008 39800 34128 6 ccff_tail
port 2 nsew signal output
rlabel metal2 s 14186 200 14242 800 6 chany_bottom_in[0]
port 3 nsew signal input
rlabel metal3 s 200 20408 800 20528 6 chany_bottom_in[10]
port 4 nsew signal input
rlabel metal3 s 200 22448 800 22568 6 chany_bottom_in[11]
port 5 nsew signal input
rlabel metal3 s 39200 5448 39800 5568 6 chany_bottom_in[12]
port 6 nsew signal input
rlabel metal3 s 39200 24488 39800 24608 6 chany_bottom_in[13]
port 7 nsew signal input
rlabel metal3 s 39200 26528 39800 26648 6 chany_bottom_in[14]
port 8 nsew signal input
rlabel metal2 s 39302 200 39358 800 6 chany_bottom_in[15]
port 9 nsew signal input
rlabel metal2 s 19982 39200 20038 39800 6 chany_bottom_in[16]
port 10 nsew signal input
rlabel metal3 s 200 31968 800 32088 6 chany_bottom_in[17]
port 11 nsew signal input
rlabel metal3 s 200 19048 800 19168 6 chany_bottom_in[18]
port 12 nsew signal input
rlabel metal2 s 36082 200 36138 800 6 chany_bottom_in[1]
port 13 nsew signal input
rlabel metal3 s 39200 7488 39800 7608 6 chany_bottom_in[2]
port 14 nsew signal input
rlabel metal2 s 9034 200 9090 800 6 chany_bottom_in[3]
port 15 nsew signal input
rlabel metal2 s 23202 39200 23258 39800 6 chany_bottom_in[4]
port 16 nsew signal input
rlabel metal3 s 39200 29928 39800 30048 6 chany_bottom_in[5]
port 17 nsew signal input
rlabel metal2 s 34150 200 34206 800 6 chany_bottom_in[6]
port 18 nsew signal input
rlabel metal2 s 34150 39200 34206 39800 6 chany_bottom_in[7]
port 19 nsew signal input
rlabel metal2 s 32218 200 32274 800 6 chany_bottom_in[8]
port 20 nsew signal input
rlabel metal2 s 27066 39200 27122 39800 6 chany_bottom_in[9]
port 21 nsew signal input
rlabel metal2 s 7102 39200 7158 39800 6 chany_bottom_out[0]
port 22 nsew signal output
rlabel metal2 s 18050 39200 18106 39800 6 chany_bottom_out[10]
port 23 nsew signal output
rlabel metal3 s 200 24488 800 24608 6 chany_bottom_out[11]
port 24 nsew signal output
rlabel metal3 s 39200 12928 39800 13048 6 chany_bottom_out[12]
port 25 nsew signal output
rlabel metal3 s 200 7488 800 7608 6 chany_bottom_out[13]
port 26 nsew signal output
rlabel metal3 s 200 30608 800 30728 6 chany_bottom_out[14]
port 27 nsew signal output
rlabel metal3 s 200 3408 800 3528 6 chany_bottom_out[15]
port 28 nsew signal output
rlabel metal3 s 200 14968 800 15088 6 chany_bottom_out[16]
port 29 nsew signal output
rlabel metal3 s 39200 28568 39800 28688 6 chany_bottom_out[17]
port 30 nsew signal output
rlabel metal3 s 39200 14968 39800 15088 6 chany_bottom_out[18]
port 31 nsew signal output
rlabel metal2 s 21270 39200 21326 39800 6 chany_bottom_out[1]
port 32 nsew signal output
rlabel metal3 s 39200 36048 39800 36168 6 chany_bottom_out[2]
port 33 nsew signal output
rlabel metal3 s 200 38088 800 38208 6 chany_bottom_out[3]
port 34 nsew signal output
rlabel metal2 s 28998 39200 29054 39800 6 chany_bottom_out[4]
port 35 nsew signal output
rlabel metal3 s 200 10888 800 11008 6 chany_bottom_out[5]
port 36 nsew signal output
rlabel metal2 s 1306 39200 1362 39800 6 chany_bottom_out[6]
port 37 nsew signal output
rlabel metal2 s 38014 39200 38070 39800 6 chany_bottom_out[7]
port 38 nsew signal output
rlabel metal3 s 200 34008 800 34128 6 chany_bottom_out[8]
port 39 nsew signal output
rlabel metal2 s 25134 200 25190 800 6 chany_bottom_out[9]
port 40 nsew signal output
rlabel metal3 s 39200 31968 39800 32088 6 chany_top_in[0]
port 41 nsew signal input
rlabel metal2 s 10322 39200 10378 39800 6 chany_top_in[10]
port 42 nsew signal input
rlabel metal2 s 3238 200 3294 800 6 chany_top_in[11]
port 43 nsew signal input
rlabel metal2 s 10322 200 10378 800 6 chany_top_in[12]
port 44 nsew signal input
rlabel metal2 s 30286 200 30342 800 6 chany_top_in[13]
port 45 nsew signal input
rlabel metal3 s 39200 10888 39800 11008 6 chany_top_in[14]
port 46 nsew signal input
rlabel metal3 s 39200 3408 39800 3528 6 chany_top_in[15]
port 47 nsew signal input
rlabel metal2 s 23202 200 23258 800 6 chany_top_in[16]
port 48 nsew signal input
rlabel metal2 s 18 39200 74 39800 6 chany_top_in[17]
port 49 nsew signal input
rlabel metal2 s 38014 200 38070 800 6 chany_top_in[18]
port 50 nsew signal input
rlabel metal2 s 12254 39200 12310 39800 6 chany_top_in[1]
port 51 nsew signal input
rlabel metal3 s 39200 8848 39800 8968 6 chany_top_in[2]
port 52 nsew signal input
rlabel metal3 s 200 1368 800 1488 6 chany_top_in[3]
port 53 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 chany_top_in[4]
port 54 nsew signal input
rlabel metal3 s 200 26528 800 26648 6 chany_top_in[5]
port 55 nsew signal input
rlabel metal3 s 200 9528 800 9648 6 chany_top_in[6]
port 56 nsew signal input
rlabel metal2 s 16118 39200 16174 39800 6 chany_top_in[7]
port 57 nsew signal input
rlabel metal2 s 18050 200 18106 800 6 chany_top_in[8]
port 58 nsew signal input
rlabel metal2 s 18 200 74 800 6 chany_top_in[9]
port 59 nsew signal input
rlabel metal3 s 200 17008 800 17128 6 chany_top_out[0]
port 60 nsew signal output
rlabel metal2 s 14186 39200 14242 39800 6 chany_top_out[10]
port 61 nsew signal output
rlabel metal2 s 25134 39200 25190 39800 6 chany_top_out[11]
port 62 nsew signal output
rlabel metal2 s 36082 39200 36138 39800 6 chany_top_out[12]
port 63 nsew signal output
rlabel metal3 s 200 28568 800 28688 6 chany_top_out[13]
port 64 nsew signal output
rlabel metal2 s 5170 200 5226 800 6 chany_top_out[14]
port 65 nsew signal output
rlabel metal2 s 1306 200 1362 800 6 chany_top_out[15]
port 66 nsew signal output
rlabel metal2 s 39302 39200 39358 39800 6 chany_top_out[16]
port 67 nsew signal output
rlabel metal2 s 30286 39200 30342 39800 6 chany_top_out[17]
port 68 nsew signal output
rlabel metal2 s 16118 200 16174 800 6 chany_top_out[18]
port 69 nsew signal output
rlabel metal3 s 39200 38088 39800 38208 6 chany_top_out[1]
port 70 nsew signal output
rlabel metal3 s 39200 1368 39800 1488 6 chany_top_out[2]
port 71 nsew signal output
rlabel metal2 s 5170 39200 5226 39800 6 chany_top_out[3]
port 72 nsew signal output
rlabel metal3 s 39200 20408 39800 20528 6 chany_top_out[4]
port 73 nsew signal output
rlabel metal2 s 7102 200 7158 800 6 chany_top_out[5]
port 74 nsew signal output
rlabel metal2 s 12254 200 12310 800 6 chany_top_out[6]
port 75 nsew signal output
rlabel metal2 s 19338 200 19394 800 6 chany_top_out[7]
port 76 nsew signal output
rlabel metal3 s 39200 22448 39800 22568 6 chany_top_out[8]
port 77 nsew signal output
rlabel metal2 s 21270 200 21326 800 6 chany_top_out[9]
port 78 nsew signal output
rlabel metal3 s 200 5448 800 5568 6 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 79 nsew signal output
rlabel metal2 s 32218 39200 32274 39800 6 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 80 nsew signal output
rlabel metal2 s 3238 39200 3294 39800 6 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 81 nsew signal output
rlabel metal2 s 9034 39200 9090 39800 6 pReset
port 82 nsew signal input
rlabel metal2 s 27066 200 27122 800 6 prog_clk
port 83 nsew signal input
rlabel metal3 s 200 12928 800 13048 6 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
port 84 nsew signal output
rlabel metal3 s 200 36048 800 36168 6 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 85 nsew signal output
rlabel metal3 s 39200 19048 39800 19168 6 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 86 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 88 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1259810
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/cby_1__1_/runs/22_12_30_10_10/results/signoff/cby_1__1_.magic.gds
string GDS_START 134360
<< end >>

