magic
tech sky130A
magscale 1 2
timestamp 1672416552
<< obsli1 >>
rect 1104 2159 36892 37553
<< obsm1 >>
rect 14 1912 37430 37584
<< metal2 >>
rect 1306 39200 1362 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 24490 39200 24546 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 7746 200 7802 800
rect 9678 200 9734 800
rect 10966 200 11022 800
rect 12898 200 12954 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 24490 200 24546 800
rect 26422 200 26478 800
rect 27710 200 27766 800
rect 29642 200 29698 800
rect 30930 200 30986 800
rect 32862 200 32918 800
rect 34150 200 34206 800
rect 36082 200 36138 800
<< obsm2 >>
rect 20 39144 1250 39545
rect 1418 39144 3182 39545
rect 3350 39144 4470 39545
rect 4638 39144 6402 39545
rect 6570 39144 7690 39545
rect 7858 39144 9622 39545
rect 9790 39144 10910 39545
rect 11078 39144 12842 39545
rect 13010 39144 14774 39545
rect 14942 39144 16062 39545
rect 16230 39144 17994 39545
rect 18162 39144 19282 39545
rect 19450 39144 21214 39545
rect 21382 39144 22502 39545
rect 22670 39144 24434 39545
rect 24602 39144 26366 39545
rect 26534 39144 27654 39545
rect 27822 39144 29586 39545
rect 29754 39144 30874 39545
rect 31042 39144 32806 39545
rect 32974 39144 34094 39545
rect 34262 39144 36026 39545
rect 36194 39144 37314 39545
rect 20 856 37424 39144
rect 130 144 1250 856
rect 1418 144 3182 856
rect 3350 144 4470 856
rect 4638 144 6402 856
rect 6570 144 7690 856
rect 7858 144 9622 856
rect 9790 144 10910 856
rect 11078 144 12842 856
rect 13010 144 14774 856
rect 14942 144 16062 856
rect 16230 144 17994 856
rect 18162 144 19282 856
rect 19450 144 21214 856
rect 21382 144 22502 856
rect 22670 144 24434 856
rect 24602 144 26366 856
rect 26534 144 27654 856
rect 27822 144 29586 856
rect 29754 144 30874 856
rect 31042 144 32806 856
rect 32974 144 34094 856
rect 34262 144 36026 856
rect 36194 144 37424 856
rect 20 31 37424 144
<< metal3 >>
rect 200 39448 800 39568
rect 200 38088 800 38208
rect 37200 38088 37800 38208
rect 200 36048 800 36168
rect 37200 36048 37800 36168
rect 200 34688 800 34808
rect 37200 34688 37800 34808
rect 200 32648 800 32768
rect 37200 32648 37800 32768
rect 200 31288 800 31408
rect 37200 31288 37800 31408
rect 200 29248 800 29368
rect 37200 29248 37800 29368
rect 200 27888 800 28008
rect 37200 27888 37800 28008
rect 200 25848 800 25968
rect 37200 25848 37800 25968
rect 200 23808 800 23928
rect 37200 23808 37800 23928
rect 200 22448 800 22568
rect 37200 22448 37800 22568
rect 200 20408 800 20528
rect 37200 20408 37800 20528
rect 200 19048 800 19168
rect 37200 19048 37800 19168
rect 200 17008 800 17128
rect 37200 17008 37800 17128
rect 200 15648 800 15768
rect 37200 15648 37800 15768
rect 200 13608 800 13728
rect 37200 13608 37800 13728
rect 200 11568 800 11688
rect 37200 11568 37800 11688
rect 200 10208 800 10328
rect 37200 10208 37800 10328
rect 200 8168 800 8288
rect 37200 8168 37800 8288
rect 200 6808 800 6928
rect 37200 6808 37800 6928
rect 200 4768 800 4888
rect 37200 4768 37800 4888
rect 200 3408 800 3528
rect 37200 3408 37800 3528
rect 200 1368 800 1488
rect 37200 1368 37800 1488
rect 37200 8 37800 128
<< obsm3 >>
rect 880 39368 37200 39541
rect 800 38288 37200 39368
rect 880 38008 37120 38288
rect 800 36248 37200 38008
rect 880 35968 37120 36248
rect 800 34888 37200 35968
rect 880 34608 37120 34888
rect 800 32848 37200 34608
rect 880 32568 37120 32848
rect 800 31488 37200 32568
rect 880 31208 37120 31488
rect 800 29448 37200 31208
rect 880 29168 37120 29448
rect 800 28088 37200 29168
rect 880 27808 37120 28088
rect 800 26048 37200 27808
rect 880 25768 37120 26048
rect 800 24008 37200 25768
rect 880 23728 37120 24008
rect 800 22648 37200 23728
rect 880 22368 37120 22648
rect 800 20608 37200 22368
rect 880 20328 37120 20608
rect 800 19248 37200 20328
rect 880 18968 37120 19248
rect 800 17208 37200 18968
rect 880 16928 37120 17208
rect 800 15848 37200 16928
rect 880 15568 37120 15848
rect 800 13808 37200 15568
rect 880 13528 37120 13808
rect 800 11768 37200 13528
rect 880 11488 37120 11768
rect 800 10408 37200 11488
rect 880 10128 37120 10408
rect 800 8368 37200 10128
rect 880 8088 37120 8368
rect 800 7008 37200 8088
rect 880 6728 37120 7008
rect 800 4968 37200 6728
rect 880 4688 37120 4968
rect 800 3608 37200 4688
rect 880 3328 37120 3608
rect 800 1568 37200 3328
rect 880 1288 37120 1568
rect 800 208 37200 1288
rect 800 35 37120 208
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 14963 2347 19488 37093
rect 19968 2347 27725 37093
<< labels >>
rlabel metal2 s 34150 39200 34206 39800 6 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
port 1 nsew signal output
rlabel metal3 s 37200 25848 37800 25968 6 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
port 2 nsew signal output
rlabel metal2 s 36082 200 36138 800 6 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
port 3 nsew signal output
rlabel metal2 s 14830 200 14886 800 6 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
port 4 nsew signal output
rlabel metal2 s 26422 39200 26478 39800 6 ccff_head
port 5 nsew signal input
rlabel metal3 s 37200 10208 37800 10328 6 ccff_tail
port 6 nsew signal output
rlabel metal2 s 12898 39200 12954 39800 6 chanx_left_in[0]
port 7 nsew signal input
rlabel metal2 s 16118 39200 16174 39800 6 chanx_left_in[10]
port 8 nsew signal input
rlabel metal3 s 37200 27888 37800 28008 6 chanx_left_in[11]
port 9 nsew signal input
rlabel metal3 s 200 38088 800 38208 6 chanx_left_in[12]
port 10 nsew signal input
rlabel metal3 s 37200 31288 37800 31408 6 chanx_left_in[13]
port 11 nsew signal input
rlabel metal2 s 19338 39200 19394 39800 6 chanx_left_in[14]
port 12 nsew signal input
rlabel metal3 s 37200 34688 37800 34808 6 chanx_left_in[15]
port 13 nsew signal input
rlabel metal3 s 200 4768 800 4888 6 chanx_left_in[16]
port 14 nsew signal input
rlabel metal3 s 200 1368 800 1488 6 chanx_left_in[17]
port 15 nsew signal input
rlabel metal3 s 37200 36048 37800 36168 6 chanx_left_in[18]
port 16 nsew signal input
rlabel metal3 s 37200 32648 37800 32768 6 chanx_left_in[1]
port 17 nsew signal input
rlabel metal3 s 200 32648 800 32768 6 chanx_left_in[2]
port 18 nsew signal input
rlabel metal3 s 37200 4768 37800 4888 6 chanx_left_in[3]
port 19 nsew signal input
rlabel metal2 s 1306 39200 1362 39800 6 chanx_left_in[4]
port 20 nsew signal input
rlabel metal3 s 200 20408 800 20528 6 chanx_left_in[5]
port 21 nsew signal input
rlabel metal2 s 27710 200 27766 800 6 chanx_left_in[6]
port 22 nsew signal input
rlabel metal3 s 200 19048 800 19168 6 chanx_left_in[7]
port 23 nsew signal input
rlabel metal3 s 37200 29248 37800 29368 6 chanx_left_in[8]
port 24 nsew signal input
rlabel metal3 s 37200 8 37800 128 6 chanx_left_in[9]
port 25 nsew signal input
rlabel metal2 s 22558 39200 22614 39800 6 chanx_left_out[0]
port 26 nsew signal output
rlabel metal3 s 200 39448 800 39568 6 chanx_left_out[10]
port 27 nsew signal output
rlabel metal3 s 37200 17008 37800 17128 6 chanx_left_out[11]
port 28 nsew signal output
rlabel metal3 s 200 15648 800 15768 6 chanx_left_out[12]
port 29 nsew signal output
rlabel metal2 s 7746 200 7802 800 6 chanx_left_out[13]
port 30 nsew signal output
rlabel metal3 s 37200 20408 37800 20528 6 chanx_left_out[14]
port 31 nsew signal output
rlabel metal2 s 14830 39200 14886 39800 6 chanx_left_out[15]
port 32 nsew signal output
rlabel metal3 s 37200 8168 37800 8288 6 chanx_left_out[16]
port 33 nsew signal output
rlabel metal2 s 24490 39200 24546 39800 6 chanx_left_out[17]
port 34 nsew signal output
rlabel metal2 s 37370 39200 37426 39800 6 chanx_left_out[18]
port 35 nsew signal output
rlabel metal2 s 34150 200 34206 800 6 chanx_left_out[1]
port 36 nsew signal output
rlabel metal2 s 18050 39200 18106 39800 6 chanx_left_out[2]
port 37 nsew signal output
rlabel metal2 s 30930 200 30986 800 6 chanx_left_out[3]
port 38 nsew signal output
rlabel metal3 s 200 3408 800 3528 6 chanx_left_out[4]
port 39 nsew signal output
rlabel metal2 s 10966 200 11022 800 6 chanx_left_out[5]
port 40 nsew signal output
rlabel metal3 s 200 27888 800 28008 6 chanx_left_out[6]
port 41 nsew signal output
rlabel metal3 s 37200 15648 37800 15768 6 chanx_left_out[7]
port 42 nsew signal output
rlabel metal2 s 4526 200 4582 800 6 chanx_left_out[8]
port 43 nsew signal output
rlabel metal3 s 200 13608 800 13728 6 chanx_left_out[9]
port 44 nsew signal output
rlabel metal3 s 200 31288 800 31408 6 chanx_right_in[0]
port 45 nsew signal input
rlabel metal3 s 200 6808 800 6928 6 chanx_right_in[10]
port 46 nsew signal input
rlabel metal3 s 200 29248 800 29368 6 chanx_right_in[11]
port 47 nsew signal input
rlabel metal2 s 6458 39200 6514 39800 6 chanx_right_in[12]
port 48 nsew signal input
rlabel metal2 s 3238 200 3294 800 6 chanx_right_in[13]
port 49 nsew signal input
rlabel metal2 s 9678 200 9734 800 6 chanx_right_in[14]
port 50 nsew signal input
rlabel metal2 s 32862 200 32918 800 6 chanx_right_in[15]
port 51 nsew signal input
rlabel metal3 s 37200 13608 37800 13728 6 chanx_right_in[16]
port 52 nsew signal input
rlabel metal3 s 37200 6808 37800 6928 6 chanx_right_in[17]
port 53 nsew signal input
rlabel metal2 s 24490 200 24546 800 6 chanx_right_in[18]
port 54 nsew signal input
rlabel metal3 s 200 36048 800 36168 6 chanx_right_in[1]
port 55 nsew signal input
rlabel metal3 s 37200 1368 37800 1488 6 chanx_right_in[2]
port 56 nsew signal input
rlabel metal3 s 200 8168 800 8288 6 chanx_right_in[3]
port 57 nsew signal input
rlabel metal3 s 37200 11568 37800 11688 6 chanx_right_in[4]
port 58 nsew signal input
rlabel metal3 s 200 23808 800 23928 6 chanx_right_in[5]
port 59 nsew signal input
rlabel metal2 s 29642 200 29698 800 6 chanx_right_in[6]
port 60 nsew signal input
rlabel metal3 s 200 17008 800 17128 6 chanx_right_in[7]
port 61 nsew signal input
rlabel metal2 s 9678 39200 9734 39800 6 chanx_right_in[8]
port 62 nsew signal input
rlabel metal2 s 4526 39200 4582 39800 6 chanx_right_in[9]
port 63 nsew signal input
rlabel metal2 s 18050 200 18106 800 6 chanx_right_out[0]
port 64 nsew signal output
rlabel metal2 s 18 200 74 800 6 chanx_right_out[10]
port 65 nsew signal output
rlabel metal2 s 22558 200 22614 800 6 chanx_right_out[11]
port 66 nsew signal output
rlabel metal2 s 10966 39200 11022 39800 6 chanx_right_out[12]
port 67 nsew signal output
rlabel metal2 s 21270 39200 21326 39800 6 chanx_right_out[13]
port 68 nsew signal output
rlabel metal2 s 32862 39200 32918 39800 6 chanx_right_out[14]
port 69 nsew signal output
rlabel metal3 s 200 25848 800 25968 6 chanx_right_out[15]
port 70 nsew signal output
rlabel metal3 s 200 22448 800 22568 6 chanx_right_out[16]
port 71 nsew signal output
rlabel metal2 s 1306 200 1362 800 6 chanx_right_out[17]
port 72 nsew signal output
rlabel metal2 s 36082 39200 36138 39800 6 chanx_right_out[18]
port 73 nsew signal output
rlabel metal2 s 27710 39200 27766 39800 6 chanx_right_out[1]
port 74 nsew signal output
rlabel metal2 s 16118 200 16174 800 6 chanx_right_out[2]
port 75 nsew signal output
rlabel metal3 s 37200 38088 37800 38208 6 chanx_right_out[3]
port 76 nsew signal output
rlabel metal3 s 37200 3408 37800 3528 6 chanx_right_out[4]
port 77 nsew signal output
rlabel metal3 s 200 10208 800 10328 6 chanx_right_out[5]
port 78 nsew signal output
rlabel metal3 s 37200 22448 37800 22568 6 chanx_right_out[6]
port 79 nsew signal output
rlabel metal2 s 6458 200 6514 800 6 chanx_right_out[7]
port 80 nsew signal output
rlabel metal2 s 12898 200 12954 800 6 chanx_right_out[8]
port 81 nsew signal output
rlabel metal2 s 19338 200 19394 800 6 chanx_right_out[9]
port 82 nsew signal output
rlabel metal3 s 37200 23808 37800 23928 6 pReset
port 83 nsew signal input
rlabel metal2 s 21270 200 21326 800 6 prog_clk
port 84 nsew signal input
rlabel metal2 s 30930 39200 30986 39800 6 top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
port 85 nsew signal output
rlabel metal2 s 29642 39200 29698 39800 6 top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_
port 86 nsew signal output
rlabel metal2 s 3238 39200 3294 39800 6 top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_
port 87 nsew signal output
rlabel metal2 s 7746 39200 7802 39800 6 top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_
port 88 nsew signal output
rlabel metal2 s 26422 200 26478 800 6 top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_
port 89 nsew signal output
rlabel metal3 s 200 11568 800 11688 6 top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_
port 90 nsew signal output
rlabel metal3 s 200 34688 800 34808 6 top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_
port 91 nsew signal output
rlabel metal3 s 37200 19048 37800 19168 6 top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_
port 92 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 93 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 93 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 94 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 38000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1937274
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/cbx_1__4_/runs/22_12_30_10_08/results/signoff/cbx_1__4_.magic.gds
string GDS_START 152304
<< end >>

